�NUMPY v {'descr': '<f8', 'fortran_order': False, 'shape': (3, 10000, 5), }                                                   
������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�%@=��ٿ}��
 ��@�ݰ��3@�`��L�!?ExxL��@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�F��ٿ�f�����@�i���3@&�� �!?�����@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�IK��ٿړ�����@Tg���3@�o��!?������@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@�ۙٿ�������@U�Ӝ��3@Q]�F;�!?��^���@m��ؙٿ�v�����@B�c��3@��VC�!?µ����@m��ؙٿ�v�����@B�c��3@��VC�!?µ����@m��ؙٿ�v�����@B�c��3@��VC�!?µ����@m��ؙٿ�v�����@B�c��3@��VC�!?µ����@m��ؙٿ�v�����@B�c��3@��VC�!?µ����@^x3�Йٿ.d,����@�JG���3@�<3e�!?'����@^x3�Йٿ.d,����@�JG���3@�<3e�!?'����@^x3�Йٿ.d,����@�JG���3@�<3e�!?'����@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@��kؙٿFZ�����@����3@3��q�!?��  ��@O�c9ڙٿ�������@a�\���3@�YT�I�!? �i���@⻽Gיٿ	�����@K^��  4@-�u�!?A�d���@⻽Gיٿ	�����@K^��  4@-�u�!?A�d���@⻽Gיٿ	�����@K^��  4@-�u�!?A�d���@��eT�ٿ�+����@S*|��3@6�ݏ!?v�����@��eT�ٿ�+����@S*|��3@6�ݏ!?v�����@��eT�ٿ�+����@S*|��3@6�ݏ!?v�����@����ٿ������@[�'  4@�
�	�!?�UH���@��Z��ٿ9q9����@Z�����3@
�Ȱ�!?�C���@��Z��ٿ9q9����@Z�����3@
�Ȱ�!?�C���@|)�ܙٿ2�J����@�&����3@~FQ�p�!?i�����@|)�ܙٿ2�J����@�&����3@~FQ�p�!?i�����@|)�ܙٿ2�J����@�&����3@~FQ�p�!?i�����@q9f��ٿ}������@�d%  4@�*o�b�!?_�B���@q9f��ٿ}������@�d%  4@�*o�b�!?_�B���@q9f��ٿ}������@�d%  4@�*o�b�!?_�B���@q9f��ٿ}������@�d%  4@�*o�b�!?_�B���@q9f��ٿ}������@�d%  4@�*o�b�!?_�B���@��-ܙٿ�*־���@�4�  4@X�ߌ�!?6%O���@��-ܙٿ�*־���@�4�  4@X�ߌ�!?6%O���@��7��ٿ1	����@D;0���3@y��+2�!?�j����@��N�ٿ<�����@��RI��3@�r.�>�!?hE���@k���ٿ�n�����@~����3@ȧ���!?�ꃿ��@_����ٿ`�m����@������3@|-1�[�!?��-���@�V���ٿ�U׺���@��3���3@CY�!?'B����@�V���ٿ�U׺���@��3���3@CY�!?'B����@\rD#�ٿ��a����@�����3@BQO�;�!?����@\rD#�ٿ��a����@�����3@BQO�;�!?����@�!ax�ٿIڳ����@�w'4��3@k#d�!?�@[���@A@�;ߙٿ�H_����@U����3@R-W�!?��m���@A@�;ߙٿ�H_����@U����3@R-W�!?��m���@A@�;ߙٿ�H_����@U����3@R-W�!?��m���@G3ݙٿ4������@�<U���3@>z�C�!?�2P���@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@x�0�ޙٿ]������@�#e��3@�ằ`�!?�����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@:h%�ٿ�}�����@��ق��3@�9),��!?�[����@���^ޙٿ�9�����@�à{��3@�H~L��!?o@����@?���יٿ�������@\Z����3@�/CL�!?0y'���@?���יٿ�������@\Z����3@�/CL�!?0y'���@GNәٿW������@ҪZ���3@���$�!?�<����@GNәٿW������@ҪZ���3@���$�!?�<����@��vԙٿ��c����@�;���3@	��r�!?��m���@W�3יٿ8������@!RR��3@���z�!?P�����@z��ٙٿ~������@[����3@

�7T�!?��A���@z��ٙٿ~������@[����3@

�7T�!?��A���@o�ʒיٿ�xy����@��w��3@�)v�!?Y�D���@w8��ٙٿ04�����@i>�S��3@0b��L�!?����@w8��ٙٿ04�����@i>�S��3@0b��L�!?����@���ۙٿ��Q����@� ���3@| %2�!?l�N���@t~�uܙٿ*%�����@D~-���3@t_��!?p���@����ܙٿ�jR����@�	����3@�<%�ڏ!?�c^���@����ܙٿ�jR����@�	����3@�<%�ڏ!?�c^���@U��ۙٿ������@�AT��3@&���!?�5����@�4�Oݙٿ������@?����3@�~�l3�!?�#����@)� �ٿT�����@��$:��3@�@��}�!?������@)� �ٿT�����@��$:��3@�@��}�!?������@)� �ٿT�����@��$:��3@�@��}�!?������@�	�ٿ+\ο���@({k���3@Ϣ�J�!?q�����@V��H�ٿ�&�����@vɾ���3@JUm�!?*����@V��H�ٿ�&�����@vɾ���3@JUm�!?*����@i��H�ٿ�z����@Q-2���3@"5g�!?5����@��b��ٿ4�˻���@�7���3@2�D�!?�1C���@��b��ٿ4�˻���@�7���3@2�D�!?�1C���@��b��ٿ4�˻���@�7���3@2�D�!?�1C���@��b��ٿ4�˻���@�7���3@2�D�!?�1C���@��#�ٿLD����@�b���3@����G�!?�l����@�]��ٿ�YA����@B0����3@!�u�<�!?�ۺ��@P���ٿѴ6����@vr:���3@PP8�!?�����@�!�6�ٿw�R����@�q�(��3@�/�e�!?��C���@�!�6�ٿw�R����@�q�(��3@�/�e�!?��C���@5
���ٿ������@�����3@����?�!?��	���@5
���ٿ������@�����3@����?�!?��	���@-����ٿ������@'����3@Q�0r*�!?�����@�'H�ٿQ�7����@����3@�6Ԉ�!?��y���@�'H�ٿQ�7����@����3@�6Ԉ�!?��y���@�'H�ٿQ�7����@����3@�6Ԉ�!?��y���@y8��ٿ_�����@mvÖ��3@j��U��!?tR����@� >��ٿ�(ܴ���@��N��3@�`>�!?�4���@㸍�ٿ.�����@�_Ii��3@o5o�v�!?�dT���@ lП�ٿ��д���@?�����3@��ٮ��!?�����@�΢��ٿ�/����@Z�d���3@��O]�!?d����@8[���ٿ4۴���@���)��3@Xp4��!?a����@��`�ٿ(���@�`�(��3@�T�"��!?7D����@��Z��ٿI�����@��@��3@<�W�|�!?N՛���@;�1d��ٿU`<����@�*U���3@f���!?������@�Y��ߙٿ�nٶ���@N4m��3@i7�Z�!?����@�vG���ٿ{�t����@gK_���3@�~̧`�!?�|����@�_�ٿ4�F����@v_�C  4@�����!?�b���@�_�ٿ4�F����@v_�C  4@�����!?�b���@�KɎ��ٿ<�ڶ���@�0�  4@�z�Tu�!?�-����@�|�ٿ�:����@���+ 4@�l�!?�����@[���ٿ?������@ض�y 4@O��s�!?����@?"I�ٿ �����@U'3 4@�	�!?8���@?"I�ٿ �����@U'3 4@�	�!?8���@����ٿ��_����@�ڶ  4@�X+�!?�|����@�����ٿKw����@wC;}  4@T�`7<�!?2�j���@�����ٿKw����@wC;}  4@T�`7<�!?2�j���@�����ٿKw����@wC;}  4@T�`7<�!?2�j���@,��H�ٿ-�
����@ʧg@  4@v��lQ�!?h����@,��H�ٿ-�
����@ʧg@  4@v��lQ�!?h����@|
�ٿ�="����@�e���3@��dC~�!?��@���@R�z��ٿ}.C����@�>��3@���p�!?[�f���@�yJs�ٿ�x�����@8�B���3@�Gl]�!?�J����@�u�O�ٿ�8�����@yu�H  4@G����!?�(����@�4$�ٿ7a�����@�7�t  4@�}X�#�!?������@��|�ٿ̐J����@�|X��3@,J�I��!?����@ӱ"&�ٿ7�����@1)z��3@t�߁��!?����@���ٿ��.����@�6l���3@a0��g�!?��)���@�W�d�ٿ7Q9����@����3@q<�Y�!?v/����@iBd�ٿ2V����@�ށN��3@��!�+�!?�����@���l�ٿ
�]����@/�Fh��3@�Z�~R�!?bN����@�9�)�ٿ _#����@�s����3@ϹX|��!?�I����@�9�)�ٿ _#����@�s����3@ϹX|��!?�I����@���ٿM����@� ����3@Qp��V�!?>J-���@�Z���ٿR������@ӿ����3@9�t8�!?1�X���@����ٿ7Nh����@��O���3@B1,�!?��R���@�hR�ٿBb����@�o  4@{h�'�!?�>|���@׸&�ٿ��'����@�/����3@!�*�!?�f����@5d��ٿ�������@��ax��3@�X��!?II���@���ٿ�<����@@.���3@�Lg�_�!?i r���@���ٿ�����@��{^��3@�q�q�!?�n���@��`�ٿ������@?����3@H�ڇ��!?��U���@x�e��ٿ�������@������3@�d�S��!?�ץ���@jɮ��ٿX�����@GUp��3@wX�`�!?�g���@�����ٿ��8����@G'����3@���@�!?<4X���@�jQ��ٿE죿���@G�F$��3@v��&�!?Ɯ����@�*|8�ٿ;G�����@���g��3@�d�8�!?�*���@&�?��ٿZ�4����@����3@�ق�!?�l���@��R�ٿ�&�����@]��?��3@��Zn�!?�� ���@U�	r�ٿ�����@�j��3@F<�@�!?������@��|��ٿWƽ���@�9����3@��3��!?�����@�c?.ߙٿ�P�����@�
����3@Y�j*�!?h����@-jV��ٿ2�I����@0l\��3@k���7�!?v-����@�A�&�ٿ.ua����@��R��3@ayy'f�!?7k���@�Q��ٿ�o�����@�q��3@�6U-��!?fe,���@J�O��ٿH�t����@\]���3@�����!?�(����@�,���ٿb�,����@9w����3@)^"��!?z"����@�m�m�ٿ%����@*t,  4@\�}��!?+�����@T�K��ٿsR˻���@(�.  4@�WNs�!?�Z����@�Ǌ.�ٿ�/;����@�Y]u  4@��_�!?�`h���@*-��ٿmx�����@Zy  4@�d 7�!?�x����@nǌP�ٿ�fc����@�0[���3@j��G�!?
�����@ń��ٿ	������@��m���3@��IPD�!?������@��|�ٿ�5����@V�  4@���R�!?`%���@��|�ٿ�5����@V�  4@���R�!?`%���@��j�ٿ�<����@�S��  4@f5Vi9�!?�;���@Hb�Eߙٿ=E�����@�U��  4@E�\�e�!?������@�x�ڙٿ�-@����@u��  4@B�7�l�!?׍���@��V�֙ٿ��n����@�gu  4@�O����!?�k}���@� �֙ٿM�L����@4��  4@�5�!?)����@�ި�ϙٿ_�M����@|WR5 4@6;-���!?������@�>�|Йٿ��V����@c h 4@e��I��!?y����@�>�|Йٿ��V����@c h 4@e��I��!?y����@QηљٿZ�G����@��� 4@�~3���!?:,��@QηљٿZ�G����@��� 4@�~3���!?:,��@`�{Uәٿ�Ա����@Ч�� 4@���G͐!?���7��@FE��̙ٿR�����@�ǌ< 4@�\��!?.kA<��@FE��̙ٿR�����@�ǌ< 4@�\��!?.kA<��@�١ٿ��2����@���� 4@:�6̐!?�e�O��@J$�[ęٿ�v����@퇱� 4@�X��}�!?���C��@J$�[ęٿ�v����@퇱� 4@�X��}�!?���C��@�]h��ٿW�����@[�w 4@��3��!?"T��@��]ϵ�ٿ�Z�����@��G� 4@�(��!?g�6:��@ �R-��ٿD8�����@z7^ 4@���oo�!?�~1��@ �R-��ٿD8�����@z7^ 4@���oo�!?�~1��@����ٿ6�����@ptMZ 4@��ᛊ�!?�/��@'u赙ٿj�:����@sH�� 4@�d|��!?���+��@
����ٿ�����@p�j; 4@�^�Ɛ!?��D6��@ߤ�V��ٿ�s4����@Wbu 4@F:R�ߐ!?t�gD��@�ˤ�ٿ�°����@��I 4@dE���!?Q�y��@�=aÙٿ��հ���@��� 4@�.x��!?���(��@�=aÙٿ��հ���@��� 4@�.x��!?���(��@�=aÙٿ��հ���@��� 4@�.x��!?���(��@n}�Ǚٿ��s����@*��� 4@�'i��!?�y���@�S=Ùٿ�3����@^�s 4@A��U��!?7��@���lșٿ�к���@bp(> 4@��-p�!?5�����@��ϙٿVDϼ���@��܄��3@`;�L�!?�7���@A|>�ϙٿyMý���@4����3@u��o5�!?k���@�j�0��ٿ�� ����@����  4@M}l q�!?S����@�ӂ���ٿP	c����@�0��  4@s9�L�!?����@=dg��ٿ�j�����@c: 4@.	�v��!?�n5��@=dg��ٿ�j�����@c: 4@.	�v��!?�n5��@��A��ٿ�d����@$�� 4@e����!?6����@	ûO��ٿb�����@(�I 4@�}�䝐!?�E���@	ûO��ٿb�����@(�I 4@�}�䝐!?�E���@v�����ٿ�ֻ����@8� 4@�m��!?��,��@v�����ٿ�ֻ����@8� 4@�m��!?��,��@l�c��ٿ�������@��-/ 4@����ː!?	S��@��GК�ٿ����@���f 4@��!?��zj��@��GК�ٿ����@���f 4@��!?��zj��@��GК�ٿ����@���f 4@��!?��zj��@��GК�ٿ����@���f 4@��!?��zj��@+�Ne��ٿ7�M����@!+f 4@`N���!?������@+�Ne��ٿ7�M����@!+f 4@`N���!?������@+�Ne��ٿ7�M����@!+f 4@`N���!?������@s'�<��ٿ��5����@Y52� 4@z��!?�ڸB��@uݧ�ܙٿ:����@�o� 4@��d���!?�G�C��@��OיٿTI����@l� 4@���^�!?o�\U��@��OיٿTI����@l� 4@���^�!?o�\U��@����ٿ�Ի����@(�g 4@��3�!?_?�{��@����ٿ�Ի����@(�g 4@��3�!?_?�{��@��-��ٿV������@~�� 4@�$d�U�!?Ӓ����@�W���ٿ�
����@_�!� 4@�fI�0�!?K�l��@����ٿ�
N����@��~ 4@lr�M �!?C6wF��@v �'�ٿY�����@��m�  4@բ-�k�!?�q���@��e7��ٿ0�պ���@Ф��  4@���}�!?Jl%��@�dv�)�ٿ�|�����@AY�	��3@��
WP�!?��5#��@v��$�ٿ<ª����@h�]g��3@��(bS�!?�����@����f�ٿ������@��@��3@-�r
>�!?��%��@I:C]:�ٿ�[����@�����3@��S�!?�����@I:C]:�ٿ�[����@�����3@��S�!?�����@/��p�ٿٚp����@�}?y��3@'�:�!?�bC���@��v(=�ٿ�ӑ����@�����3@��1�!?[�}X��@w���ٿ�h�����@��:���3@v�턔�!?�uxb��@1h�ԙٿ�A����@��&���3@�;���!?�u�v��@1h�ԙٿ�A����@��&���3@�;���!?�u�v��@�ͧ:יٿ��/����@t"����3@Fڂw��!?��%��@�ͧ:יٿ��/����@t"����3@Fڂw��!?��%��@�wО��ٿ˓.����@�I����3@v��̓�!?�S���@����ٿn�G����@;�$��3@�kۜP�!?÷����@����ٿn�G����@;�$��3@�kۜP�!?÷����@�.�Uڙٿ��_����@ ����3@8&�gp�!?/. l��@J���ٿLOr����@/�W��3@�o�Y�!?�ʼ��@Qe|��ٿ@�%����@���k��3@�8�/�!?y�`$��@��7�'�ٿTC����@�����3@�e��s�!?*<�k��@g�C�ٙٿK�����@��Ÿ��3@^ZzG��!?����@3����ٿO������@��ƴ��3@���r�!?�m��@�����ٿ6������@�$,8��3@E�w�[�!?S2�2��@�����ٿ6������@�$,8��3@E�w�[�!?S2�2��@�<.S�ٿDcw ��@�Hx��3@��qt?�!?�r6��@��w��ٿ>�c! ��@�\�=��3@�3]�!?r`���@���ٚٿf#@& ��@�Sֿ�3@ո�$�!?>�b��@�Ov��ٿq�~! ��@
�%���3@�كP�!?������@��m�h�ٿ�TyW ��@�P�d��3@�ƦFj�!?��]���@8�E"x�ٿxb�W ��@H��ܠ�3@	���!?�e����@t[b��ٿ�F<K ��@(�����3@q��?�!?V�d���@����ٿjQ�D ��@o��`��3@Z�@�!?��Z��@>���K�ٿ<G ��@������3@�����!?�����@|/�#�ٿ�� ��@�>��3@%��|��!?�B��@��q<.�ٿf�9����@�s��3@p9e���!?����@�Q�}��ٿ������@�uj" 4@�~z��!?�c_���@��ݯ�ٿK����@ ����3@Y0��F�!?�g���@��ݯ�ٿK����@ ����3@Y0��F�!?�g���@��ݯ�ٿK����@ ����3@Y0��F�!?�g���@��a$��ٿ�������@)-H��3@���n�!?�->���@F�1�D�ٿc�t����@��K���3@���w�!?Ů�5��@F�1�D�ٿc�t����@��K���3@���w�!?Ů�5��@F�1�D�ٿc�t����@��K���3@���w�!?Ů�5��@h: �5�ٿ	�}����@z���3@�=߉�!?+�q��@h: �5�ٿ	�}����@z���3@�=߉�!?+�q��@h: �5�ٿ	�}����@z���3@�=߉�!?+�q��@���^��ٿ5�J���@ ��S 4@�ucxB�!?�~����@�1��ߘٿ-@���@�M,| 4@��)0E�!?
] ]��@�1��ߘٿ-@���@�M,| 4@��)0E�!?
] ]��@]6/ޘٿ������@H��e 4@^2��!?L<��@]6/ޘٿ������@H��e 4@^2��!?L<��@]6/ޘٿ������@H��e 4@^2��!?L<��@� U��ٿLږ����@Vy� 4@44�U*�!?c�=��@� U��ٿLږ����@Vy� 4@44�U*�!?c�=��@� U��ٿLږ����@Vy� 4@44�U*�!?c�=��@��vAǘٿp%�����@wL�Ĩ 4@6�o�!?�����@F�KY]�ٿ�� 8���@)���\ 4@3ٜ�0�!?c���@F�KY]�ٿ�� 8���@)���\ 4@3ٜ�0�!?c���@�Cw%�ٿ-w�	���@@A�{ 4@�g6G�!?ݼ���@�Cw%�ٿ-w�	���@@A�{ 4@�g6G�!?ݼ���@���?+�ٿ�y���@:���� 4@�t1s!�!?׃<��@���?+�ٿ�y���@:���� 4@�t1s!�!?׃<��@]L�]H�ٿ0!�;���@%��=O 4@���Q�!?0�Q_��@]L�]H�ٿ0!�;���@%��=O 4@���Q�!?0�Q_��@Md#�#�ٿymJ^���@�C�2 4@6_i�C�!?��t~��@<��<��ٿ��T���@{ղ�0 4@�����!?��J��@<��<��ٿ��T���@{ղ�0 4@�����!?��J��@<��<��ٿ��T���@{ղ�0 4@�����!?��J��@�;��A�ٿ�!%����@�xe� 4@�}�	#�!?��ˏ��@�;��A�ٿ�!%����@�xe� 4@�}�	#�!?��ˏ��@�;��A�ٿ�!%����@�xe� 4@�}�	#�!?��ˏ��@�;��A�ٿ�!%����@�xe� 4@�}�	#�!?��ˏ��@2Γ��ٿ������@��w 4@�C+�A�!?�R!a��@{�KE�ٿ��/d���@HP=�& 4@4"��!?������@#�YA�ٿ�c�����@����^ 4@��=��!?�����@�"8a�ٿ�$4���@Ye��< 4@���ᒐ!?4�����@��yM��ٿ����@GTe 4@2 ��>�!?����@��yM��ٿ����@GTe 4@2 ��>�!?����@�D�&��ٿ������@�܄� 4@zN%�!?��j=��@�D�&��ٿ������@�܄� 4@zN%�!?��j=��@��6�B�ٿb�~���@S���� 4@�B��!?�n�u�@�ך��ٿ���.���@-+w)B 4@j��$P�!?��+���@w�
!�ٿ�wg���@��t& 4@�61�f�!?d�c;��@��4�ٿ�a,���@�}$= 4@�_.%W�!?��d��@<ʆH-�ٿJaO���@疧 4@<P�no�!?�-~��@<ʆH-�ٿJaO���@疧 4@<P�no�!?�-~��@<ʆH-�ٿJaO���@疧 4@<P�no�!?�-~��@<ʆH-�ٿJaO���@疧 4@<P�no�!?�-~��@<ʆH-�ٿJaO���@疧 4@<P�no�!?�-~��@K�wŘٿa�͙���@ӖG���3@ɧWx�!?�>����@K�wŘٿa�͙���@ӖG���3@ɧWx�!?�>����@K�wŘٿa�͙���@ӖG���3@ɧWx�!?�>����@K�wŘٿa�͙���@ӖG���3@ɧWx�!?�>����@Z�Y�,�ٿ&�w���@"����3@a��L��!?��w��@ƻӢ��ٿ�� ��@k���3@�ʹ���!?��fX��@ƻӢ��ٿ�� ��@k���3@�ʹ���!?��fX��@�2�Ԗٿ��
}���@[.�v��3@Cs�2L�!?v����@�2�Ԗٿ��
}���@[.�v��3@Cs�2L�!?v����@�2�Ԗٿ��
}���@[.�v��3@Cs�2L�!?v����@�2�Ԗٿ��
}���@[.�v��3@Cs�2L�!?v����@7�K�ٿU#�2���@�n�� 4@M-B��!?�y"��@Cƌᾘٿ|4���@��v�t 4@����!?/?���@Cƌᾘٿ|4���@��v�t 4@����!?/?���@Cƌᾘٿ|4���@��v�t 4@����!?/?���@ע�Fؘٿ�G]����@z��^o 4@���Ǐ!?�}���@ע�Fؘٿ�G]����@z��^o 4@���Ǐ!?�}���@��9�ŘٿĿ�����@4
��3@�H*bZ�!?���k��@�M�o�ٿ}"� ��@m<,�h�3@M�ku�!?㵣���@�M�o�ٿ}"� ��@m<,�h�3@M�ku�!?㵣���@�ٻ,��ٿ��" ��@qY:
��3@�_�p�!?"d����@�ٻ,��ٿ��" ��@qY:
��3@�_�p�!?"d����@�ٻ,��ٿ��" ��@qY:
��3@�_�p�!?"d����@�ٻ,��ٿ��" ��@qY:
��3@�_�p�!?"d����@}Ue9+�ٿe�7 ��@o��A&�3@i��K�!?��E���@��Q�ٿ�B�T ��@�˧�N�3@طߏ�!?,3���@��F_��ٿ��� ��@A��غ�3@���Z�!?,ސ��@��F_��ٿ��� ��@A��غ�3@���Z�!?,ސ��@��F_��ٿ��� ��@A��غ�3@���Z�!?,ސ��@��F_��ٿ��� ��@A��غ�3@���Z�!?,ސ��@��F_��ٿ��� ��@A��غ�3@���Z�!?,ސ��@=Б��ٿ�#����@H�4q��3@�=�6�!?O�c��@=Б��ٿ�#����@H�4q��3@�=�6�!?O�c��@=Б��ٿ�#����@H�4q��3@�=�6�!?O�c��@=Б��ٿ�#����@H�4q��3@�=�6�!?O�c��@Ee����ٿ�1. ��@1�F]l�3@"9�7|�!?�x�L��@�����ٿɡ�����@�!�P��3@l�9�w�!?]y[���@���zƜٿ&�����@�C�� 4@wI�h�!?S�VV��@���zƜٿ&�����@�C�� 4@wI�h�!?S�VV��@���zƜٿ&�����@�C�� 4@wI�h�!?S�VV��@���zƜٿ&�����@�C�� 4@wI�h�!?S�VV��@�_/^�ٿ��|� ��@%����3@+,Rp�!?ov���@�_/^�ٿ��|� ��@%����3@+,Rp�!?ov���@�_/^�ٿ��|� ��@%����3@+,Rp�!?ov���@G?*�G�ٿ�\����@#��t��3@�o�<|�!?��01��@G?*�G�ٿ�\����@#��t��3@�o�<|�!?��01��@�KE�ٿ�%; ��@0��,�3@�_z���!?�Rp��@�KE�ٿ�%; ��@0��,�3@�_z���!?�Rp��@�KE�ٿ�%; ��@0��,�3@�_z���!?�Rp��@�i[?�ٿ�����@��Q��3@��\�!?�?3���@�i[?�ٿ�����@��Q��3@��\�!?�?3���@���'�ٿV̞���@��l���3@�1mnP�!?:�����@���'�ٿV̞���@��l���3@�1mnP�!?:�����@���'�ٿV̞���@��l���3@�1mnP�!?:�����@���'�ٿV̞���@��l���3@�1mnP�!?:�����@�ܺT�ٿ������@t�;�? 4@�gSl��!?�j6N��@a�c�ٿ���l���@���"4@�_��w�!?�ŏ�@a�c�ٿ���l���@���"4@�_��w�!?�ŏ�@a�c�ٿ���l���@���"4@�_��w�!?�ŏ�@a�c�ٿ���l���@���"4@�_��w�!?�ŏ�@n�M���ٿwJ�����@�!��� 4@���vw�!?�����@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@r��Cr�ٿG�����@����1 4@��(C��!?R8hz��@��8��ٿh�����@񜫨� 4@c�ĚR�!?�/���@��8��ٿh�����@񜫨� 4@c�ĚR�!?�/���@�1K[�ٿ$�, ��@�-k���3@�z\�j�!?A,
j��@�1K[�ٿ$�, ��@�-k���3@�z\�j�!?A,
j��@�1K[�ٿ$�, ��@�-k���3@�z\�j�!?A,
j��@�1K[�ٿ$�, ��@�-k���3@�z\�j�!?A,
j��@�1K[�ٿ$�, ��@�-k���3@�z\�j�!?A,
j��@g�&�ٿ�������@0y����3@/j��W�!?Q�����@�r@�Әٿ�� ��@�ŋ(�3@FQFJ�!?�p����@�r@�Әٿ�� ��@�ŋ(�3@FQFJ�!?�p����@�r@�Әٿ�� ��@�ŋ(�3@FQFJ�!?�p����@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@i�{$ɛٿd,�� ��@U��O��3@2R���!?F�k���@��.KF�ٿ1�fx ��@U��l��3@9l�8�!?�h!���@�iZO��ٿ��U ��@��3�! 4@�ټ�#�!?������@�iZO��ٿ��U ��@��3�! 4@�ټ�#�!?������@_T.�ٿ��R[���@��^r4@"�,�K�!?z6W+�@_T.�ٿ��R[���@��^r4@"�,�K�!?z6W+�@_T.�ٿ��R[���@��^r4@"�,�K�!?z6W+�@/wK
�ٿ�8,���@�;��<4@�r���!?�B(�@�&ӟٿy8���@�;�;� 4@�>�F#�!?z޸@�@�&ӟٿy8���@�;�;� 4@�>�F#�!?z޸@�@�V�ۻ�ٿ���� ��@� (�Y�3@z8�;�!?�4����@�V�ۻ�ٿ���� ��@� (�Y�3@z8�;�!?�4����@��b'�ٿbq4��@2�����3@V�ykY�!?�
u<��@��b'�ٿbq4��@2�����3@V�ykY�!?�
u<��@��b'�ٿbq4��@2�����3@V�ykY�!?�
u<��@���4�ٿCX� ��@Q�Uk�3@;|V��!?G�n���@���4�ٿCX� ��@Q�Uk�3@;|V��!?G�n���@�B�ٿ�\����@ռ.| 4@{�����!?TYr��@��J��ٿ�Tdy��@���'��3@d��`�!?�r����@HU&�&�ٿ/��8��@uX	��3@|���g�!?�Rb��@HU&�&�ٿ/��8��@uX	��3@|���g�!?�Rb��@HU&�&�ٿ/��8��@uX	��3@|���g�!?�Rb��@HU&�&�ٿ/��8��@uX	��3@|���g�!?�Rb��@HU&�&�ٿ/��8��@uX	��3@|���g�!?�Rb��@�3�֝ٿ���-��@;&���3@���o�!?h*���@�}�B�ٿ�V���@b��[��3@:�+�!?�M���@�}�B�ٿ�V���@b��[��3@:�+�!?�M���@�}�B�ٿ�V���@b��[��3@:�+�!?�M���@�g�ٿK�2v��@	�Y)1�3@�m��]�!?p±S��@�g�ٿK�2v��@	�Y)1�3@�m��]�!?p±S��@����ٿ���}���@Hwb��4@�+q�w�!?�Ң7�@����ٿ���}���@Hwb��4@�+q�w�!?�Ң7�@����ٿ���}���@Hwb��4@�+q�w�!?�Ң7�@�/g���ٿU�f����@c��f4@��M���!?nb��@����o�ٿ��]���@�־�	4@��tC{�!?������@��n�U�ٿ>�m����@(f�+4@��P~�!?�!C��@h aB��ٿ�$%����@���#4@^�!Aw�!?�ݠ}�@��p��ٿt�?���@�i��A�3@�TW�o�!?UZd��@��p��ٿt�?���@�i��A�3@�TW�o�!?UZd��@��p��ٿt�?���@�i��A�3@�TW�o�!?UZd��@?��>��ٿ8�v����@ʗ-���3@��\�z�!?�X+��@|�d�
�ٿγ�����@�P��3@�"f��!?!�� �@�ry��ٿ��L����@D&H`�4@IM�|�!?��f#��@*<NRf�ٿh������@��ګ<	4@Ʃ��K�!?e�li��@*<NRf�ٿh������@��ګ<	4@Ʃ��K�!?e�li��@�JC��ٿ�o��@����E4@��5��!?x�"s�@�JC��ٿ�o��@����E4@��5��!?x�"s�@����h�ٿ<�	9���@�',g:4@g/�1�!?��ک��@����h�ٿ<�	9���@�',g:4@g/�1�!?��ک��@����h�ٿ<�	9���@�',g:4@g/�1�!?��ک��@E�-�ٿL����@f�z�d4@�{�pD�!?��Xʯ�@h�4&�ٿ���4��@�.���4@�ЂB'�!?�����@h�4&�ٿ���4��@�.���4@�ЂB'�!?�����@h�4&�ٿ���4��@�.���4@�ЂB'�!?�����@�ؼN�ٿ�ә-��@��6��4@�W�d�!?3m6x��@�ؼN�ٿ�ә-��@��6��4@�W�d�!?3m6x��@�ؼN�ٿ�ә-��@��6��4@�W�d�!?3m6x��@�ؼN�ٿ�ә-��@��6��4@�W�d�!?3m6x��@�G�g�ٿ#Tޙ���@��%Uh4@8[P�u�!?a6�
�@�G�g�ٿ#Tޙ���@��%Uh4@8[P�u�!?a6�
�@��S�0�ٿ}�6���@��z�4@�ȅ1�!?<�Q�@��S�0�ٿ}�6���@��z�4@�ȅ1�!?<�Q�@	�/�o�ٿl���@e��H4@�VG�
�!?-�u��@	�/�o�ٿl���@e��H4@�VG�
�!?-�u��@	�/�o�ٿl���@e��H4@�VG�
�!?-�u��@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@`mΔ�ٿ��>��@Kc1J4@�1�}7�!?Z�	7�@�D���ٿW+�?��@�"���4@U�Y�!?C�}w�@�D���ٿW+�?��@�"���4@U�Y�!?C�}w�@�D���ٿW+�?��@�"���4@U�Y�!?C�}w�@�D���ٿW+�?��@�"���4@U�Y�!?C�}w�@�V�۟ٿ Mk-և�@�(9ig.4@GJ����!?�!��J�@�|F)[�ٿ��S·�@�iB944@��x?�!?��È��@7xSc��ٿ6/�݇�@r)�m$4@Ș�j&�!?�"�/a�@OjL76�ٿ�Ŀ%��@�af�4@��K�Ԑ!?�`��+�@M̂��ٿ��Q�ȇ�@��x�A4@2�,А!?�t�]
�@M̂��ٿ��Q�ȇ�@��x�A4@2�,А!?�t�]
�@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@-�U9Ϡٿ��U���@kS4@(��4�!?p4O��@��I�ٿ����Ӈ�@e@�6�;4@Y$���!?���&m	�@7Y���ٿ���^���@�
�j	c4@����2�!?�����@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@��f��ٿJ�@����@"���P4@,�0�n�!?�"Np�@�)�$(�ٿ��S���@}����3@s3ZO�!?;-�@�)�$(�ٿ��S���@}����3@s3ZO�!?;-�@�)�$(�ٿ��S���@}����3@s3ZO�!?;-�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@ �7�ٿ���1��@�����4@&��ZB�!?Iu�xL�@�Ί���ٿ�-�����@}���h4@:�㆐!?��b��@�Ί���ٿ�-�����@}���h4@:�㆐!?��b��@���}�ٿ)&б���@/�MgbL4@(����!?[VF#�@���}�ٿ)&б���@/�MgbL4@(����!?[VF#�@���}�ٿ)&б���@/�MgbL4@(����!?[VF#�@���}�ٿ)&б���@/�MgbL4@(����!?[VF#�@���}�ٿ)&б���@/�MgbL4@(����!?[VF#�@<��c�ٿ����@b�p}��3@�5�]Տ!?�"�@RR�h��ٿ­����@@5^u��3@jDB���!?Ԉ
H��@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@�]>��ٿ��nd���@#+)�"�3@�ʸ���!?�8����@���!�ٿ������@�[#�b�3@�+K��!?�Ȥʳ�@�%cT�ٿ:��a��@w�m�4@c,�zU�!?&�8�P�@�%cT�ٿ:��a��@w�m�4@c,�zU�!?&�8�P�@�%cT�ٿ:��a��@w�m�4@c,�zU�!?&�8�P�@�%cT�ٿ:��a��@w�m�4@c,�zU�!?&�8�P�@�%cT�ٿ:��a��@w�m�4@c,�zU�!?&�8�P�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@+f����ٿ�e�����@#
ݱI4@�]�2��!?�w�T�
�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@�/-[[�ٿ9������@NG�d�4@��2F�!?���]�@܀����ٿ�of\���@�
ڱ4@L�[�u�!?:�4���@܀����ٿ�of\���@�
ڱ4@L�[�u�!?:�4���@܀����ٿ�of\���@�
ڱ4@L�[�u�!?:�4���@܀����ٿ�of\���@�
ڱ4@L�[�u�!?:�4���@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@\�M�o�ٿ�����@���3@6q��i�!?i~�^��@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@�57錙ٿ���؇�@�����74@�F��!?%�		�@t b��ٿ����@�x��B4@�2���!?���@t b��ٿ����@�x��B4@�2���!?���@t b��ٿ����@�x��B4@�2���!?���@t b��ٿ����@�x��B4@�2���!?���@t b��ٿ����@�x��B4@�2���!?���@pǏ�ٿ�[Q����@y�RJ<
4@���պ�!?W�T��@pǏ�ٿ�[Q����@y�RJ<
4@���պ�!?W�T��@pǏ�ٿ�[Q����@y�RJ<
4@���պ�!?W�T��@pǏ�ٿ�[Q����@y�RJ<
4@���պ�!?W�T��@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@7�7`5�ٿ�~�$��@$�@�3@ג�\M�!?A�a�@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@�w;�L�ٿ=�=��@�����3@�Ȩ�P�!?��'���@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@Mƨ=�ٿ�;'�ه�@���34@= ƭR�!?Q�;��@�����ٿ��(��@QNf���3@�����!?G���@ ��Q�ٿhN.�ˇ�@$����.4@ɜ0���!?�>P�o�@���/�ٿ֖C��@���p�3@����U�!?~k�k~�@���/�ٿ֖C��@���p�3@����U�!?~k�k~�@���/�ٿ֖C��@���p�3@����U�!?~k�k~�@���/�ٿ֖C��@���p�3@����U�!?~k�k~�@���/�ٿ֖C��@���p�3@����U�!?~k�k~�@_���ٿ�y�����@f(?4@m�󢋐!?�ϕ�6�@_���ٿ�y�����@f(?4@m�󢋐!?�ϕ�6�@���ᝡٿ��T���@�����3@��Y�^�!?eqC|k �@���ᝡٿ��T���@�����3@��Y�^�!?eqC|k �@�TЍd�ٿ|<ՙ��@ݘ�t��3@Ka��!?��b��@�TЍd�ٿ|<ՙ��@ݘ�t��3@Ka��!?��b��@�����ٿ'��2��@�U�4@qa��T�!?à>ձ�@)�N�ٿ\�%���@L����3@���l/�!?cL�5
�@����ӣٿ9�����@�ة!4@����J�!?�$�;��@)��o�ٿ��HӇ�@��/zX24@qla�p�!?��6l��@)��o�ٿ��HӇ�@��/zX24@qla�p�!?��6l��@)��o�ٿ��HӇ�@��/zX24@qla�p�!?��6l��@)��o�ٿ��HӇ�@��/zX24@qla�p�!?��6l��@)��o�ٿ��HӇ�@��/zX24@qla�p�!?��6l��@�ǣ��ٿ�(&�
��@�7{�^�3@��K�!?�.����@�h���ٿ�����@ҙ���3@`�)`�!?}`���@�h���ٿ�����@ҙ���3@`�)`�!?}`���@�h���ٿ�����@ҙ���3@`�)`�!?}`���@�h���ٿ�����@ҙ���3@`�)`�!?}`���@�h���ٿ�����@ҙ���3@`�)`�!?}`���@�h���ٿ�����@ҙ���3@`�)`�!?}`���@����֘ٿr������@Ѷ��d
4@_��0�!?~���@����֘ٿr������@Ѷ��d
4@_��0�!?~���@����֘ٿr������@Ѷ��d
4@_��0�!?~���@����֘ٿr������@Ѷ��d
4@_��0�!?~���@����֘ٿr������@Ѷ��d
4@_��0�!?~���@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@C[�ٿ�����@����
4@�W��W�!?5�����@�ȟ�ٿ�����@���1�3@�7��B�!?4�����@�ȟ�ٿ�����@���1�3@�7��B�!?4�����@�ȟ�ٿ�����@���1�3@�7��B�!?4�����@�ȟ�ٿ�����@���1�3@�7��B�!?4�����@�ȟ�ٿ�����@���1�3@�7��B�!?4�����@����h�ٿ��*[��@��\���3@�-��W�!?��a��@HI�B�ٿ4�Y��@B�Y6�3@oN�R�!?����F�@HI�B�ٿ4�Y��@B�Y6�3@oN�R�!?����F�@�%{��ٿ1B�j���@�/`Q�4@kTNM��!?�84���@�%{��ٿ1B�j���@�/`Q�4@kTNM��!?�84���@��Ù�ٿ�#����@7�l�+4@��]�!?ٜ��P�@1qҢٿ���uc��@(�2�'4@d�u[�!?Ԟ�6�@1qҢٿ���uc��@(�2�'4@d�u[�!?Ԟ�6�@1qҢٿ���uc��@(�2�'4@d�u[�!?Ԟ�6�@1qҢٿ���uc��@(�2�'4@d�u[�!?Ԟ�6�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@�]��c�ٿU9.w��@��u�<	4@�^+w�!?�CQs�@��V�աٿ��r�_��@�ӷ�I)4@�\/0�!?l��o	�@��9��ٿ�չ��@z�� !4@���	�!?,,8�x�@��9��ٿ�չ��@z�� !4@���	�!?,,8�x�@��9��ٿ�չ��@z�� !4@���	�!?,,8�x�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@�|X�Θٿ�K0d��@�;��3@�T~%�!?�(:�_�@q�N��ٿ�MU���@�%�_�3@zǁ�-�!?i�N"�@q�N��ٿ�MU���@�%�_�3@zǁ�-�!?i�N"�@q�N��ٿ�MU���@�%�_�3@zǁ�-�!?i�N"�@q�N��ٿ�MU���@�%�_�3@zǁ�-�!?i�N"�@[<�/�ٿ�S�Li��@����I�3@$�=q�!??�S� �@[<�/�ٿ�S�Li��@����I�3@$�=q�!??�S� �@[<�/�ٿ�S�Li��@����I�3@$�=q�!??�S� �@��;��ٿ�l!��@i�����3@���m�!?��HX�@�����ٿ���=���@�O`�3@jw�ˬ�!?���+= �@�����ٿ���=���@�O`�3@jw�ˬ�!?���+= �@�����ٿ���=���@�O`�3@jw�ˬ�!?���+= �@�����ٿ���=���@�O`�3@jw�ˬ�!?���+= �@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@W��P�ٿ���CЇ�@����3@�H��U�!?�TOzS�@��;:*�ٿ�L[��@�{��K�3@:����!?��Z��@��;:*�ٿ�L[��@�{��K�3@:����!?��Z��@��;:*�ٿ�L[��@�{��K�3@:����!?��Z��@�?f�ٿc�*Q���@v*φ��3@��ɧ�!? �a��@�?f�ٿc�*Q���@v*φ��3@��ɧ�!? �a��@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@R�+�^�ٿ\Wf�9��@���8�3@�Jڬ�!?��p �@j�2���ٿ !?��@�$�:a4@B�
�!?��w �@j�2���ٿ !?��@�$�:a4@B�
�!?��w �@j�2���ٿ !?��@�$�:a4@B�
�!?��w �@j�2���ٿ !?��@�$�:a4@B�
�!?��w �@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@CMh��ٿ=.S���@d�~!�3@O����!?P!Mh��@P:�As�ٿKͱ���@�)Fz�3@��h�!?������@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@ �a�ٿ��A$��@[!� �4@���If�!?V���3�@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@⃯�L�ٿ��^z���@_?F�e"4@Ǫ�l��!?|gK���@7?N��ٿ �_:��@U�L�jR4@���gv�!?��qv��@Tm�ٿ{^�8n��@�s�I�4@X����!?)����@Tm�ٿ{^�8n��@�s�I�4@X����!?)����@���A�ٿk��S��@�2��3@M����!?�f��@���A�ٿk��S��@�2��3@M����!?�f��@��4w�ٿ}:�����@��MU3&4@��׫6�!?�,�m�@��4w�ٿ}:�����@��MU3&4@��׫6�!?�,�m�@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@�ׅ�ٿPL���@+�&��j4@��h�!?n���@���V�ٿ���N��@6��{e�3@5����!?�� �T�@���V�ٿ���N��@6��{e�3@5����!?�� �T�@���V�ٿ���N��@6��{e�3@5����!?�� �T�@���V�ٿ���N��@6��{e�3@5����!?�� �T�@���V�ٿ���N��@6��{e�3@5����!?�� �T�@��X�ٿ��S؇�@}pu64@��]N�!?7<�"<�@��X�ٿ��S؇�@}pu64@��]N�!?7<�"<�@6�_5F�ٿ��7g��@N�!G"-4@WƉ�+�!?��Ѿ��@6�_5F�ٿ��7g��@N�!G"-4@WƉ�+�!?��Ѿ��@��ٿ7�6�5��@��;��3@Q��y5�!?�eǴ}�@��ٿ7�6�5��@��;��3@Q��y5�!?�eǴ}�@��ٿ7�6�5��@��;��3@Q��y5�!?�eǴ}�@��ٿ7�6�5��@��;��3@Q��y5�!?�eǴ}�@�)q��ٿA5w���@�����3@��S�G�!?-�i��@�)q��ٿA5w���@�����3@��S�G�!?-�i��@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�תY+�ٿ��p��@�����4@aHrt�!?F��^�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�2՞Мٿ�\ ���@�f�ھ4@������!?�'S�
�@�i}�9�ٿL�ཇ�@��@*�3@��>(M�!?�.<~j�@�i}�9�ٿL�ཇ�@��@*�3@��>(M�!?�.<~j�@�i}�9�ٿL�ཇ�@��@*�3@��>(M�!?�.<~j�@�i}�9�ٿL�ཇ�@��@*�3@��>(M�!?�.<~j�@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@NUz�ٿ~�z��@BezS��3@��
3�!?�����@=��}�ٿ5~�}���@�o�aZ�3@%�=	�!?u�N^C��@��ύ�ٿ?�^����@�8�&�3@tM�=�!?�,�E��@��ύ�ٿ?�^����@�8�&�3@tM�=�!?�,�E��@��ύ�ٿ?�^����@�8�&�3@tM�=�!?�,�E��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@y�i�ٿ�F9z���@=V��D4@���@,�!?�X¦��@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@IN�O�ٿH���@��S��)4@����F�!?xn�� �@�6b_��ٿ,d~hy��@9��a�4@J{��G�!?��>]�@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@��Qߘٿ�]x7w��@���$�4@-+��!?|EJ�	��@Ά*ĝٿv�w����@":�r�4@I�=�!?��r���@Ά*ĝٿv�w����@":�r�4@I�=�!?��r���@Ά*ĝٿv�w����@":�r�4@I�=�!?��r���@Bcp%��ٿ� ���@�1Wv�X4@v�r�!?Q�Y�@Bcp%��ٿ� ���@�1Wv�X4@v�r�!?Q�Y�@Bcp%��ٿ� ���@�1Wv�X4@v�r�!?Q�Y�@���0��ٿ����@N�'bi�3@,+�a1�!?Ǐ@���@���0��ٿ����@N�'bi�3@,+�a1�!?Ǐ@���@���.�ٿS�1~8��@�-�o/�3@N&܂�!?z���@���.�ٿS�1~8��@�-�o/�3@N&܂�!?z���@���.�ٿS�1~8��@�-�o/�3@N&܂�!?z���@j�I<��ٿ�T1a���@5` b_�3@��l)B�!?Gϟϊ�@j�I<��ٿ�T1a���@5` b_�3@��l)B�!?Gϟϊ�@;,� ��ٿ�V�B���@k
5�!�3@_� �.�!?����v	�@����ٿuh����@���TWF4@�m`��!?�_.^��@����ٿuh����@���TWF4@�m`��!?�_.^��@����ٿuh����@���TWF4@�m`��!?�_.^��@����ٿuh����@���TWF4@�m`��!?�_.^��@<Z�ɖٿu1��ބ�@)��h�3@L}F���!?�f�m�
�@<Z�ɖٿu1��ބ�@)��h�3@L}F���!?�f�m�
�@<Z�ɖٿu1��ބ�@)��h�3@L}F���!?�f�m�
�@���9�ٿ=�����@=S!� 4@�%��!?U>}�q�@���9�ٿ=�����@=S!� 4@�%��!?U>}�q�@�����ٿ>p �߅�@6>.�'4@h�72�!?;)�ٰ�@�F_Τٿ&��.���@*݂�4@��z�8�!?dh=���@�F_Τٿ&��.���@*݂�4@��z�8�!?dh=���@�F_Τٿ&��.���@*݂�4@��z�8�!?dh=���@�F_Τٿ&��.���@*݂�4@��z�8�!?dh=���@�F_Τٿ&��.���@*݂�4@��z�8�!?dh=���@2�z���ٿ}�eJ���@��lD��3@�4ؿ_�!?r*���@2�z���ٿ}�eJ���@��lD��3@�4ؿ_�!?r*���@2�z���ٿ}�eJ���@��lD��3@�4ؿ_�!?r*���@2�z���ٿ}�eJ���@��lD��3@�4ؿ_�!?r*���@2�z���ٿ}�eJ���@��lD��3@�4ؿ_�!?r*���@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�l�Ks�ٿ�
���@�+q�)�3@�~�f�!?g�1^��@�:\�ٿ}�)���@��G�r54@W�O��!?p	��@�:\�ٿ}�)���@��G�r54@W�O��!?p	��@�:\�ٿ}�)���@��G�r54@W�O��!?p	��@���^��ٿ�**6���@2w�/��3@a��)��!?�>2�@,J���ٿH"E����@�^%4@��?CP�!?ou�62ޖ@,J���ٿH"E����@�^%4@��?CP�!?ou�62ޖ@,J���ٿH"E����@�^%4@��?CP�!?ou�62ޖ@,J���ٿH"E����@�^%4@��?CP�!?ou�62ޖ@,J���ٿH"E����@�^%4@��?CP�!?ou�62ޖ@��/ʕ�ٿ�X���@���1�3@q�t��!?��p�Eɖ@I+:��ٿm|�$��@���?�3@P`6���!?��)(��@I+:��ٿm|�$��@���?�3@P`6���!?��)(��@I+:��ٿm|�$��@���?�3@P`6���!?��)(��@I+:��ٿm|�$��@���?�3@P`6���!?��)(��@I+:��ٿm|�$��@���?�3@P`6���!?��)(��@.��K��ٿ1��:��@�&�T�C4@�+�8k�!?�O�
���@.��K��ٿ1��:��@�&�T�C4@�+�8k�!?�O�
���@.��K��ٿ1��:��@�&�T�C4@�+�8k�!?�O�
���@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@c��T�ٿ�nv���@���Mh4@��씐!?4�;.~�@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@�|��ٿR�vW.��@0�X2,4@��F'�!?��Ux��@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@���ݛٿ�C���@pX7#��3@�����!?�(�-y�@Xˎ��ٿ1��{ٶ�@W�k�4@�Qy?M�!?�B�;��@Xˎ��ٿ1��{ٶ�@W�k�4@�Qy?M�!?�B�;��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@1�!�͚ٿkAv�6�@�Ծ�(4@�o0!�!?H�U��@����S�ٿ�z2v��@E�>�Y4@6���y�!?�[[���@����S�ٿ�z2v��@E�>�Y4@6���y�!?�[[���@����S�ٿ�z2v��@E�>�Y4@6���y�!?�[[���@����S�ٿ�z2v��@E�>�Y4@6���y�!?�[[���@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@#����ٿ��Ί���@� ���
4@Uf�&�!?�����_�@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��au�ٿ���T.��@'�"#��3@LS��!?\ ]c��@��ڒa�ٿ�+���@h�!�~�3@�@�$8�!?\GZS�@��ڒa�ٿ�+���@h�!�~�3@�@�$8�!?\GZS�@��ڒa�ٿ�+���@h�!�~�3@�@�$8�!?\GZS�@��ڒa�ٿ�+���@h�!�~�3@�@�$8�!?\GZS�@��j �ٿL�4�"��@z�Y��3@-/�f�!?A�7`�@��j �ٿL�4�"��@z�Y��3@-/�f�!?A�7`�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�AnO�ٿo�7����@�3$��3@W�}!�!?D��.�e�@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�� �ٿ~�O����@�)V�3@Y�Ԅ�!?�DQ��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�-v�՞ٿe����@dѤ��-4@�W����!?Q48��@�V�ӣٿ��nH��@)�?��3@�$%+�!?��ll�@�V�ӣٿ��nH��@)�?��3@�$%+�!?��ll�@�V�ӣٿ��nH��@)�?��3@�$%+�!?��ll�@՞R��ٿ���[��@ud��>4@f�kZ�!?`���7]�@՞R��ٿ���[��@ud��>4@f�kZ�!?`���7]�@՞R��ٿ���[��@ud��>4@f�kZ�!?`���7]�@՞R��ٿ���[��@ud��>4@f�kZ�!?`���7]�@����ٿ�������@�)��I4@V���!?�h<'�2�@��(�ٿ������@�xظo*4@�Up�d�!?�=�V��@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@p� ���ٿv�l��@��ph�4@��M1�!?��گ'�@����͝ٿ����q��@5Z�u��3@<R���!?��� �S�@����͝ٿ����q��@5Z�u��3@<R���!?��� �S�@����͝ٿ����q��@5Z�u��3@<R���!?��� �S�@>��L��ٿb�����@:�	�=4@�l��!?���B>_�@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��"��ٿf��_��@�� [�3@W�Ε�!?j�oX/ �@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@��)�ڜٿ«ƛ���@�Z}�:�3@oc�p�!?KLv�2�@&��,�ٿ	��6/�@� �e84@�N��l�!?����!��@&��,�ٿ	��6/�@� �e84@�N��l�!?����!��@&��,�ٿ	��6/�@� �e84@�N��l�!?����!��@V)��V�ٿ
m	���@b|���3@F�v��!?!��9�!�@V)��V�ٿ
m	���@b|���3@F�v��!?!��9�!�@V)��V�ٿ
m	���@b|���3@F�v��!?!��9�!�@�CJLk�ٿ���)(�@�̛�W�3@٨�n��!?w-�+W�@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@u��ܢٿ�/"��@�@y�3@�2thP�!?��-�=��@h��E�ٿN�L{��@���M�4@1����!?A��\�@h��E�ٿN�L{��@���M�4@1����!?A��\�@�-f�Ǘٿ%�-:���@mw0�4@���!?��\���@x���z�ٿ�M!���@}��lQ,4@��-[�!?��U�֕@x���z�ٿ�M!���@}��lQ,4@��-[�!?��U�֕@x���z�ٿ�M!���@}��lQ,4@��-[�!?��U�֕@x���z�ٿ�M!���@}��lQ,4@��-[�!?��U�֕@x���z�ٿ�M!���@}��lQ,4@��-[�!?��U�֕@�ru[�ٿf8�����@���x#4@��? �!?�30b��@�ru[�ٿf8�����@���x#4@��? �!?�30b��@�ru[�ٿf8�����@���x#4@��? �!?�30b��@�ru[�ٿf8�����@���x#4@��? �!?�30b��@�ru[�ٿf8�����@���x#4@��? �!?�30b��@�ru[�ٿf8�����@���x#4@��? �!?�30b��@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@Z`ؠ�ٿ�@�?���@I)��#4@��L�9�!?�j���@B�şٿf�X��@.�V��3@�J�;�!?޳�éȕ@B�şٿf�X��@.�V��3@�J�;�!?޳�éȕ@��'<��ٿ�����@b��(��3@�!���!? ��/r��@��'<��ٿ�����@b��(��3@�!���!? ��/r��@��'<��ٿ�����@b��(��3@�!���!? ��/r��@O���ٿ��'!��@����3@G~�ת�!?�Jiq�@O���ٿ��'!��@����3@G~�ת�!?�Jiq�@O���ٿ��'!��@����3@G~�ת�!?�Jiq�@O���ٿ��'!��@����3@G~�ת�!?�Jiq�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@O
����ٿ{6K��@J>�I�3@��Ȁ�!?�6��0�@�D\��ٿw�-����@8UC8��3@���Z|�!?,����3�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@��{��ٿ�M���@�
��'�3@v�ͻ�!?���3K�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@NC�\��ٿR"����@��Tf�3@��ci�!?y���?	�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@�A��ٿ(����@
�	`k�3@亚>��!?�{�B�=�@����ٿ�c8_B��@�����3@����!?��k��F�@����ٿ�c8_B��@�����3@����!?��k��F�@�x�ٿ2t��1�@rF�w�4@B�D^�!?���
o��@�x�ٿ2t��1�@rF�w�4@B�D^�!?���
o��@�x�ٿ2t��1�@rF�w�4@B�D^�!?���
o��@�x�ٿ2t��1�@rF�w�4@B�D^�!?���
o��@�x�ٿ2t��1�@rF�w�4@B�D^�!?���
o��@�%�g��ٿaZ/���@Ju��4@m~bP��!?�n��8C�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@hxkŜٿKb�v�@��=*�4@� J9�!?���Ĥ�@���L)�ٿT��>j��@ohj�5�3@>�G>G�!?_ŝ׽2�@���L)�ٿT��>j��@ohj�5�3@>�G>G�!?_ŝ׽2�@���L)�ٿT��>j��@ohj�5�3@>�G>G�!?_ŝ׽2�@���L)�ٿT��>j��@ohj�5�3@>�G>G�!?_ŝ׽2�@���L)�ٿT��>j��@ohj�5�3@>�G>G�!?_ŝ׽2�@:���b�ٿ$�[����@ǚ�)O4@��y��!?(o�֕@�^9i��ٿ��Y����@^��(I
4@
N��!?��b��@�^9i��ٿ��Y����@^��(I
4@
N��!?��b��@�^9i��ٿ��Y����@^��(I
4@
N��!?��b��@U��{�ٿ�(;���@��-4@�X�M�!?_��G�V�@U��{�ٿ�(;���@��-4@�X�M�!?_��G�V�@U��{�ٿ�(;���@��-4@�X�M�!?_��G�V�@U��{�ٿ�(;���@��-4@�X�M�!?_��G�V�@U��{�ٿ�(;���@��-4@�X�M�!?_��G�V�@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@�2|�q�ٿ�@w����@պ|�?4@��
�n�!?rh�J���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@d�=2�ٿ!/&����@���g4@9�Fb*�!?^��U���@�Wۜٿ�f�����@�v�9/4@˅�=�!?]%����@*j�\[�ٿF��̉��@�k�g4@K�����!?j���^ؕ@s5��ģٿ�+>��@l#���4@���>]�!?���D��@s5��ģٿ�+>��@l#���4@���>]�!?���D��@s5��ģٿ�+>��@l#���4@���>]�!?���D��@s5��ģٿ�+>��@l#���4@���>]�!?���D��@���ă�ٿ|1b���@��LD$4@����9�!?�x%b��@���ă�ٿ|1b���@��LD$4@����9�!?�x%b��@b��ٖٿS�/r��@}�&z�3@�m>Ԉ�!?t^��S�@b��ٖٿS�/r��@}�&z�3@�m>Ԉ�!?t^��S�@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@���G�ٿ��$���@nA�5&�3@���`�!?�w�땕@<aw-[�ٿ͑p����@HG�!4@���_�!?\�'w:�@<aw-[�ٿ͑p����@HG�!4@���_�!?\�'w:�@<aw-[�ٿ͑p����@HG�!4@���_�!?\�'w:�@�!Q!�ٿZ,����@vG�p��3@��/%�!?�������@�!Q!�ٿZ,����@vG�p��3@��/%�!?�������@�!Q!�ٿZ,����@vG�p��3@��/%�!?�������@�!Q!�ٿZ,����@vG�p��3@��/%�!?�������@a��ޜٿM�B����@*�;���3@�:���!?�Ѓ�s��@a��ޜٿM�B����@*�;���3@�:���!?�Ѓ�s��@�c��	�ٿM�%��@�g:C��3@�J�:�!?�����@�c��	�ٿM�%��@�g:C��3@�J�:�!?�����@�c��	�ٿM�%��@�g:C��3@�J�:�!?�����@Dή�-�ٿ�L(>��@�٪�\�3@�TlW�!?�˵^�@Dή�-�ٿ�L(>��@�٪�\�3@�TlW�!?�˵^�@Dή�-�ٿ�L(>��@�٪�\�3@�TlW�!?�˵^�@Dή�-�ٿ�L(>��@�٪�\�3@�TlW�!?�˵^�@Dή�-�ٿ�L(>��@�٪�\�3@�TlW�!?�˵^�@F�}�ڝٿ�U����@��vc)4@���;�!?�zw%2�@F�}�ڝٿ�U����@��vc)4@���;�!?�zw%2�@F�}�ڝٿ�U����@��vc)4@���;�!?�zw%2�@F�}�ڝٿ�U����@��vc)4@���;�!?�zw%2�@F�}�ڝٿ�U����@��vc)4@���;�!?�zw%2�@��a��ٿ�2S׈��@�ٿ)�(4@=���.�!?ʙ��{��@��a��ٿ�2S׈��@�ٿ)�(4@=���.�!?ʙ��{��@��a��ٿ�2S׈��@�ٿ)�(4@=���.�!?ʙ��{��@��a��ٿ�2S׈��@�ٿ)�(4@=���.�!?ʙ��{��@Wk�-%�ٿh�U�)�@|~3�4@�Fr��!?Y���@Wk�-%�ٿh�U�)�@|~3�4@�Fr��!?Y���@Wk�-%�ٿh�U�)�@|~3�4@�Fr��!?Y���@Wk�-%�ٿh�U�)�@|~3�4@�Fr��!?Y���@g�5\��ٿ���N#��@ts+��3@��f��!?4�]�^Ε@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@e��)�ٿ��`��@���t�4@a@��O�!?>������@c"kO�ٿ����ˑ�@�q,�%�3@�CP7Q�!?� x�A��@�ܤ��ٿ�w���%�@�#ue�3@Ռn�,�!?,����@N���Ҡٿ���s���@����3@��
8�!?b:�b�@N���Ҡٿ���s���@����3@��
8�!?b:�b�@N���Ҡٿ���s���@����3@��
8�!?b:�b�@۽�G��ٿ�r�
 ��@�E}�U�3@����!�!?V�	e�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@|�Y�ҞٿL�w��b�@�b5� 4@p1�1�!?�?O_�@�b�� �ٿ��i�E(�@q�Q�4@���x�!?�Jn�S��@�b�� �ٿ��i�E(�@q�Q�4@���x�!?�Jn�S��@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���M�ٿ���QN�@ֈ�'�3@a��k�!?�c�5]ϕ@���lC�ٿr��ϲ!�@ݪp�4@�H��;�!?�Z��ѥ�@&���ǜٿ��~y�v�@��7�3@�\�Ɛ!?��BV��@3��ԝٿ(�:J�'�@�95UF�3@+�K�!?	RIf�@3��ԝٿ(�:J�'�@�95UF�3@+�K�!?	RIf�@3��ԝٿ(�:J�'�@�95UF�3@+�K�!?	RIf�@3��ԝٿ(�:J�'�@�95UF�3@+�K�!?	RIf�@�g��ٿ�Kbk���@��`'4@���D��!?���e�ԕ@�g��ٿ�Kbk���@��`'4@���D��!?���e�ԕ@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@��^W՚ٿ.��I��@��%
�&4@.a�B�!?�1�*��@�[C氠ٿ(�uN��@ߒ�w�4@���S�!?�A�-�V�@�� �ٿz1�^��@ �\D4@i��?#�!?�u�Hޕ@[���¤ٿKsQa�@�W�ԛ�3@�-g�N�!?�̐	J-�@j'�ˮ�ٿ~�Ԡ�2�@c3��V4@N��7/�!?�+���@��Rܠٿ�Ɏ��@s��Gr:4@�
yM8�!?�P��?�@�L��Ңٿp�.���@�F)C<�3@3���\�!?��=ڸ��@�L��Ңٿp�.���@�F)C<�3@3���\�!?��=ڸ��@�L��Ңٿp�.���@�F)C<�3@3���\�!?��=ڸ��@��U���ٿr��O-�@1Ph/4@LX	�!?09�w��@��U���ٿr��O-�@1Ph/4@LX	�!?09�w��@��U���ٿr��O-�@1Ph/4@LX	�!?09�w��@��U���ٿr��O-�@1Ph/4@LX	�!?09�w��@��U���ٿr��O-�@1Ph/4@LX	�!?09�w��@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@4'Mp�ٿ����^�@�/YL�4@*
�N�!?��s�@�V�F �ٿ	������@;T�.4@�L��|�!?W�2d�̕@�V�F �ٿ	������@;T�.4@�L��|�!?W�2d�̕@�V�F �ٿ	������@;T�.4@�L��|�!?W�2d�̕@�V�F �ٿ	������@;T�.4@�L��|�!?W�2d�̕@�V�F �ٿ	������@;T�.4@�L��|�!?W�2d�̕@�ށ�֜ٿ�%��%��@��=���3@PLO�!?��Gc�@�ށ�֜ٿ�%��%��@��=���3@PLO�!?��Gc�@��=��ٿR$聶�@��
�[
4@IR&�!?I�]��Е@q���áٿ9����@�R�1�3@|f��W�!?�+d4�͕@q���áٿ9����@�R�1�3@|f��W�!?�+d4�͕@q���áٿ9����@�R�1�3@|f��W�!?�+d4�͕@q���áٿ9����@�R�1�3@|f��W�!?�+d4�͕@q���áٿ9����@�R�1�3@|f��W�!?�+d4�͕@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@!a�/u�ٿ��\� �@Y��6��3@{'^Ȑ!?��*r��@������ٿ�8��o��@�S_��3@��[�!?�I��p�@������ٿ�8��o��@�S_��3@��[�!?�I��p�@������ٿ�8��o��@�S_��3@��[�!?�I��p�@������ٿ�8��o��@�S_��3@��[�!?�I��p�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@>`�:��ٿ�u�E��@�OLm��3@�8ũt�!?���n�@����ٿD�k|��@��I@�3@��4L-�!?y�z�E�@����ٿD�k|��@��I@�3@��4L-�!?y�z�E�@����ٿD�k|��@��I@�3@��4L-�!?y�z�E�@^s�q��ٿ?
 0�5�@>��34@^���.�!?���z	'�@^s�q��ٿ?
 0�5�@>��34@^���.�!?���z	'�@^s�q��ٿ?
 0�5�@>��34@^���.�!?���z	'�@&��u�ٿ��O��@-\��?4@�R��K�!?��@���@&��u�ٿ��O��@-\��?4@�R��K�!?��@���@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@׷��٘ٿ���=v:�@(9���4@�.ᤐ!?��P5O�@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@7���ʖٿ��`�Q�@�g���3@�V�!?��+Õ@��먟�ٿSN��`��@���Z�	4@��P�U�!?�yy�C�@��먟�ٿSN��`��@���Z�	4@��P�U�!?�yy�C�@��@E4�ٿ��Y�@�O��_4@b�6�I�!?n�gY&��@��@E4�ٿ��Y�@�O��_4@b�6�I�!?n�gY&��@��@E4�ٿ��Y�@�O��_4@b�6�I�!?n�gY&��@��N�ٿ������@��,c4@����!?U�0����@����ٿ�Ka���@���&en4@@Q0�ݏ!?5�C F�@����ٿ�Ka���@���&en4@@Q0�ݏ!?5�C F�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@J
�DV�ٿ�����@�r���3@b��B�!?:��=�2�@�cA�ܖٿs�K�v��@�(��lT4@���?�!?�m��
�@�cA�ܖٿs�K�v��@�(��lT4@���?�!?�m��
�@�cA�ܖٿs�K�v��@�(��lT4@���?�!?�m��
�@�cA�ܖٿs�K�v��@�(��lT4@���?�!?�m��
�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@@H��ٿl4�']�@�p�e4@������!?H� CV}�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�@�#ݙٿ��4��@_���<a4@��~S�!?�.?,E�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@�կ�ٿ@�"��@�[[��24@�Ad�N�!?P��s�@�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@���՟ٿpG3 5��@�1ɭ4@?�>@�!?4m�a�@��h�қٿ��:��@�5e:�24@�˭�4�!?_�+�і@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@C\�()�ٿ��� �4�@`p�zi4@rړU�!?��$[�p�@񤦂A�ٿ8�C�@����14@��:D�!?�0]�_��@񤦂A�ٿ8�C�@����14@��:D�!?�0]�_��@񤦂A�ٿ8�C�@����14@��:D�!?�0]�_��@񤦂A�ٿ8�C�@����14@��:D�!?�0]�_��@񤦂A�ٿ8�C�@����14@��:D�!?�0]�_��@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@�7��ٿz7�\�@K4 g4@>�#.�!?+�D�d�@��?̖�ٿM��A��@�rY�4@~�dԏ!?1���i8�@��?̖�ٿM��A��@�rY�4@~�dԏ!?1���i8�@lzz"D�ٿ�{f���@���4@m��:Ə!?ДHq*�@lzz"D�ٿ�{f���@���4@m��:Ə!?ДHq*�@>|P׶�ٿꥦ5I&�@��⍠$4@� ��!?���9�ە@>|P׶�ٿꥦ5I&�@��⍠$4@� ��!?���9�ە@>|P׶�ٿꥦ5I&�@��⍠$4@� ��!?���9�ە@nC�1�ٿ��F��@�/v��3@�z#s�!?�w��Q�@nC�1�ٿ��F��@�/v��3@�z#s�!?�w��Q�@nC�1�ٿ��F��@�/v��3@�z#s�!?�w��Q�@nC�1�ٿ��F��@�/v��3@�z#s�!?�w��Q�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@U���a�ٿ���8�c�@kdO��,4@�^�EN�!?�ԮJ�L�@���b�ٿ�F�֙�@�i:�3@�4w�:�!?H�q�?��@���b�ٿ�F�֙�@�i:�3@�4w�:�!?H�q�?��@���b�ٿ�F�֙�@�i:�3@�4w�:�!?H�q�?��@���b�ٿ�F�֙�@�i:�3@�4w�:�!?H�q�?��@����;�ٿlF5LҰ�@����'4@<^·��!?{�_�Qו@����;�ٿlF5LҰ�@����'4@<^·��!?{�_�Qו@����;�ٿlF5LҰ�@����'4@<^·��!?{�_�Qו@����;�ٿlF5LҰ�@����'4@<^·��!?{�_�Qו@����;�ٿlF5LҰ�@����'4@<^·��!?{�_�Qו@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@O�mٿ)��f!c�@!�p��H4@=�+�!?���hF�@��})��ٿS��j9#�@�
���4@O� ���!?�A�7��@��})��ٿS��j9#�@�
���4@O� ���!?�A�7��@��})��ٿS��j9#�@�
���4@O� ���!?�A�7��@��})��ٿS��j9#�@�
���4@O� ���!?�A�7��@��})��ٿS��j9#�@�
���4@O� ���!?�A�7��@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@���F��ٿ�U;�@[YJ�04@e~H�6�!?^��F�@�kn�'�ٿ�an�r�@(#`��4@'�HKp�!?t�AS�_�@�kn�'�ٿ�an�r�@(#`��4@'�HKp�!?t�AS�_�@�kn�'�ٿ�an�r�@(#`��4@'�HKp�!?t�AS�_�@�kn�'�ٿ�an�r�@(#`��4@'�HKp�!?t�AS�_�@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@�6)cƛٿ�a�f�9�@!�J�3@N�F��!?̖�M��@���N��ٿ��89�@r��Y14@h�
3�!?p�tHf�@���N��ٿ��89�@r��Y14@h�
3�!?p�tHf�@�ڸ��ٿl���N.�@y��<"M4@-���<�!?pV�^�@�ڸ��ٿl���N.�@y��<"M4@-���<�!?pV�^�@�ڸ��ٿl���N.�@y��<"M4@-���<�!?pV�^�@�ڸ��ٿl���N.�@y��<"M4@-���<�!?pV�^�@�ڸ��ٿl���N.�@y��<"M4@-���<�!?pV�^�@�5�:��ٿ�0M��@�P*;I4@�eb��!?�¶.F�@�5�:��ٿ�0M��@�P*;I4@�eb��!?�¶.F�@�5�:��ٿ�0M��@�P*;I4@�eb��!?�¶.F�@�5�:��ٿ�0M��@�P*;I4@�eb��!?�¶.F�@N�,)�ٿ�vň�@JҚ�W�3@B�%\�!?@$�K@N�,)�ٿ�vň�@JҚ�W�3@B�%\�!?@$�K@i�</��ٿ�"�u��@C�-�v�3@/���!?�7���*�@ʑ�:��ٿ�/Me���@(h0-�3@�H�A!�!?�+[�ӕ@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@�v��ٿ(n?}�@5W���4@�P�Y��!?\�g�O�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@��큝ٿ��@��@+�9p��3@�]�"|�!?ᷕ�9�@%�"��ٿ�.m�05�@]�44@'��3�!?�>�	�.�@%�"��ٿ�.m�05�@]�44@'��3�!?�>�	�.�@%�"��ٿ�.m�05�@]�44@'��3�!?�>�	�.�@�O���ٿ��1���@W�(x#4@��|*N�!?� ��X�@�O���ٿ��1���@W�(x#4@��|*N�!?� ��X�@�O���ٿ��1���@W�(x#4@��|*N�!?� ��X�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@Z���8�ٿ���Zw�@W#�A4@�KYW�!?;<�9J.�@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�M݂�ٿU6w��@���ñ4@�g*U�!?A.����@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@�Sz��ٿQhIu��@�l�P�)4@F��PR�!?����g�@���2��ٿGQ�^�@ƀ�_.4@D���&�!?y80�ڕ@���2��ٿGQ�^�@ƀ�_.4@D���&�!?y80�ڕ@���2��ٿGQ�^�@ƀ�_.4@D���&�!?y80�ڕ@z;�I��ٿ�����@"��a4@��~X�!?�T>�@z;�I��ٿ�����@"��a4@��~X�!?�T>�@z;�I��ٿ�����@"��a4@��~X�!?�T>�@z;�I��ٿ�����@"��a4@��~X�!?�T>�@z;�I��ٿ�����@"��a4@��~X�!?�T>�@�}|��ٿ��l���@0�f���3@g�
,��!?�u$l��@ѻ�>��ٿ�o�U���@&��B%4@�P�u�!?I�ҕ@ѻ�>��ٿ�o�U���@&��B%4@�P�u�!?I�ҕ@ѻ�>��ٿ�o�U���@&��B%4@�P�u�!?I�ҕ@ѻ�>��ٿ�o�U���@&��B%4@�P�u�!?I�ҕ@�9���ٿ%B����@����3@��X�!?~%]��3�@�9���ٿ%B����@����3@��X�!?~%]��3�@�9���ٿ%B����@����3@��X�!?~%]��3�@�a�?�ٿzL9]��@ v	4@��?��!?J3P��ŕ@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�fѰ��ٿzt+[��@�'[��4@[.��!?,��g�T�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@�6Y�Ĝٿ�^+���@]e�H!4@��Sf�!?(_�5�\�@-2�3�ٿ.i%�S&�@�U��U�3@��&1��!?�#'ONP�@-2�3�ٿ.i%�S&�@�U��U�3@��&1��!?�#'ONP�@-2�3�ٿ.i%�S&�@�U��U�3@��&1��!?�#'ONP�@Tw�y�ٿCW�ǿ�@�X K*4@@}q�g�!?7B�g2,�@Tw�y�ٿCW�ǿ�@�X K*4@@}q�g�!?7B�g2,�@Tw�y�ٿCW�ǿ�@�X K*4@@}q�g�!?7B�g2,�@Tw�y�ٿCW�ǿ�@�X K*4@@}q�g�!?7B�g2,�@Tw�y�ٿCW�ǿ�@�X K*4@@}q�g�!?7B�g2,�@�5q&)�ٿ�"���	�@���\^4@��ue�!?m���f�@���-�ٿ��D��V�@nK?4@{�l�!?�Ԋ�k��@���-�ٿ��D��V�@nK?4@{�l�!?�Ԋ�k��@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@��(#��ٿzJʴD��@�s0j4@�*-�i�!?3���T�@�1��0�ٿ$͏C�z�@?:_<p'4@���Tu�!?a�[%O�@�1��0�ٿ$͏C�z�@?:_<p'4@���Tu�!?a�[%O�@�1��0�ٿ$͏C�z�@?:_<p'4@���Tu�!?a�[%O�@�1��0�ٿ$͏C�z�@?:_<p'4@���Tu�!?a�[%O�@6/�+u�ٿ�y`n� �@n�v��H4@���4��!?3�_@ �@6/�+u�ٿ�y`n� �@n�v��H4@���4��!?3�_@ �@m�ǟٿ��ص��@3u3��4@���J�!?b�V� �@m�ǟٿ��ص��@3u3��4@���J�!?b�V� �@2Mev#�ٿ������@iF�O�3@�~�}�!?�W�7eٕ@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@�q4?�ٿ�h�+7d�@�'i{`�3@��ˍO�!?4�\k���@���2�ٿ���A�@3&g�k14@��^�q�!?��T�!�@���2�ٿ���A�@3&g�k14@��^�q�!?��T�!�@���2�ٿ���A�@3&g�k14@��^�q�!?��T�!�@���2�ٿ���A�@3&g�k14@��^�q�!?��T�!�@���2�ٿ���A�@3&g�k14@��^�q�!?��T�!�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@/�e�a�ٿ� �
=%�@�I���H4@4CHP�!?�dA�4(�@2H�ۅ�ٿ�o�c�@���ڜ�3@�DD�P�!?'K�:��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@k�� ^�ٿ�")jp�@�k֌�3@��u_G�!?"d5ޱ��@��b��ٿ�|���&�@�5ş4@��	|��!?�(����@��b��ٿ�|���&�@�5ş4@��	|��!?�(����@��b��ٿ�|���&�@�5ş4@��	|��!?�(����@��b��ٿ�|���&�@�5ş4@��	|��!?�(����@0�#���ٿ�Mح���@�W��j�3@�2q���!?σ�c�Օ@���j��ٿ١���@[<�R)�3@�b����!?�-=�@Q���;�ٿgXK-��@��"E<4@m�Q�j�!??⤀#�@Q���;�ٿgXK-��@��"E<4@m�Q�j�!??⤀#�@Q���;�ٿgXK-��@��"E<4@m�Q�j�!??⤀#�@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@P^���ٿ�\U6'��@��m14@�M~�!?�Hs4 �@�����ٿ8��[ߙ�@��"4@"�*�e�!?�0F31?�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@l��%�ٿ�zh����@x� �4@�j�pq�!?��)�@�@��e	�ٿ��l��p�@�u{�3@����l�!?_�y�C2�@��e	�ٿ��l��p�@�u{�3@����l�!?_�y�C2�@�\�f%�ٿ>�{���@�R0d�
4@q��v.�!?��s��@�\�f%�ٿ>�{���@�R0d�
4@q��v.�!?��s��@q-�͞ٿ�/c��7�@�7g1�3@�t��+�!?���0r_�@q-�͞ٿ�/c��7�@�7g1�3@�t��+�!?���0r_�@d���ٿ�h��w�@�����3@�]-�v�!?6��|�@d���ٿ�h��w�@�����3@�]-�v�!?6��|�@d���ٿ�h��w�@�����3@�]-�v�!?6��|�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@r�ov��ٿC:>~V(�@O �+�3@�H��q�!?u�[�@yh����ٿL��/���@���]�3@�qz�!?)����@yh����ٿL��/���@���]�3@�qz�!?)����@yh����ٿL��/���@���]�3@�qz�!?)����@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@rr��!�ٿ�)���@���*�%4@�`!�,�!?���|��@�F���ٿ�8f����@�7h�#4@����x�!?%�o|��@�F���ٿ�8f����@�7h�#4@����x�!?%�o|��@�F���ٿ�8f����@�7h�#4@����x�!?%�o|��@�F���ٿ�8f����@�7h�#4@����x�!?%�o|��@�F���ٿ�8f����@�7h�#4@����x�!?%�o|��@TD�~�ٿ"�<��+�@&�K4@���g�!?h��ҕ@TD�~�ٿ"�<��+�@&�K4@���g�!?h��ҕ@�7tň�ٿ�9�u�5�@���{�,4@c?�a1�!?�ő[�8�@�7tň�ٿ�9�u�5�@���{�,4@c?�a1�!?�ő[�8�@�7tň�ٿ�9�u�5�@���{�,4@c?�a1�!?�ő[�8�@�7tň�ٿ�9�u�5�@���{�,4@c?�a1�!?�ő[�8�@��+@�ٿ�!k�b�@O��44@*��4�!?z�>����@��+@�ٿ�!k�b�@O��44@*��4�!?z�>����@��+@�ٿ�!k�b�@O��44@*��4�!?z�>����@�׶]��ٿ�I����@�Hf�=4@��+���!?�w7���@�Y���ٿ�����\�@�>�ju4@P�< �!?R?�e�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@HL =>�ٿ����~�@]�b|^4@�8��!?���P�v�@�r�z)�ٿ��'�kR�@�?L�h?4@)8��N�!?�[��^q�@�r�z)�ٿ��'�kR�@�?L�h?4@)8��N�!?�[��^q�@�r�z)�ٿ��'�kR�@�?L�h?4@)8��N�!?�[��^q�@�r�z)�ٿ��'�kR�@�?L�h?4@)8��N�!?�[��^q�@X��*M�ٿ�0ƈ7�@��R�4@8�V�!?x�_�@���ֳ�ٿ�x�v�@��c^4�3@+����!?���W�@���ֳ�ٿ�x�v�@��c^4�3@+����!?���W�@���ֳ�ٿ�x�v�@��c^4�3@+����!?���W�@���ֳ�ٿ�x�v�@��c^4�3@+����!?���W�@���:�ٿ�p%q��@�o\Y�3@������!?�j����@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@�~~d�ٿ?��!��@��3�&4@n�\k\�!?���
�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@ʻ�r7�ٿf_1Q��@{R���3@{��X�!?��|�S�@�AXT'�ٿ�~3T_��@�֮��4@$Q�n�!?�3r����@�AXT'�ٿ�~3T_��@�֮��4@$Q�n�!?�3r����@�AXT'�ٿ�~3T_��@�֮��4@$Q�n�!?�3r����@�AXT'�ٿ�~3T_��@�֮��4@$Q�n�!?�3r����@�AXT'�ٿ�~3T_��@�֮��4@$Q�n�!?�3r����@vc�Vc�ٿqvґg��@�!�Q!4@�&h��!?]����@vc�Vc�ٿqvґg��@�!�Q!4@�&h��!?]����@vc�Vc�ٿqvґg��@�!�Q!4@�&h��!?]����@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@��m�l�ٿ�M�f��@�D��64@zd^��!?]��7���@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@�eӅj�ٿ��	�cJ�@�M���
4@�f��z�!?��^�7ĕ@{�8F��ٿ����y�@����4@��q�f�!?��}��@{�8F��ٿ����y�@����4@��q�f�!?��}��@{�8F��ٿ����y�@����4@��q�f�!?��}��@{�8F��ٿ����y�@����4@��q�f�!?��}��@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@lmQ	Y�ٿ���M��@of:֫.4@iA�Y�!?����8�@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�����ٿ>==3mI�@��@v4@���C��!?�[g��ӕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�1��ٿH=�9���@e�#�h4@ }I��!?>kRJҕ@�����ٿ�����@�7�m24@K�ޥ�!?+��r�@����ٿ1>v���@"�^���3@���q�!?pY��T�@����ٿ1>v���@"�^���3@���q�!?pY��T�@����ٿ1>v���@"�^���3@���q�!?pY��T�@��kx�ٿ��r���@*9�	�3@��?'�!?"w��@��kx�ٿ��r���@*9�	�3@��?'�!?"w��@��kx�ٿ��r���@*9�	�3@��?'�!?"w��@��kx�ٿ��r���@*9�	�3@��?'�!?"w��@cHg�ٿv�eڪ\�@�&Df�3@8n9z��!?/�x��-�@cHg�ٿv�eڪ\�@�&Df�3@8n9z��!?/�x��-�@cHg�ٿv�eڪ\�@�&Df�3@8n9z��!?/�x��-�@cHg�ٿv�eڪ\�@�&Df�3@8n9z��!?/�x��-�@m���L�ٿN������@߈���3@�=���!?��u/ܕ@������ٿ��ӿF �@+=�4@Ң�o��!?*�E��@������ٿ��ӿF �@+=�4@Ң�o��!?*�E��@������ٿ��ӿF �@+=�4@Ң�o��!?*�E��@������ٿ��ӿF �@+=�4@Ң�o��!?*�E��@������ٿ��ӿF �@+=�4@Ң�o��!?*�E��@� �c��ٿ�(�
O�@�5ogP4@{a�2��!?���S���@��.�L�ٿ��|� �@�/LK�N4@O����!?f�i���@��.�L�ٿ��|� �@�/LK�N4@O����!?f�i���@����ٿ!(z���@S^J��3@��6�w�!?mSk�˕@����ٿ!(z���@S^J��3@��6�w�!?mSk�˕@����ٿ!(z���@S^J��3@��6�w�!?mSk�˕@����ٿ!(z���@S^J��3@��6�w�!?mSk�˕@��6�Ǣٿ_n��5��@�|���44@D
>��!?��y@�@��6�Ǣٿ_n��5��@�|���44@D
>��!?��y@�@!�uA:�ٿ1��nj��@9ZK�Lm4@3{�0[�!?�̕(���@!�uA:�ٿ1��nj��@9ZK�Lm4@3{�0[�!?�̕(���@!�uA:�ٿ1��nj��@9ZK�Lm4@3{�0[�!?�̕(���@O�e��ٿ��W�v��@0���P4@�8���!?�RϊY�@O�e��ٿ��W�v��@0���P4@�8���!?�RϊY�@O�e��ٿ��W�v��@0���P4@�8���!?�RϊY�@_�I�ٿ���_9�@�`� �3@-IJ}�!? .!Φ�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@U��_ʛٿq�����@� ���3@'˜�M�!?�����f�@���d�ٿ�P��7�@��;�4@ǀRf$�!?T��-駕@���d�ٿ�P��7�@��;�4@ǀRf$�!?T��-駕@���d�ٿ�P��7�@��;�4@ǀRf$�!?T��-駕@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@�z��m�ٿx8�W�@�f�a4@���N�!?�K*�`�@m��c�ٿ���2��@._Zx'4@U��a"�!?���eו@m��c�ٿ���2��@._Zx'4@U��a"�!?���eו@m��c�ٿ���2��@._Zx'4@U��a"�!?���eו@�(�3ؔٿk�<P�@&����3@ehP(P�!?�x_k�@��p|�ٿ"��2hG�@��Q�~ 4@:tL�Ɛ!?XB��k�@�&��ٿF2J��@��-��3@D �1��!?��ц��@�&��ٿF2J��@��-��3@D �1��!?��ц��@�&��ٿF2J��@��-��3@D �1��!?��ц��@�&��ٿF2J��@��-��3@D �1��!?��ц��@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�M���ٿ�[�X<�@����;4@����!?�n���@�
�*ʜٿ��vs��@c����4@�x��]�!?\A^V1͕@3���?�ٿJ�/����@�]R�/4@wN7�@�!?%4"m��@3���?�ٿJ�/����@�]R�/4@wN7�@�!?%4"m��@3���?�ٿJ�/����@�]R�/4@wN7�@�!?%4"m��@3���?�ٿJ�/����@�]R�/4@wN7�@�!?%4"m��@��PR�ٿ�y[�u��@��CiB4@�xF=%�!?�]�
�@`<��ٿ.���r��@�:�4@�R)���!?HЬQG��@`<��ٿ.���r��@�:�4@�R)���!?HЬQG��@`<��ٿ.���r��@�:�4@�R)���!?HЬQG��@0P7��ٿpT9�cx�@����nF4@H�E�T�!?އ�Õ@0P7��ٿpT9�cx�@����nF4@H�E�T�!?އ�Õ@0P7��ٿpT9�cx�@����nF4@H�E�T�!?އ�Õ@�+�u�ٿ���Z@�@Ys/h4@��C8b�!?�'�ۓl�@�+�u�ٿ���Z@�@Ys/h4@��C8b�!?�'�ۓl�@�+�u�ٿ���Z@�@Ys/h4@��C8b�!?�'�ۓl�@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@P��+��ٿ��\h��@qQN4@��ݦ��!?�����@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@_ã8�ٿx��N ��@�*.4@;��B^�!?jL;lR�@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@ ��ٿyx@���@����64@�9�B\�!?k����@2}��Ǡٿ�<V��7�@�r6�4@ ���!?�|:���@�ux�ٿb���5�@+���D4@��t�!?B����@�]Kq�ٿ�ʭ!�"�@��'*��3@��_���!?���@�]Kq�ٿ�ʭ!�"�@��'*��3@��_���!?���@�]Kq�ٿ�ʭ!�"�@��'*��3@��_���!?���@�]Kq�ٿ�ʭ!�"�@��'*��3@��_���!?���@�]Kq�ٿ�ʭ!�"�@��'*��3@��_���!?���@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�dK��ٿF@@���@�K�1v	4@%�G\�!?�Z����@�n5�X�ٿ�F��C�@������3@4�+���!?��o�-�@���1�ٿ��z]��@��I�5�3@��Y�c�!?G��q���@���1�ٿ��z]��@��I�5�3@��Y�c�!?G��q���@���1�ٿ��z]��@��I�5�3@��Y�c�!?G��q���@�WM�{�ٿU�3���@ts�)(4@�8(8�!?s[E��@�WM�{�ٿU�3���@ts�)(4@�8(8�!?s[E��@�WM�{�ٿU�3���@ts�)(4@�8(8�!?s[E��@�WM�{�ٿU�3���@ts�)(4@�8(8�!?s[E��@�@��?�ٿ���"(�@IU�Z34@{���%�!?;/��Õ@�@��?�ٿ���"(�@IU�Z34@{���%�!?;/��Õ@�@��?�ٿ���"(�@IU�Z34@{���%�!?;/��Õ@/��ʹ�ٿ,^Lw�y�@;( ��3@L�0%�!?���>䓕@/��ʹ�ٿ,^Lw�y�@;( ��3@L�0%�!?���>䓕@/��ʹ�ٿ,^Lw�y�@;( ��3@L�0%�!?���>䓕@/��ʹ�ٿ,^Lw�y�@;( ��3@L�0%�!?���>䓕@L����ٿ�����@��\���3@�9�%�!?9o�H�Y�@dśٿ��jٸ��@H\y�*4@��9S�!?�Tr�@�>��ٿOYٝ�@�$�t��3@8���h�!?cHW�w�@�>��ٿOYٝ�@�$�t��3@8���h�!?cHW�w�@���q��ٿ��)�@}tD�4@0��V��!?Pw��@���q��ٿ��)�@}tD�4@0��V��!?Pw��@���q��ٿ��)�@}tD�4@0��V��!?Pw��@R'�p�ٿ�j}>���@}>�g�B4@�{��L�!?-�?@�@;ֹ�Ϡٿ�=n _W�@�K�4@Oe�!��!?�d�<��@;ֹ�Ϡٿ�=n _W�@�K�4@Oe�!��!?�d�<��@;ֹ�Ϡٿ�=n _W�@�K�4@Oe�!��!?�d�<��@;ֹ�Ϡٿ�=n _W�@�K�4@Oe�!��!?�d�<��@;ֹ�Ϡٿ�=n _W�@�K�4@Oe�!��!?�d�<��@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@���㝟ٿ������@S�CdL4@H�'q��!?�vԕ@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@Zi¶�ٿ��<�d�@��~J�4@-�$��!?��lG뵕@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@���]A�ٿ �z�@�<��4@���tv�!?�
dqy��@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@N�c��ٿ�0p�t��@�ʊP��3@���G�!?���|�@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�����ٿ6�4ٗ�@���o �3@��QT�!?������@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@�'�	Ԡٿ�|6L���@3�n'4@9x�}]�!?�0�Zs�@��zv�ٿ�Ï�7��@+דH4@�K�gu�!?��t�N��@i(�{�ٿ������@C�ǣE�3@`�m�,�!?�5;��@i(�{�ٿ������@C�ǣE�3@`�m�,�!?�5;��@i(�{�ٿ������@C�ǣE�3@`�m�,�!?�5;��@�os-�ٿi� ݪ��@I/H�4@��@�h�!?!�+��@�os-�ٿi� ݪ��@I/H�4@��@�h�!?!�+��@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L��s��ٿ�� ֪C�@
1�4@U�q�P�!?�4ױI�@L7j��ٿq'}+���@��]h(4@�/>�G�!?e�1��@L7j��ٿq'}+���@��]h(4@�/>�G�!?e�1��@L7j��ٿq'}+���@��]h(4@�/>�G�!?e�1��@L7j��ٿq'}+���@��]h(4@�/>�G�!?e�1��@��uƥ�ٿ��c��@7n���]4@���+Q�!?cꝹ9ە@��uƥ�ٿ��c��@7n���]4@���+Q�!?cꝹ9ە@��uƥ�ٿ��c��@7n���]4@���+Q�!?cꝹ9ە@��uƥ�ٿ��c��@7n���]4@���+Q�!?cꝹ9ە@��uƥ�ٿ��c��@7n���]4@���+Q�!?cꝹ9ە@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@��9�ٿ5o��C��@�9+;>84@�7�<�!?ݦm�~��@7�ɛ��ٿ�I_w��@߬�6�j4@*��P�!?���Aѕ@7�ɛ��ٿ�I_w��@߬�6�j4@*��P�!?���Aѕ@�0�w�ٿ�%Q��t�@�6g�A4@��?,+�!?��].��@�0�w�ٿ�%Q��t�@�6g�A4@��?,+�!?��].��@�0�w�ٿ�%Q��t�@�6g�A4@��?,+�!?��].��@�q�0��ٿ���0|��@���w.4@�`�=Ϗ!?�����@�q�0��ٿ���0|��@���w.4@�`�=Ϗ!?�����@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@��/���ٿcIa"��@
V���3@X��|R�!?D(84�@<�TJ�ٿ��$.��@�z�] 4@k���C�!?6�i�mϕ@<�TJ�ٿ��$.��@�z�] 4@k���C�!?6�i�mϕ@�cQ�ٿ<�9���@�x�#4@Fٺ�H�!?c)����@�cQ�ٿ<�9���@�x�#4@Fٺ�H�!?c)����@�cQ�ٿ<�9���@�x�#4@Fٺ�H�!?c)����@X�7�јٿHr6x��@M�4@���{T�!?��i1��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@̰;���ٿ pf���@j���
4@_�;mX�!?uH+W��@��l��ٿH����@?r��A4@�F�m�!?�"Uɕ@��l��ٿH����@?r��A4@�F�m�!?�"Uɕ@��l��ٿH����@?r��A4@�F�m�!?�"Uɕ@��l��ٿH����@?r��A4@�F�m�!?�"Uɕ@��l��ٿH����@?r��A4@�F�m�!?�"Uɕ@.��ٿ,�7���@	l�T.4@s�f]�!?��N{�@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�f���ٿĠ ���@�.�&4@k-�=:�!?§�%�ӕ@�Yp�|�ٿ�˪��@�hI�Q4@Z�3�9�!?d��ځ��@�Yp�|�ٿ�˪��@�hI�Q4@Z�3�9�!?d��ځ��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@X {���ٿ��B1��@g��>14@)�;�l�!?����3��@�O���ٿ�V�D�@�{�&�u4@��s��!?��k_��@�O���ٿ�V�D�@�{�&�u4@��s��!?��k_��@�O���ٿ�V�D�@�{�&�u4@��s��!?��k_��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@���e�ٿ�p���@�g�Wxi4@�;ܦ�!?3�0��@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@I)?�ԝٿ�2�O��@�|e���3@��焐!?�m
�@P��Yo�ٿ���0�W�@ ��/4@�6J�}�!?SG#��ە@P��Yo�ٿ���0�W�@ ��/4@�6J�}�!?SG#��ە@P��Yo�ٿ���0�W�@ ��/4@�6J�}�!?SG#��ە@P��Yo�ٿ���0�W�@ ��/4@�6J�}�!?SG#��ە@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@�s��ٿ����k��@���E4@���u�!?��ـ̗�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@��R��ٿ�#� �@�y�D=4@�[�ֆ�!?��r�K>�@E��ٿ��_�B��@���4A 4@^���P�!?����2&�@E��ٿ��_�B��@���4A 4@^���P�!?����2&�@�����ٿCi�h�)�@�(�3:4@و�Aw�!?�%k��@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@4❠�ٿ!c%pE��@kݼz�4@�f$Q�!?F�Uޕ@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@��YKc�ٿ��Vo�@��`�p4@n�M�!?�r�r�ו@.~�yI�ٿ��iN�k�@�chw�U4@m��U@�!?G�h ��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@�b�c��ٿ0H��(�@2Յ��^4@J)�W��!?�A�e��@9w�aיٿ4ī�J�@1���R4@)Q޾��!?�)��H�@9w�aיٿ4ī�J�@1���R4@)Q޾��!?�)��H�@b� ��ٿ��խ��@���'�*4@6���j�!?�3O�ɕ@���4�ٿ�J�w���@U����4@�-4�[�!?��m.��@���4�ٿ�J�w���@U����4@�-4�[�!?��m.��@���]�ٿ�R�-�W�@��	u$4@�L��Q�!?8�UF4�@���]�ٿ�R�-�W�@��	u$4@�L��Q�!?8�UF4�@���]�ٿ�R�-�W�@��	u$4@�L��Q�!?8�UF4�@���]�ٿ�R�-�W�@��	u$4@�L��Q�!?8�UF4�@�Ǿ��ٿ�zT6��@Ɍ+�G4@�?��T�!?&NU��!�@�Ǿ��ٿ�zT6��@Ɍ+�G4@�?��T�!?&NU��!�@�Ǿ��ٿ�zT6��@Ɍ+�G4@�?��T�!?&NU��!�@z�Wy��ٿ��r��Y�@8Ku��#4@E8(zP�!?�'7�w�@z�Wy��ٿ��r��Y�@8Ku��#4@E8(zP�!?�'7�w�@z�Wy��ٿ��r��Y�@8Ku��#4@E8(zP�!?�'7�w�@z�Wy��ٿ��r��Y�@8Ku��#4@E8(zP�!?�'7�w�@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@��|ۢٿwB@��7�@<�<[D4@��G�~�!?�[p�r��@?'*�ٿh�u�2�@c�X,��3@���m�!?��D����@?'*�ٿh�u�2�@c�X,��3@���m�!?��D����@i'�W*�ٿ�5���@)x4@
?/$��!?HZ
��@u�� $�ٿ2S����@$$��4@gA�o�!?4o��ƕ@u�� $�ٿ2S����@$$��4@gA�o�!?4o��ƕ@u�� $�ٿ2S����@$$��4@gA�o�!?4o��ƕ@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@j0�ٿ��<��@�^��~4@Jg�T�!?FC��h��@�����ٿ���8�G�@�m���4@0(Q��!?J���@�rV}z�ٿ1V�Ny��@EIx��3@Pv�d��!?e��w��@�rV}z�ٿ1V�Ny��@EIx��3@Pv�d��!?e��w��@�rV}z�ٿ1V�Ny��@EIx��3@Pv�d��!?e��w��@�rV}z�ٿ1V�Ny��@EIx��3@Pv�d��!?e��w��@�rV}z�ٿ1V�Ny��@EIx��3@Pv�d��!?e��w��@�B\׭�ٿ�#�K���@:h�R 4@o6��y�!?�eәܕ@�B\׭�ٿ�#�K���@:h�R 4@o6��y�!?�eәܕ@�B\׭�ٿ�#�K���@:h�R 4@o6��y�!?�eәܕ@�B\׭�ٿ�#�K���@:h�R 4@o6��y�!?�eәܕ@�B\׭�ٿ�#�K���@:h�R 4@o6��y�!?�eәܕ@�?P�c�ٿxKEE>�@��^�4@����Ð!?6��-��@�?P�c�ٿxKEE>�@��^�4@����Ð!?6��-��@�?P�c�ٿxKEE>�@��^�4@����Ð!?6��-��@]&����ٿ\��I3��@ K���3@��uՐ�!?���W���@]&����ٿ\��I3��@ K���3@��uՐ�!?���W���@]&����ٿ\��I3��@ K���3@��uՐ�!?���W���@]&����ٿ\��I3��@ K���3@��uՐ�!?���W���@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@ӟ}��ٿ��vc;
�@oC�-4@m�?�^�!?h��@�ו@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@)�ሙ�ٿš1)g-�@�
G��-4@Y��Db�!?��TA��@-3����ٿ�5�{�x�@���4@�q��!?A�,�c��@2ˀ�l�ٿ�
�>��@oo�Wk;4@�dHᦐ!?˄kȕ@2ˀ�l�ٿ�
�>��@oo�Wk;4@�dHᦐ!?˄kȕ@2ˀ�l�ٿ�
�>��@oo�Wk;4@�dHᦐ!?˄kȕ@2ˀ�l�ٿ�
�>��@oo�Wk;4@�dHᦐ!?˄kȕ@%��z�ٿ��++A�@�ۿJ
4@vO�ʐ�!?�7�$���@%��z�ٿ��++A�@�ۿJ
4@vO�ʐ�!?�7�$���@[���ٗٿ�jz�@����*4@�ޥP`�!?<˫>��@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�.��ٿ�.��ȡ�@`ESk�'4@��@b�!?���בc�@�1��r�ٿ�2�[T��@i��1>4@�o�gb�!?��w�}�@�1��r�ٿ�2�[T��@i��1>4@�o�gb�!?��w�}�@�1��r�ٿ�2�[T��@i��1>4@�o�gb�!?��w�}�@�1��r�ٿ�2�[T��@i��1>4@�o�gb�!?��w�}�@�ͦC�ٿ��悀�@i�.(_4@�C��U�!?�(�mR6�@�����ٿs屿L�@ˮ��'a4@���2C�!?�s���@�����ٿs屿L�@ˮ��'a4@���2C�!?�s���@�����ٿs屿L�@ˮ��'a4@���2C�!?�s���@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@��C�#�ٿ�~�"�@���2�L4@!6��!?
��u�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@����ٿ8@^���@�{F�

4@��K�!?�� ��-�@��
��ٿU����@v˭��84@ ���!?��M�+�@��
��ٿU����@v˭��84@ ���!?��M�+�@��
��ٿU����@v˭��84@ ���!?��M�+�@�)��u�ٿ��"��@�O�j�)4@ �F7+�!?������@�)��u�ٿ��"��@�O�j�)4@ �F7+�!?������@�)��u�ٿ��"��@�O�j�)4@ �F7+�!?������@�)��u�ٿ��"��@�O�j�)4@ �F7+�!?������@�)��u�ٿ��"��@�O�j�)4@ �F7+�!?������@�4m���ٿl���	��@�܊��#4@Fu`�l�!?�ǽb.�@�4m���ٿl���	��@�܊��#4@Fu`�l�!?�ǽb.�@�4m���ٿl���	��@�܊��#4@Fu`�l�!?�ǽb.�@���9ΝٿPDM���@G�QY:(4@H��as�!? |����@�%�R��ٿ>}PFt��@W�w�_4@T��d�!?�2,A:�@�%�R��ٿ>}PFt��@W�w�_4@T��d�!?�2,A:�@-�߳:�ٿ���2�+�@ݚ$��y4@b�/\�!?�^n��@-�߳:�ٿ���2�+�@ݚ$��y4@b�/\�!?�^n��@zD$�ٿ'��R���@�)��84@�U�E��!?'����@zD$�ٿ'��R���@�)��84@�U�E��!?'����@zD$�ٿ'��R���@�)��84@�U�E��!?'����@N����ٿ�嵋k�@��E/=4@A�R7��!?.��	�@N����ٿ�嵋k�@��E/=4@A�R7��!?.��	�@� �2��ٿ<�ݟ��@�̲Y4@hUא!?߯��	�@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@���F�ٿ�`wL+�@a��B>4@�x˵��!?֕���@�� ��ٿ:���k8�@�!�߽4@�Y[�q�!?ҎJ5@�� ��ٿ:���k8�@�!�߽4@�Y[�q�!?ҎJ5@�� ��ٿ:���k8�@�!�߽4@�Y[�q�!?ҎJ5@�� ��ٿ:���k8�@�!�߽4@�Y[�q�!?ҎJ5@�� ��ٿ:���k8�@�!�߽4@�Y[�q�!?ҎJ5@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@B�%�ٿ`��=�@p'���/4@^�z��!?FS��Օ@*�`=&�ٿ������@6�if,$4@�U��g�!?�ܥY|/�@*�`=&�ٿ������@6�if,$4@�U��g�!?�ܥY|/�@*�`=&�ٿ������@6�if,$4@�U��g�!?�ܥY|/�@*�`=&�ٿ������@6�if,$4@�U��g�!?�ܥY|/�@]Fv3�ٿ(��B���@lD�`�4@f-ȍ��!?�s��@]Fv3�ٿ(��B���@lD�`�4@f-ȍ��!?�s��@]Fv3�ٿ(��B���@lD�`�4@f-ȍ��!?�s��@]Fv3�ٿ(��B���@lD�`�4@f-ȍ��!?�s��@]Fv3�ٿ(��B���@lD�`�4@f-ȍ��!?�s��@J ���ٿ^,�S�P�@��s_e24@�Y�ȣ�!?2�m��Õ@J ���ٿ^,�S�P�@��s_e24@�Y�ȣ�!?2�m��Õ@J ���ٿ^,�S�P�@��s_e24@�Y�ȣ�!?2�m��Õ@J ���ٿ^,�S�P�@��s_e24@�Y�ȣ�!?2�m��Õ@J ���ٿ^,�S�P�@��s_e24@�Y�ȣ�!?2�m��Õ@���p�ٿo�rJ�@Yw���'4@P�T�!?��Yc�@���p�ٿo�rJ�@Yw���'4@P�T�!?��Yc�@��Lp~�ٿ+Y�Y��@��$?��3@��h�U�!?Иl�+^�@3�E�ٿ��V��-�@�П64@��t��!? �j=�@�S���ٿ���0��@�4��v	4@�6���!?�\q5���@�S���ٿ���0��@�4��v	4@�6���!?�\q5���@�W����ٿې�߃X�@�pA>�Q4@���a�!?�>�P��@�W����ٿې�߃X�@�pA>�Q4@���a�!?�>�P��@�W����ٿې�߃X�@�pA>�Q4@���a�!?�>�P��@�W����ٿې�߃X�@�pA>�Q4@���a�!?�>�P��@�W����ٿې�߃X�@�pA>�Q4@���a�!?�>�P��@[�,���ٿ7�(��M�@�{�-24@V�߷�!?~���@[�,���ٿ7�(��M�@�{�-24@V�߷�!?~���@[�,���ٿ7�(��M�@�{�-24@V�߷�!?~���@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@#zy�{�ٿ��
C�M�@~�w�m'4@�����!?%\�I��@�5@D�ٿ�A!=MZ�@L򔩂E4@�7�겐!?Q��ΐ֕@�5@D�ٿ�A!=MZ�@L򔩂E4@�7�겐!?Q��ΐ֕@�5@D�ٿ�A!=MZ�@L򔩂E4@�7�겐!?Q��ΐ֕@s�D���ٿU66|�@�2��14@���z��!?bgd���@s�D���ٿU66|�@�2��14@���z��!?bgd���@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@ �F�:�ٿ�S"����@*�(�#4@/KzL�!?�~`=-��@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@�>*yӚٿ�(��;��@[�B-I4@b�Krj�!?rX�}���@߄���ٿ^<��8�@��E4@���Lv�!?"~Q����@�;ݙ�ٿ�y�����@���2�/4@��sy~�!?�"��.��@�;ݙ�ٿ�y�����@���2�/4@��sy~�!?�"��.��@�;ݙ�ٿ�y�����@���2�/4@��sy~�!?�"��.��@�;ݙ�ٿ�y�����@���2�/4@��sy~�!?�"��.��@�;ݙ�ٿ�y�����@���2�/4@��sy~�!?�"��.��@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@7(]Ϝٿ����o�@���h!4@Ù�Z�!?�F�yu0�@ �*��ٿ{����@2C5<]4@(CzL�!?��s��@ �*��ٿ{����@2C5<]4@(CzL�!?��s��@rG�7ԡٿZ���H�@���X4@�\�Z?�!?�	�!zd�@rG�7ԡٿZ���H�@���X4@�\�Z?�!?�	�!zd�@�I0d�ٿ���#���@c�φ_'4@k0�G"�!?�?Jp�n�@�I0d�ٿ���#���@c�φ_'4@k0�G"�!?�?Jp�n�@��9�ٿL�1�@y�;��4@Y�?]�!?������@��9�ٿL�1�@y�;��4@Y�?]�!?������@��9�ٿL�1�@y�;��4@Y�?]�!?������@��9�ٿL�1�@y�;��4@Y�?]�!?������@��9�ٿL�1�@y�;��4@Y�?]�!?������@$��Cl�ٿ�dۇO�@YD"a#4@�U���!?���>��@$��Cl�ٿ�dۇO�@YD"a#4@�U���!?���>��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@�e����ٿ�h��@�v4@Fؔ���!?Q#r��@-З��ٿnx3G>�@���a�44@>Ւr�!?����o�@ǻ��M�ٿ�_�jü�@w^�?�/4@����q�!?gz�@ǻ��M�ٿ�_�jü�@w^�?�/4@����q�!?gz�@ǻ��M�ٿ�_�jü�@w^�?�/4@����q�!?gz�@�����ٿpRwc{�@8b �#'4@kBa��!?�&OlO&�@�����ٿpRwc{�@8b �#'4@kBa��!?�&OlO&�@�����ٿpRwc{�@8b �#'4@kBa��!?�&OlO&�@�����ٿpRwc{�@8b �#'4@kBa��!?�&OlO&�@��J�ٿNb�j���@�?�(14@	��d�!?��Z��*�@��J�ٿNb�j���@�?�(14@	��d�!?��Z��*�@8����ٿ���8�@�˲�S?4@�UȚE�!?x�_��@ b���ٿ���Ț��@LSd�� 4@4WA��!?DO�=�@�����ٿ����z�@�#���)4@�Q�S��!?��+���@�����ٿ����z�@�#���)4@�Q�S��!?��+���@��%n�ٿ`3Ne�@��15D4@>\!�|�!?݈j5��@��%n�ٿ`3Ne�@��15D4@>\!�|�!?݈j5��@��%n�ٿ`3Ne�@��15D4@>\!�|�!?݈j5��@��%n�ٿ`3Ne�@��15D4@>\!�|�!?݈j5��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@���*�ٿY��0��@ۭN�;C4@��ڈ��!?$>�A��@�����ٿ^i��K\�@��6�4@�✐!?3ӂ���@�����ٿ^i��K\�@��6�4@�✐!?3ӂ���@�����ٿ^i��K\�@��6�4@�✐!?3ӂ���@�����ٿ^i��K\�@��6�4@�✐!?3ӂ���@�`>u��ٿZS�铻�@�굷�4@�p6X��!?i%J��@
�T�јٿ��\&nV�@��>���3@�~r(��!?���ө�@
�T�јٿ��\&nV�@��>���3@�~r(��!?���ө�@
�T�јٿ��\&nV�@��>���3@�~r(��!?���ө�@
�T�јٿ��\&nV�@��>���3@�~r(��!?���ө�@/�ٿ���3��@�����3@�N�S�!?�I)X�a�@/�ٿ���3��@�����3@�N�S�!?�I)X�a�@�.^=�ٿ��h���@�un�4@����5�!?bG�����@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@z1����ٿ�J��:�@K־Ce4@�����!?ndj^�@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@�����ٿ������@�f�N`4@v�ܼl�!?g� p���@����ٿ�R��'��@Ê��a4@�ʺ���!?xi/E��@����ٿJ3����@�ϙ��m4@��#5�!?��a§�@b�u��ٿح+��U�@�C�)*�3@�6K�M�!?X���a�@b�u��ٿح+��U�@�C�)*�3@�6K�M�!?X���a�@b�u��ٿح+��U�@�C�)*�3@�6K�M�!?X���a�@b�u��ٿح+��U�@�C�)*�3@�6K�M�!?X���a�@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@���ٿ�K�D
��@�B�=G94@}c��!?���PD��@[�@�ϘٿS����@����74@^�z]L�!?�f��v�@�?۾J�ٿ"'�UT,�@?[���Y4@N,�	�!?;�W�u�@�?۾J�ٿ"'�UT,�@?[���Y4@N,�	�!?;�W�u�@�?۾J�ٿ"'�UT,�@?[���Y4@N,�	�!?;�W�u�@��J �ٿ
�0Y���@q�A��V4@��6�!?�A��@��J �ٿ
�0Y���@q�A��V4@��6�!?�A��@��J �ٿ
�0Y���@q�A��V4@��6�!?�A��@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@"�5��ٿ|��hj�@�q���L4@[�D6�!?��/!�ϕ@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@�Q�9��ٿh ��|��@t�V�64@2��#5�!?D�c����@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@���G�ٿm�����@]n�ߦF4@����c�!?�㛷ٕ@�=����ٿ�v�21/�@�����3@�#x��!?	��׬�@(j�lM�ٿ<Tv��@t��A�4@�$�+��!?��0�wޕ@(j�lM�ٿ<Tv��@t��A�4@�$�+��!?��0�wޕ@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@C�;�ٿݵ�A�
�@�>���3@9N4���!?����u��@x�<�ٿt� ��@3i<
��3@��	ߠ�!?H� ��@x�<�ٿt� ��@3i<
��3@��	ߠ�!?H� ��@���pƚٿV�~|��@c�8E4@��x�!?!�B���@���pƚٿV�~|��@c�8E4@��x�!?!�B���@���pƚٿV�~|��@c�8E4@��x�!?!�B���@���pƚٿV�~|��@c�8E4@��x�!?!�B���@���H�ٿ7�}@ה�@VP&C�*4@���_��!?��%�Wϕ@���H�ٿ7�}@ה�@VP&C�*4@���_��!?��%�Wϕ@���H�ٿ7�}@ה�@VP&C�*4@���_��!?��%�Wϕ@���H�ٿ7�}@ה�@VP&C�*4@���_��!?��%�Wϕ@���H�ٿ7�}@ה�@VP&C�*4@���_��!?��%�Wϕ@v��.�ٿFᯁ�c�@X��_ �3@�n@]�!?P�ytՕ@v��.�ٿFᯁ�c�@X��_ �3@�n@]�!?P�ytՕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@�Z�ןٿ�:���@u��?4@P3��4�!?�h��0ȕ@����k�ٿ/� 5��@~�:i�3@��{f�!?z�/u�*�@����k�ٿ/� 5��@~�:i�3@��{f�!?z�/u�*�@�
��ٿ)������@��@��3@ 7�o�!?�O��ϕ@Nt+��ٿt�Jh���@�C�I��3@dB�o�!?� �7!��@Nt+��ٿt�Jh���@�C�I��3@dB�o�!?� �7!��@ b酀�ٿ)�2ذ|�@N1�)4@a��V�!?n+����@*+k��ٿ��#z���@��	�-4@�l,WJ�!??��A�@4�=��ٿ��=����@�/
��54@)�2d�!?&��@4�=��ٿ��=����@�/
��54@)�2d�!?&��@��@{i�ٿ�����@6��/(4@S��!T�!?X:,5{�@��@{i�ٿ�����@6��/(4@S��!T�!?X:,5{�@ҚsH�ٿ��7|_�@8��;�3@��5r�!??��@ҚsH�ٿ��7|_�@8��;�3@��5r�!??��@ҚsH�ٿ��7|_�@8��;�3@��5r�!??��@ҚsH�ٿ��7|_�@8��;�3@��5r�!??��@�e��x�ٿE����@Ѿ&�3@�;8|�!?v���˕@�e��x�ٿE����@Ѿ&�3@�;8|�!?v���˕@�e��x�ٿE����@Ѿ&�3@�;8|�!?v���˕@�e��x�ٿE����@Ѿ&�3@�;8|�!?v���˕@\��r�ٿ)K֯���@��)�3@6�ٌ�!?N��5�@\��r�ٿ)K֯���@��)�3@6�ٌ�!?N��5�@\��r�ٿ)K֯���@��)�3@6�ٌ�!?N��5�@\��r�ٿ)K֯���@��)�3@6�ٌ�!?N��5�@E��br�ٿ5�-nĦ�@��N ��3@M��zM�!?#��w>�@E��br�ٿ5�-nĦ�@��N ��3@M��zM�!?#��w>�@l�s2��ٿ�����@�Mu6;�3@��m���!?tYҘ)�@`��T͜ٿ��A{�3�@6\����3@h�Q�`�!?���/��@os#��ٿ�<|M,�@����3@�D�2�!?�e�ȅΕ@os#��ٿ�<|M,�@����3@�D�2�!?�e�ȅΕ@�Λʜٿ��n�0�@����3@ F�*�!?l!��ҕ@�Λʜٿ��n�0�@����3@ F�*�!?l!��ҕ@�Λʜٿ��n�0�@����3@ F�*�!?l!��ҕ@�Λʜٿ��n�0�@����3@ F�*�!?l!��ҕ@1�!��ٿ-�j��@�m|T)4@��zT�!?��X�E�@1�!��ٿ-�j��@�m|T)4@��zT�!?��X�E�@1�!��ٿ-�j��@�m|T)4@��zT�!?��X�E�@P�MN��ٿFq���@��8��3@i�_�2�!?�}-��@P�MN��ٿFq���@��8��3@i�_�2�!?�}-��@P�MN��ٿFq���@��8��3@i�_�2�!?�}-��@���
�ٿ�uC��P�@�dD4@ǌ��A�!?�=C���@���
�ٿ�uC��P�@�dD4@ǌ��A�!?�=C���@���
�ٿ�uC��P�@�dD4@ǌ��A�!?�=C���@�]�H�ٿ�U�*5b�@t:f��4@#w�D�!?�Os�_�@��aA�ٿn��6�@۸==�3@GI��Z�!?����c�@��aA�ٿn��6�@۸==�3@GI��Z�!?����c�@��aA�ٿn��6�@۸==�3@GI��Z�!?����c�@ē?0��ٿ�Y>�/�@��%�b�3@���c�!?u	��x\�@F���ٿt�
��@JL���3@�W �h�!?���ݶ�@F���ٿt�
��@JL���3@�W �h�!?���ݶ�@F���ٿt�
��@JL���3@�W �h�!?���ݶ�@F���ٿt�
��@JL���3@�W �h�!?���ݶ�@F���ٿt�
��@JL���3@�W �h�!?���ݶ�@W�����ٿ�[Y�	��@0љ��3@����!?ߋ���@W�����ٿ�[Y�	��@0љ��3@����!?ߋ���@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@�O�n��ٿaiAߏ:�@&�w@�3@�x7�W�!?��Lܩ�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@<�����ٿ��v�p��@{�$RJ4@y�k�!?���W(9�@��(_��ٿ+���j�@���"4@n��=�!?���&�@��(_��ٿ+���j�@���"4@n��=�!?���&�@��(_��ٿ+���j�@���"4@n��=�!?���&�@��(_��ٿ+���j�@���"4@n��=�!?���&�@��(_��ٿ+���j�@���"4@n��=�!?���&�@��(_��ٿ+���j�@���"4@n��=�!?���&�@�ioz��ٿ��J�np�@����"4@G�r�-�!?aў4ɕ@�ioz��ٿ��J�np�@����"4@G�r�-�!?aў4ɕ@@q�]{�ٿbi����@�w_�,4@Y�$MI�!?n)�L�@���ݺ�ٿi��G#�@��l,4@ԕr�!?�jQ��@�t3���ٿΰT&���@�Ȋ׈)4@n��]�!?��O��@�t3���ٿΰT&���@�Ȋ׈)4@n��]�!?��O��@�t3���ٿΰT&���@�Ȋ׈)4@n��]�!?��O��@4�\Rs�ٿֺ�_m�@�ϫ��4@����Y�!?&1��4ѕ@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@'ȼ�c�ٿQH2��@�]�y�3@mo�hP�!?�Yk��%�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@zx�0"�ٿ�sg��b�@��}�4@�h�x��!?a�p3w_�@�ʠ&g�ٿw���W��@�:��k4@�p��x�!?F)�V���@�ʠ&g�ٿw���W��@�:��k4@�p��x�!?F)�V���@�ʠ&g�ٿw���W��@�:��k4@�p��x�!?F)�V���@��]��ٿ3d�i���@��|*54@�|��!?�ښ�T�@��]��ٿ3d�i���@��|*54@�|��!?�ښ�T�@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@¹\��ٿvp�P<�@�Y��)T4@PX1��!?Ť�k���@�I�X�ٿ,./����@�L~��,4@����c�!?B���M�@�I�X�ٿ,./����@�L~��,4@����c�!?B���M�@�I�X�ٿ,./����@�L~��,4@����c�!?B���M�@�I�X�ٿ,./����@�L~��,4@����c�!?B���M�@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@��-Ď�ٿ}ft"���@+���/4@\Z@V�!?M)�(fו@n�mJޙٿ�1�T��@ ��U�&4@9S�!?
��t���@*|(�d�ٿ:�r����@�mV�4@��\�g�!?�+�:+Q�@*|(�d�ٿ:�r����@�mV�4@��\�g�!?�+�:+Q�@^!��H�ٿ ���w2�@���4@Խz+z�!?l*�,�@^!��H�ٿ ���w2�@���4@Խz+z�!?l*�,�@D�.�ٿNK��r�@��nl4@�V�Mb�!?a��5�	�@�և���ٿH/���@���f84@�^��}�!?7d=�c�@ ���ٿ����J�@�G��^4@@�7�!?�^���@ ���ٿ����J�@�G��^4@@�7�!?�^���@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@�V4��ٿ��c�d�@m��TK4@<�p\�!?�C��^�@��P���ٿ�9�~��@"�A�qa4@_�A���!?%,%����@��P���ٿ�9�~��@"�A�qa4@_�A���!?%,%����@��P���ٿ�9�~��@"�A�qa4@_�A���!?%,%����@��P���ٿ�9�~��@"�A�qa4@_�A���!?%,%����@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@���!�ٿ<:Vj�&�@f/f�V]4@�����!?hs�%ԕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@����ٿ��5�'�@N���4@Eׯo�!?�v��ŕ@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�ڭ{��ٿ,�c�@����'�3@��RW�!?K7Sm���@�g�K�ٿ���!�@T��z"4@���f�!?��5����@���ĕٿ�1K!�@��)�3@�ٍ�N�!?�A��D�@���ĕٿ�1K!�@��)�3@�ٍ�N�!?�A��D�@���ĕٿ�1K!�@��)�3@�ٍ�N�!?�A��D�@���ĕٿ�1K!�@��)�3@�ٍ�N�!?�A��D�@GZ%�Ӛٿ"�d�m!�@��O��3@���I�!?���+{�@GZ%�Ӛٿ"�d�m!�@��O��3@���I�!?���+{�@GZ%�Ӛٿ"�d�m!�@��O��3@���I�!?���+{�@��?Z�ٿ�����	�@�bQ�C4@W6V ��!?,M�M�@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@�Q <��ٿ3ܨ���@�ș�"�3@T�Fw�!?�m���@���Οٿ��5n�J�@+�H�4<4@\��)m�!?���� o�@���Οٿ��5n�J�@+�H�4<4@\��)m�!?���� o�@��l��ٿh�/.��@��t�34@�#RHd�!?Y��3D�@�w4<L�ٿT��ч�@;���*4@��o���!?�@�A%�@�w4<L�ٿT��ч�@;���*4@��o���!?�@�A%�@r�%m�ٿ1̯�݌�@��4Q4@D�"�_�!?8E��6�@��e �ٿ3�64�A�@n��y�4@��C>�!? 6�u�K�@��e �ٿ3�64�A�@n��y�4@��C>�!? 6�u�K�@��e �ٿ3�64�A�@n��y�4@��C>�!? 6�u�K�@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@�h��\�ٿ�e]	��@ߴ��4@؅�6D�!?�S�ݕ@B{�9�ٿ��5���@A�o#�B4@�֋0r�!?�
#�:��@B{�9�ٿ��5���@A�o#�B4@�֋0r�!?�
#�:��@B{�9�ٿ��5���@A�o#�B4@�֋0r�!?�
#�:��@�^�'�ٿ�	�`�@�s���4@����V�!?����@�^�'�ٿ�	�`�@�s���4@����V�!?����@�^�'�ٿ�	�`�@�s���4@����V�!?����@�^�'�ٿ�	�`�@�s���4@����V�!?����@��$q�ٿ2$S���@McB`�3@��?
��!?�aIҡ��@!:H%>�ٿlݤ�@�WQj�3@1bۃd�!?kFLh�@!:H%>�ٿlݤ�@�WQj�3@1bۃd�!?kFLh�@!:H%>�ٿlݤ�@�WQj�3@1bۃd�!?kFLh�@ex��%�ٿ-%b>��@㓹�D�3@��yL�!?w�c�mO�@ex��%�ٿ-%b>��@㓹�D�3@��yL�!?w�c�mO�@�VQ��ٿ�l~��@�e�S��3@��s��!?�u���@�VQ��ٿ�l~��@�e�S��3@��s��!?�u���@�VQ��ٿ�l~��@�e�S��3@��s��!?�u���@نV��ٿ�4Y���@dP`a4@`�X9h�!?<�m%��@��?i�ٿ0������@�5��{	4@�ɀ��!?Q�Z�ĕ@��?i�ٿ0������@�5��{	4@�ɀ��!?Q�Z�ĕ@��?i�ٿ0������@�5��{	4@�ɀ��!?Q�Z�ĕ@��?i�ٿ0������@�5��{	4@�ɀ��!?Q�Z�ĕ@��?i�ٿ0������@�5��{	4@�ɀ��!?Q�Z�ĕ@=�u���ٿ���|e��@��:�F4@������!?�&p���@=�u���ٿ���|e��@��:�F4@������!?�&p���@=�u���ٿ���|e��@��:�F4@������!?�&p���@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@)�Jx�ٿ�s�+�@Z�?cP44@K��^w�!?��G?��@|^�N��ٿ��bM���@;f����3@��Ǐ��!?L��,��@|^�N��ٿ��bM���@;f����3@��Ǐ��!?L��,��@|^�N��ٿ��bM���@;f����3@��Ǐ��!?L��,��@;��|Πٿ&�GJ���@6M��!4@y�fq�!?9SV�Re�@;��|Πٿ&�GJ���@6M��!4@y�fq�!?9SV�Re�@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@T�l��ٿ�0��'�@�\@4@�q��U�!?0+���@��� �ٿKaUHT�@r1��4@ezd c�!?�É����@��� �ٿKaUHT�@r1��4@ezd c�!?�É����@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@���	�ٿoo�`'��@�p�D��3@���ޗ�!?�d�ƕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�]���ٿҢ�a�&�@,��v4@׺�h�!?_��ԕ@�L̂�ٿ(��%Wo�@�<�Y�;4@̂H0��!?y�|��ԕ@�L̂�ٿ(��%Wo�@�<�Y�;4@̂H0��!?y�|��ԕ@�L̂�ٿ(��%Wo�@�<�Y�;4@̂H0��!?y�|��ԕ@�L̂�ٿ(��%Wo�@�<�Y�;4@̂H0��!?y�|��ԕ@�X�|�ٿ`s�"M�@�����b4@�"�ĉ�!?�!�D�@�X�|�ٿ`s�"M�@�����b4@�"�ĉ�!?�!�D�@�X�|�ٿ`s�"M�@�����b4@�"�ĉ�!?�!�D�@�X�|�ٿ`s�"M�@�����b4@�"�ĉ�!?�!�D�@�J�ؤٿ���;��@n��S%4@qٯ��!?�C{g0ٕ@�J�ؤٿ���;��@n��S%4@qٯ��!?�C{g0ٕ@�J�ؤٿ���;��@n��S%4@qٯ��!?�C{g0ٕ@�mB�ٿ�����@���H_�3@n�t��!?���1�ҕ@�mB�ٿ�����@���H_�3@n�t��!?���1�ҕ@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@���^�ٿN�O�+��@��<*��3@u�8=��!?��qn��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@<�7�ٿ/Al�@�~"K	4@s�˚�!?
͕��@,���ٿ�<�3M�@*S�֭�3@�܄�h�!?��4��@Vԗ���ٿt�����@�}z�X4@���j�!?_��|=6�@Vԗ���ٿt�����@�}z�X4@���j�!?_��|=6�@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@���ٿ�)�>~��@��͂�4@!%�/p�!?#��z���@��~�ٿA��4.D�@~̰k4@�S�w�!?�v,Dx1�@��~�ٿA��4.D�@~̰k4@�S�w�!?�v,Dx1�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@�3��D�ٿx���ί�@Zt^��3@��"eW�!?���}�#�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@j|I��ٿ<����@kE��74@&I2�!?��_7�)�@\���A�ٿȾ�:W��@Uͽ�4@?`�.�!?
���?�@\���A�ٿȾ�:W��@Uͽ�4@?`�.�!?
���?�@י�ܝ�ٿZ��@�@�uX�4@Q7�&j�!?-�����@י�ܝ�ٿZ��@�@�uX�4@Q7�&j�!?-�����@�-8�՜ٿ���u(�@.�]m64@Rx�{^�!?ۀ�z͕@�-8�՜ٿ���u(�@.�]m64@Rx�{^�!?ۀ�z͕@�-8�՜ٿ���u(�@.�]m64@Rx�{^�!?ۀ�z͕@�-8�՜ٿ���u(�@.�]m64@Rx�{^�!?ۀ�z͕@�B��ٿ�7P���@�u�x�3@;`�D�!?U����@�B��ٿ�7P���@�u�x�3@;`�D�!?U����@�B��ٿ�7P���@�u�x�3@;`�D�!?U����@�B��ٿ�7P���@�u�x�3@;`�D�!?U����@�B��ٿ�7P���@�u�x�3@;`�D�!?U����@�Ig;'�ٿr���&��@F��E'4@Wqvw�!?��7\W��@�Ig;'�ٿr���&��@F��E'4@Wqvw�!?��7\W��@�Ig;'�ٿr���&��@F��E'4@Wqvw�!?��7\W��@�Ig;'�ٿr���&��@F��E'4@Wqvw�!?��7\W��@�{n�+�ٿEx���@��v��3@ǧ�s�!?Y�8N�@�<��!�ٿ����7a�@��M�3@#p�/m�!?z�/����@ ��§ٿ/��P!�@/ӓ��Y4@ڞTP�!?�-l*��@ ��§ٿ/��P!�@/ӓ��Y4@ڞTP�!?�-l*��@ ��§ٿ/��P!�@/ӓ��Y4@ڞTP�!?�-l*��@ ��§ٿ/��P!�@/ӓ��Y4@ڞTP�!?�-l*��@��$�l�ٿ����@�tۧ�h4@kF�l�!?P�u
|�@
(5A��ٿGu���g�@��T34@�U=>�!?>r�'3�@
(5A��ٿGu���g�@��T34@�U=>�!?>r�'3�@);Aa�ٿ^� <���@mW�,�4@.I7&�!?�Y����@);Aa�ٿ^� <���@mW�,�4@.I7&�!?�Y����@);Aa�ٿ^� <���@mW�,�4@.I7&�!?�Y����@);Aa�ٿ^� <���@mW�,�4@.I7&�!?�Y����@���5d�ٿ�O�P�@�'0�64@C���s�!?&�:
��@�}�£ٿ�j����@W���:4@�Ce��!?����̑�@��Ow��ٿ"=��(�@?㯲�;4@�����!?����]�@~����ٿ�F���@^�,��"4@�Ѝ��!?��y�EY�@������ٿ"B`���@j$��B4@��� r�!?��\�6�@������ٿ"B`���@j$��B4@��� r�!?��\�6�@p&"ڡٿCu���@�w�1�4@\�x��!?g���Õ@p&"ڡٿCu���@�w�1�4@\�x��!?g���Õ@�
Ls�ٿ������@���s�4@%Ɩ�h�!?D|��˕@�
Ls�ٿ������@���s�4@%Ɩ�h�!?D|��˕@�
Ls�ٿ������@���s�4@%Ɩ�h�!?D|��˕@�
Ls�ٿ������@���s�4@%Ɩ�h�!?D|��˕@�
Ls�ٿ������@���s�4@%Ɩ�h�!?D|��˕@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@��ξ3�ٿ	_�B7Q�@Q�>�'4@�~1-�!?��x�@`�`�ٿ>�z�V�@�xY&D4@�}�1�!?�� ����@`�`�ٿ>�z�V�@�xY&D4@�}�1�!?�� ����@`�`�ٿ>�z�V�@�xY&D4@�}�1�!?�� ����@`�`�ٿ>�z�V�@�xY&D4@�}�1�!?�� ����@}-X���ٿf`�E|L�@���o�4@Ax�he�!?���
%�@}-X���ٿf`�E|L�@���o�4@Ax�he�!?���
%�@}-X���ٿf`�E|L�@���o�4@Ax�he�!?���
%�@}-X���ٿf`�E|L�@���o�4@Ax�he�!?���
%�@}-X���ٿf`�E|L�@���o�4@Ax�he�!?���
%�@�Z{� �ٿ�C��ej�@u�i4@�(K�a�!?Q����A�@�Z{� �ٿ�C��ej�@u�i4@�(K�a�!?Q����A�@�x0�ٿ���&�@��0�&4@�6>��!?4�w(�@�m����ٿp���{�@�� ��3@�L����!?��:_�@�[%�ٿ,U]�mA�@Ct�G��3@�oԣ�!?8�T����@�[%�ٿ,U]�mA�@Ct�G��3@�oԣ�!?8�T����@G҇ՙٿs����b�@.jG� 4@e%�]G�!?�VrH��@G҇ՙٿs����b�@.jG� 4@e%�]G�!?�VrH��@G҇ՙٿs����b�@.jG� 4@e%�]G�!?�VrH��@G҇ՙٿs����b�@.jG� 4@e%�]G�!?�VrH��@W�^X�ٿ�3N�+�@`R{�4@�V�|�!?}i���@W�^X�ٿ�3N�+�@`R{�4@�V�|�!?}i���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@G����ٿ��=
1��@��c@74@D(a�g�!?�~���@�'�Ηٿt�cN��@�����+4@+�h�N�!?��?�@�'�Ηٿt�cN��@�����+4@+�h�N�!?��?�@l'̛ٿ�����@�n�d4@�3��b�!?ǉp��@l'̛ٿ�����@�n�d4@�3��b�!?ǉp��@l'̛ٿ�����@�n�d4@�3��b�!?ǉp��@l'̛ٿ�����@�n�d4@�3��b�!?ǉp��@l'̛ٿ�����@�n�d4@�3��b�!?ǉp��@#(ne�ٿ�)^�ǌ�@cl.��3@�(¤6�!?<�ԛ�@�C�.�ٿ>"��y�@�d!4@�d�$C�!?��U/-h�@�C�.�ٿ>"��y�@�d!4@�d�$C�!?��U/-h�@�C�.�ٿ>"��y�@�d!4@�d�$C�!?��U/-h�@�cKO�ٿ�呪.�@'��4@@B�N�!?7Nw��@Cٿ1���E�@�jh��4@1���!?���n=��@Cٿ1���E�@�jh��4@1���!?���n=��@Cٿ1���E�@�jh��4@1���!?���n=��@Cٿ1���E�@�jh��4@1���!?���n=��@Cٿ1���E�@�jh��4@1���!?���n=��@Cٿ1���E�@�jh��4@1���!?���n=��@�x.��ٿ�B�1J��@r�S� 4@�^%�ې!?��/�u�@#D,���ٿA����@�����3@Iʨ�Ð!?�o���@��,�ٿ�HӜG�@��D�3@��ȫ��!?6�w�m�@��,�ٿ�HӜG�@��D�3@��ȫ��!?6�w�m�@��,�ٿ�HӜG�@��D�3@��ȫ��!?6�w�m�@�ˠ�U�ٿY�Y�^8�@`����3@g(|�!?��9���@�ˠ�U�ٿY�Y�^8�@`����3@g(|�!?��9���@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@L�4��ٿ_�)o?��@]N����3@4�N��!?�3�ρ�@KZ~[��ٿ��^���@KI{�4@�#���!?��i���@KZ~[��ٿ��^���@KI{�4@�#���!?��i���@KZ~[��ٿ��^���@KI{�4@�#���!?��i���@KZ~[��ٿ��^���@KI{�4@�#���!?��i���@KZ~[��ٿ��^���@KI{�4@�#���!?��i���@^֬���ٿ|���,�@YF��4@��Ő!?���)R�@@Q�4v�ٿ��z���@檇�>4@8EI�Đ!?�`UL���@@Q�4v�ٿ��z���@檇�>4@8EI�Đ!?�`UL���@��c��ٿs6x8���@m���/4@W%����!?�?u�Ep�@��c��ٿs6x8���@m���/4@W%����!?�?u�Ep�@��c��ٿs6x8���@m���/4@W%����!?�?u�Ep�@-/��ǚٿ��Rz���@�ڛt%4@���c��!?QQ�po�@w�&�ٿ5�q���@��y4@ �Z9x�!?��f��@w�&�ٿ5�q���@��y4@ �Z9x�!?��f��@�t9
�ٿ���=��@�U�R�Q4@*ƌ!X�!?�������@�t9
�ٿ���=��@�U�R�Q4@*ƌ!X�!?�������@�t9
�ٿ���=��@�U�R�Q4@*ƌ!X�!?�������@�t9
�ٿ���=��@�U�R�Q4@*ƌ!X�!?�������@haڍ�ٿ�p���@�n~ 94@�ɚ�_�!?1V�eV�@haڍ�ٿ�p���@�n~ 94@�ɚ�_�!?1V�eV�@haڍ�ٿ�p���@�n~ 94@�ɚ�_�!?1V�eV�@haڍ�ٿ�p���@�n~ 94@�ɚ�_�!?1V�eV�@haڍ�ٿ�p���@�n~ 94@�ɚ�_�!?1V�eV�@�;P�j�ٿ�9)���@��CX�4@5�s�!?ϘA�'�@�;P�j�ٿ�9)���@��CX�4@5�s�!?ϘA�'�@	|x�ϜٿWgG ��@q�#��L4@��i�!?�~.�T�@GLˢ�ٿ)ÔU�
�@�w�Bk4@�}���!?g�����@�Ύޝٿ�d@o���@�����14@�2��!?c����ҕ@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@q��l�ٿ����D�@2��^�3@A=��:�!?�-O���@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@;'�,��ٿO��K
�@�c��3@5d}��!?q[�UZ�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@�CK�ٿ
�8�43�@�}$��3@�^}�5�!?�f��T�@9=�Qҙٿ�>�]f��@���Y��3@�=��h�!?��u�.�@9=�Qҙٿ�>�]f��@���Y��3@�=��h�!?��u�.�@9=�Qҙٿ�>�]f��@���Y��3@�=��h�!?��u�.�@��%�ٿ$����j�@0�ખ�3@{qaAT�!?7r�o�u�@��%�ٿ$����j�@0�ખ�3@{qaAT�!?7r�o�u�@��%�ٿ$����j�@0�ખ�3@{qaAT�!?7r�o�u�@��%�ٿ$����j�@0�ખ�3@{qaAT�!?7r�o�u�@��%�ٿ$����j�@0�ખ�3@{qaAT�!?7r�o�u�@�#��ƞٿf�?��@6B	�4@W��/<�!?ݱ�Wͺ�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@q�G��ٿ_�E� �@�0w� 4@���6P�!?%f�̢�@�H�ɑ�ٿ�����@,s��e4@3=����!?��$�@�H�ɑ�ٿ�����@,s��e4@3=����!?��$�@��ǭw�ٿ��0�I�@[]ʭ�3@�(��o�!?:�hW��@��ǭw�ٿ��0�I�@[]ʭ�3@�(��o�!?:�hW��@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@���ٿ3�VH���@Ӣ0�;4@�;i�!?��;�C �@@��{�ٿ~��A1��@��DopC4@6�	�k�!?�D/M���@@��{�ٿ~��A1��@��DopC4@6�	�k�!?�D/M���@РO��ٿ�v5=�@׷���;4@�NH�|�!?C�[ �G�@РO��ٿ�v5=�@׷���;4@�NH�|�!?C�[ �G�@РO��ٿ�v5=�@׷���;4@�NH�|�!?C�[ �G�@РO��ٿ�v5=�@׷���;4@�NH�|�!?C�[ �G�@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@�:¿��ٿlSI���@ݮ��4@�j�LH�!?*p�L�Õ@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@G<�0�ٿ~����@��Vw�4@U6�C�!?���a?��@y��"��ٿ�W��?�@�~��44@���W�!?�0�Õ@��[��ٿ]2����@2��4@�&r`f�!?� 7�iٕ@��[��ٿ]2����@2��4@�&r`f�!?� 7�iٕ@��[��ٿ]2����@2��4@�&r`f�!?� 7�iٕ@��(}��ٿ�%��A��@zD�=�4@�f�V?�!?Z5�f��@��(}��ٿ�%��A��@zD�=�4@�f�V?�!?Z5�f��@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@R�uD��ٿ(��F�@�"�b�3@·��}�!?!�&�Ε@����ٿ���@�H�`��3@�ԣ�/�!?0-{��ؕ@����ٿ���@�H�`��3@�ԣ�/�!?0-{��ؕ@����ٿ���@�H�`��3@�ԣ�/�!?0-{��ؕ@�[o���ٿ�%B^�@#��p54@�D�=�!?�r&ŗ�@�[o���ٿ�%B^�@#��p54@�D�=�!?�r&ŗ�@5�n��ٿ��2��s�@�T�{4@w$lP�!?�od*˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@���&G�ٿ�\%*<��@QX�:�4@�M͛��!?Ր�W�˕@;���T�ٿ�- ��@�/�ʊD4@S)bpϐ!?��>FB�@;���T�ٿ�- ��@�/�ʊD4@S)bpϐ!?��>FB�@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@<ʱr��ٿά�\y��@��&#4@!�[6��!?������@��z\�ٿ���%�(�@��:44@;�1��!?��Q�(�@��z\�ٿ���%�(�@��:44@;�1��!?��Q�(�@��z\�ٿ���%�(�@��:44@;�1��!?��Q�(�@U�B?��ٿ�r�Z��@��rɕa4@X�ו��!?7�ˁ�e�@U�B?��ٿ�r�Z��@��rɕa4@X�ו��!?7�ˁ�e�@U�B?��ٿ�r�Z��@��rɕa4@X�ו��!?7�ˁ�e�@U�B?��ٿ�r�Z��@��rɕa4@X�ו��!?7�ˁ�e�@ف�7B�ٿ�ޭ���@ ��(4@"b"]w�!?�v�q��@�t�D�ٿ���=EU�@���844@���[~�!?J'g��N�@�t�D�ٿ���=EU�@���844@���[~�!?J'g��N�@!�~}�ٿϽA���@���34@�ə��!?c�2�@;���7�ٿ��C�a��@s5�)�!4@�1P3ɐ!?�?�K.ȕ@�]���ٿ�F����@�I��94@M��t�!?r��j�˕@�]���ٿ�F����@�I��94@M��t�!?r��j�˕@�]���ٿ�F����@�I��94@M��t�!?r��j�˕@�]���ٿ�F����@�I��94@M��t�!?r��j�˕@�]���ٿ�F����@�I��94@M��t�!?r��j�˕@��<�ٿ�EbS��@�'���4@9[�,�!?~*�#�Օ@��<�ٿ�EbS��@�'���4@9[�,�!?~*�#�Օ@��<�ٿ�EbS��@�'���4@9[�,�!?~*�#�Օ@��<�ٿ�EbS��@�'���4@9[�,�!?~*�#�Օ@��<�ٿ�EbS��@�'���4@9[�,�!?~*�#�Օ@�y��ٿ�;o�V��@��8���3@�����!?����n�@�y��ٿ�;o�V��@��8���3@�����!?����n�@�y��ٿ�;o�V��@��8���3@�����!?����n�@�y��ٿ�;o�V��@��8���3@�����!?����n�@�y��ٿ�;o�V��@��8���3@�����!?����n�@�6�ٔٿZ��:ō�@��3�2
4@�^�
�!?M��إ�@�6�ٔٿZ��:ō�@��3�2
4@�^�
�!?M��إ�@�6�ٔٿZ��:ō�@��3�2
4@�^�
�!?M��إ�@�6�ٔٿZ��:ō�@��3�2
4@�^�
�!?M��إ�@�6�ٔٿZ��:ō�@��3�2
4@�^�
�!?M��إ�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@a�i��ٿ���%4h�@�Qe}kI4@S��J�!?yRE�n�@[��`��ٿ�Kwf��@�/���m4@(�S���!?��c/�@[��`��ٿ�Kwf��@�/���m4@(�S���!?��c/�@[��`��ٿ�Kwf��@�/���m4@(�S���!?��c/�@��8�ٿT�8����@6�/�]14@|52�M�!?7݄:NV�@��8�ٿT�8����@6�/�]14@|52�M�!?7݄:NV�@��8�ٿT�8����@6�/�]14@|52�M�!?7݄:NV�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@��ey�ٿЄV��@�`�N4@�$����!?��p�t�@���葠ٿ������@=~�R)"4@Hi4�!?f�:WÕ@���葠ٿ������@=~�R)"4@Hi4�!?f�:WÕ@���葠ٿ������@=~�R)"4@Hi4�!?f�:WÕ@���葠ٿ������@=~�R)"4@Hi4�!?f�:WÕ@���葠ٿ������@=~�R)"4@Hi4�!?f�:WÕ@�3H���ٿ~Bnx~��@�
立�3@:��j�!?���)Е@�3H���ٿ~Bnx~��@�
立�3@:��j�!?���)Е@�i�Xšٿ�o ���@8X���4@�?�DU�!?��PV;�@�i�Xšٿ�o ���@8X���4@�?�DU�!?��PV;�@~�B�ɛٿ�UQ�v��@>�jw�:4@�����!?��Y2�@~�B�ɛٿ�UQ�v��@>�jw�:4@�����!?��Y2�@~�B�ɛٿ�UQ�v��@>�jw�:4@�����!?��Y2�@~�B�ɛٿ�UQ�v��@>�jw�:4@�����!?��Y2�@�M:NC�ٿ6�����@�S��524@�0����!?D8WX�ݕ@�M:NC�ٿ6�����@�S��524@�0����!?D8WX�ݕ@�M:NC�ٿ6�����@�S��524@�0����!?D8WX�ݕ@�M:NC�ٿ6�����@�S��524@�0����!?D8WX�ݕ@�M:NC�ٿ6�����@�S��524@�0����!?D8WX�ݕ@��?�ٿ��]���@3�0T4@�t'�!?n�\����@��?�ٿ��]���@3�0T4@�t'�!?n�\����@��?�ٿ��]���@3�0T4@�t'�!?n�\����@���4�ٿ�.�-0�@t�T��54@hJK/<�!?�@
Oᾕ@���4�ٿ�.�-0�@t�T��54@hJK/<�!?�@
Oᾕ@���4�ٿ�.�-0�@t�T��54@hJK/<�!?�@
Oᾕ@���4�ٿ�.�-0�@t�T��54@hJK/<�!?�@
Oᾕ@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�fP��ٿP����@������3@����O�!?$��6L�@�����ٿ�3��@O��DV�3@�ȉe��!?T���!�@�����ٿ�3��@O��DV�3@�ȉe��!?T���!�@�����ٿ�3��@O��DV�3@�ȉe��!?T���!�@z0����ٿ2߹���@�����/4@ʊA�!?^����@�f���ٿ�*��]��@$�
�&4@)�v���!?Qf�㿕@�f���ٿ�*��]��@$�
�&4@)�v���!?Qf�㿕@t�|�ٿ�N6�� �@�����>4@1md4�!?��Ќʻ�@+mKr�ٿy�����@����K4@�� ���!?��x����@+mKr�ٿy�����@����K4@�� ���!?��x����@+mKr�ٿy�����@����K4@�� ���!?��x����@+mKr�ٿy�����@����K4@�� ���!?��x����@+mKr�ٿy�����@����K4@�� ���!?��x����@�=�w��ٿp"CB��@%�8%4M4@(�f��!?GK�k��@�=�w��ٿp"CB��@%�8%4M4@(�f��!?GK�k��@�=�w��ٿp"CB��@%�8%4M4@(�f��!?GK�k��@���ٿKV]$�o�@�A���K4@V�WM�!?�����@�����ٿٙ]O%��@ALJэI4@�����!?.�t⤕@�����ٿٙ]O%��@ALJэI4@�����!?.�t⤕@�����ٿٙ]O%��@ALJэI4@�����!?.�t⤕@�/�K��ٿe��H�X�@5Eh	�,4@E=Ÿ��!?���xg��@ب�ߞٿӒ� �Q�@�Ї'��3@��㴀�!?��4��@qq���ٿ��`�@�Ʉ	�3@�OH�!?�sd롷�@qq���ٿ��`�@�Ʉ	�3@�OH�!?�sd롷�@qq���ٿ��`�@�Ʉ	�3@�OH�!?�sd롷�@qq���ٿ��`�@�Ʉ	�3@�OH�!?�sd롷�@qq���ٿ��`�@�Ʉ	�3@�OH�!?�sd롷�@�/�ٿ�q�m���@�����3@�k,-�!?��c�	�@�/�ٿ�q�m���@�����3@�k,-�!?��c�	�@�/�ٿ�q�m���@�����3@�k,-�!?��c�	�@�/�ٿ�q�m���@�����3@�k,-�!?��c�	�@�/�ٿ�q�m���@�����3@�k,-�!?��c�	�@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@s��Ɵٿ�c1�~��@z0�$�24@�?i�7�!?�T����@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@��ߌ�ٿE!)��6�@�׊�&4@jɄ�N�!?����ە@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@�H�?�ٿl&�o9�@�dz�Z4@��9ax�!?Anm��Õ@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@R-�)��ٿcXf���@Z�7H%64@ks�؏!?�z����@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@��Z��ٿ������@E�	��C4@�MJ�!?�k�j���@e����ٿ�l�"�N�@�+�(4@r�w<=�!?�|�?�(�@e����ٿ�l�"�N�@�+�(4@r�w<=�!?�|�?�(�@�r��k�ٿ��;1��@�EV]44@	I��s�!?��:>)�@�1��ٿ��O7���@T���
4@)�k�f�!?J�j$�ܕ@$9�J�ٿ�	;	�@!!K�
4@TYjm�!?��4L�@g$�B�ٿX>����@�d�54@Nԛ���!?]�'_,�@g$�B�ٿX>����@�d�54@Nԛ���!?]�'_,�@g$�B�ٿX>����@�d�54@Nԛ���!?]�'_,�@����ٿ�,�.��@�eY��$4@9�Eu�!?Z!Ӗ�|�@i>���ٿ/�Xԡ��@���z=4@8L����!?.郻r�@i>���ٿ/�Xԡ��@���z=4@8L����!?.郻r�@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@��i�ٿ���dq�@ʇ�ѐ�3@���Z�!?�a�Ҏޕ@ђ��ɛٿ�/ ]:<�@��"{4@��T~8�!?N$_�s��@ђ��ɛٿ�/ ]:<�@��"{4@��T~8�!?N$_�s��@ђ��ɛٿ�/ ]:<�@��"{4@��T~8�!?N$_�s��@ђ��ɛٿ�/ ]:<�@��"{4@��T~8�!?N$_�s��@ђ��ɛٿ�/ ]:<�@��"{4@��T~8�!?N$_�s��@��r�7�ٿ�^'!~��@l���n4@�klt�!?�b�;� �@r�]	��ٿ6o��	��@���͎'4@O*�O�!?�-2��@r�]	��ٿ6o��	��@���͎'4@O*�O�!?�-2��@r�]	��ٿ6o��	��@���͎'4@O*�O�!?�-2��@r�]	��ٿ6o��	��@���͎'4@O*�O�!?�-2��@r�]	��ٿ6o��	��@���͎'4@O*�O�!?�-2��@c�=�5�ٿ��[��@ؼJ��44@E_٧]�!?)��8ܕ@c�=�5�ٿ��[��@ؼJ��44@E_٧]�!?)��8ܕ@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�+�қٿ̕��p��@~{�U14@O$V�!?�"U(�Е@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@�����ٿw��;��@�LN>'4@�#�슐!?d}�t���@���<ŗٿ�툫��@����4@HH�Q�!?*�+�B/�@���<ŗٿ�툫��@����4@HH�Q�!?*�+�B/�@���<ŗٿ�툫��@����4@HH�Q�!?*�+�B/�@Q�LI.�ٿ� ��u��@2��3@�8�6�!?����"�@Q�LI.�ٿ� ��u��@2��3@�8�6�!?����"�@�C� Q�ٿ���"��@r�}��3@E�*[�!?,�D'��@�C� Q�ٿ���"��@r�}��3@E�*[�!?,�D'��@;\�hM�ٿ���[���@�����3@po�!?������@;\�hM�ٿ���[���@�����3@po�!?������@;\�hM�ٿ���[���@�����3@po�!?������@;\�hM�ٿ���[���@�����3@po�!?������@;\�hM�ٿ���[���@�����3@po�!?������@e�[{�ٿ��z-�@N�K�684@>�J@�!?�t�U���@e�[{�ٿ��z-�@N�K�684@>�J@�!?�t�U���@e�[{�ٿ��z-�@N�K�684@>�J@�!?�t�U���@e�[{�ٿ��z-�@N�K�684@>�J@�!?�t�U���@e�[{�ٿ��z-�@N�K�684@>�J@�!?�t�U���@��ېW�ٿ� t�l�@|t�!�4@��;�!?z�qLH�@��ېW�ٿ� t�l�@|t�!�4@��;�!?z�qLH�@��ېW�ٿ� t�l�@|t�!�4@��;�!?z�qLH�@��ېW�ٿ� t�l�@|t�!�4@��;�!?z�qLH�@��ېW�ٿ� t�l�@|t�!�4@��;�!?z�qLH�@��B��ٿZ�t6��@�U��3@b"���!?�h���@�:%�#�ٿv�TGw��@&���D�3@$�][f�!?獇���@�:%�#�ٿv�TGw��@&���D�3@$�][f�!?獇���@�:%�#�ٿv�TGw��@&���D�3@$�][f�!?獇���@,���ٿ��̴��@�����3@���Ư�!?�.d�x�@5��켡ٿn6�_���@���F�04@��z�!?�;(�@D��r?�ٿ�'?�5�@	���84@�D8��!?�X�Tϕ@D��r?�ٿ�'?�5�@	���84@�D8��!?�X�Tϕ@��5,��ٿ���7��@x�j��14@R\�6�!?B�]���@��5,��ٿ���7��@x�j��14@R\�6�!?B�]���@��5,��ٿ���7��@x�j��14@R\�6�!?B�]���@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@�*V﹣ٿ�w5���@]��#4@���[�!?�jz��@u�C�Y�ٿ��ҽ��@^�.�'4@X9�P�!?�V�(�@u�C�Y�ٿ��ҽ��@^�.�'4@X9�P�!?�V�(�@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@I(}xw�ٿ���#�V�@p�lS�#4@1bj�S�!?��f��@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@��,�ٿ�:�����@�y�A54@���_�!?~�c~�@\��.�ٿ��J��@&����@4@֝H�!?{d8͒ߕ@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@��՚ٿ��߰��@"���\*4@���JK�!?ג;u5�@+�ӸJ�ٿ���TD�@� fW�,4@$%ӟm�!?��(�@+�ӸJ�ٿ���TD�@� fW�,4@$%ӟm�!?��(�@+�ӸJ�ٿ���TD�@� fW�,4@$%ӟm�!?��(�@f2��ٿu|r�(�@C�2�=J4@��d��!?����u�@f2��ٿu|r�(�@C�2�=J4@��d��!?����u�@f2��ٿu|r�(�@C�2�=J4@��d��!?����u�@f2��ٿu|r�(�@C�2�=J4@��d��!?����u�@f2��ٿu|r�(�@C�2�=J4@��d��!?����u�@�ܗٿ�&�5�*�@����44@��	���!?�M]ؑ��@�ܗٿ�&�5�*�@����44@��	���!?�M]ؑ��@�ܗٿ�&�5�*�@����44@��	���!?�M]ؑ��@�ܗٿ�&�5�*�@����44@��	���!?�M]ؑ��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@���ٿ��dd��@���%�X4@�}����!?�{�])��@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@y�֞=�ٿ��R�/$�@��j
��3@~H��a�!?ͷc6�@05��:�ٿ�2���@��_�
4@�q:`^�!?����JR�@05��:�ٿ�2���@��_�
4@�q:`^�!?����JR�@05��:�ٿ�2���@��_�
4@�q:`^�!?����JR�@��m�g�ٿ�=��x�@���w4@�m�Tj�!?�{�Ԙ˕@��m�g�ٿ�=��x�@���w4@�m�Tj�!?�{�Ԙ˕@��m�g�ٿ�=��x�@���w4@�m�Tj�!?�{�Ԙ˕@����ٿ~��Q��@��E:�4@��`FP�!?��
��@����ٿ~��Q��@��E:�4@��`FP�!?��
��@����ٿ~��Q��@��E:�4@��`FP�!?��
��@����ٿ~��Q��@��E:�4@��`FP�!?��
��@����ٿ~��Q��@��E:�4@��`FP�!?��
��@���U��ٿ���Zw��@8���o94@���k�!?��� O��@���U��ٿ���Zw��@8���o94@���k�!?��� O��@���U��ٿ���Zw��@8���o94@���k�!?��� O��@���U��ٿ���Zw��@8���o94@���k�!?��� O��@a~RYٿ<GIF���@m+�v<4@�(D҃�!?��S��Q�@a~RYٿ<GIF���@m+�v<4@�(D҃�!?��S��Q�@a~RYٿ<GIF���@m+�v<4@�(D҃�!?��S��Q�@a~RYٿ<GIF���@m+�v<4@�(D҃�!?��S��Q�@�ZśٿZ����@3���4@!mrs�!?�����@�ZśٿZ����@3���4@!mrs�!?�����@�ZśٿZ����@3���4@!mrs�!?�����@�ZśٿZ����@3���4@!mrs�!?�����@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@Yl�q*�ٿ,Z��]�@.�S34@��z�Ð!?�+4�V�@�#5�P�ٿ�Hv
���@���[�4@,:]��!?>���j��@�#5�P�ٿ�Hv
���@���[�4@,:]��!?>���j��@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@
����ٿ4p�����@Hz2$`�3@���]q�!?��]���@��Nt۠ٿX�b�v��@��q|�3@��!WO�!?v�w�~�@��Nt۠ٿX�b�v��@��q|�3@��!WO�!?v�w�~�@��Nt۠ٿX�b�v��@��q|�3@��!WO�!?v�w�~�@��Nt۠ٿX�b�v��@��q|�3@��!WO�!?v�w�~�@��Nt۠ٿX�b�v��@��q|�3@��!WO�!?v�w�~�@���ٿ���c�@i��J:�3@�4cw�!?ܬ���@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�jf �ٿ8}b���@}�^E�.4@�t����!?	�n�i�@�)�x�ٿ���&M�@H�:S#G4@�3p���!?{�O�֌�@�)�x�ٿ���&M�@H�:S#G4@�3p���!?{�O�֌�@~"x�7�ٿCݗ����@�Ì�4@ٗd8ΐ!?��\	��@~"x�7�ٿCݗ����@�Ì�4@ٗd8ΐ!?��\	��@~"x�7�ٿCݗ����@�Ì�4@ٗd8ΐ!?��\	��@~"x�7�ٿCݗ����@�Ì�4@ٗd8ΐ!?��\	��@~"x�7�ٿCݗ����@�Ì�4@ٗd8ΐ!?��\	��@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@�(�ٿ��l˻�@s�"�3@3Ψ�e�!?V'*0�ە@1<�ٿ�j�5���@���G�3@L� _4�!?�u�3�@1<�ٿ�j�5���@���G�3@L� _4�!?�u�3�@1<�ٿ�j�5���@���G�3@L� _4�!?�u�3�@1<�ٿ�j�5���@���G�3@L� _4�!?�u�3�@��?��ٿ��XI��@�;�#�4@�Ikg�!?yz�}�ѕ@��?��ٿ��XI��@�;�#�4@�Ikg�!?yz�}�ѕ@��?��ٿ��XI��@�;�#�4@�Ikg�!?yz�}�ѕ@��?��ٿ��XI��@�;�#�4@�Ikg�!?yz�}�ѕ@fK���ٿ��L���@��<t.4@� ;��!?�u���@��cAH�ٿ�D6�@�'�	4@���a�!?D����-�@��cAH�ٿ�D6�@�'�	4@���a�!?D����-�@��cAH�ٿ�D6�@�'�	4@���a�!?D����-�@���L�ٿ�5�êQ�@��iB 4@��k�m�!?���0P
�@���L�ٿ�5�êQ�@��iB 4@��k�m�!?���0P
�@���L�ٿ�5�êQ�@��iB 4@��k�m�!?���0P
�@���L�ٿ�5�êQ�@��iB 4@��k�m�!?���0P
�@���L�ٿ�5�êQ�@��iB 4@��k�m�!?���0P
�@�Ýa6�ٿ��u\LN�@��צ�4@��ϋG�!?A�R���@�Ýa6�ٿ��u\LN�@��צ�4@��ϋG�!?A�R���@�Ýa6�ٿ��u\LN�@��צ�4@��ϋG�!?A�R���@�Ýa6�ٿ��u\LN�@��צ�4@��ϋG�!?A�R���@�Ýa6�ٿ��u\LN�@��צ�4@��ϋG�!?A�R���@=��Sܟٿ`{�C�j�@���44@Zn0;b�!?��ˀȰ�@=��Sܟٿ`{�C�j�@���44@Zn0;b�!?��ˀȰ�@�K�Cn�ٿ�_�Ir��@BxL2!4@�ɒ���!?�ӹK��@Ф�ߝٿ��6t��@|��O|4@�N����!?�0(/��@Ф�ߝٿ��6t��@|��O|4@�N����!?�0(/��@�	� ��ٿ51��ۏ�@H�u�64@�_�B�!?�[̑P�@�	� ��ٿ51��ۏ�@H�u�64@�_�B�!?�[̑P�@�	� ��ٿ51��ۏ�@H�u�64@�_�B�!?�[̑P�@b�:�ٿ#@M'v��@u�s4@os�ml�!?��J� ˕@b�:�ٿ#@M'v��@u�s4@os�ml�!?��J� ˕@b�:�ٿ#@M'v��@u�s4@os�ml�!?��J� ˕@b�:�ٿ#@M'v��@u�s4@os�ml�!?��J� ˕@b�:�ٿ#@M'v��@u�s4@os�ml�!?��J� ˕@��+���ٿ�uL�5�@��z��K4@8�A��!?���@=�
���ٿ��ݰM�@+P�_LU4@�WS�!?q��0��@=�
���ٿ��ݰM�@+P�_LU4@�WS�!?q��0��@=�
���ٿ��ݰM�@+P�_LU4@�WS�!?q��0��@nu��J�ٿV�|hN�@��B��4@��=�!?131Hoؕ@nu��J�ٿV�|hN�@��B��4@��=�!?131Hoؕ@�㈞�ٿ �U����@�'����3@�.��E�!?��5�檕@���ٿ2�?��@�k�G��3@����!?0��!��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@*
�Jo�ٿ��Ar�@�X���3@��=�!?W@vI��@E$b�~�ٿ��a�i�@�!�L4@k����!?�^Y���@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@���i�ٿ�I"80��@B�͐24@B�%�J�!??�j����@=&�ԙ�ٿcOY���@�KXP�4@:o�k��!?�藨�@=&�ԙ�ٿcOY���@�KXP�4@:o�k��!?�藨�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@Bw��ٿ0WW׆��@�p�7	N4@��w}�!?�)�^�@5��×ٿ�-����@��3B`4@�HK\G�!?��Հ��@5��×ٿ�-����@��3B`4@�HK\G�!?��Հ��@���;��ٿp��{t�@o*��p	4@hy�*�!?)��u>�@���;��ٿp��{t�@o*��p	4@hy�*�!?)��u>�@���;��ٿp��{t�@o*��p	4@hy�*�!?)��u>�@�FكK�ٿc�z�T�@�#f�4@X6��/�!?F���w�@��=���ٿ�O�4��@Ó�r�`4@�l�Z�!?g���ו�@�/�Ǌ�ٿ�r����@39
��j4@P�/��!?!ԡ,hl�@�/�Ǌ�ٿ�r����@39
��j4@P�/��!?!ԡ,hl�@�/�Ǌ�ٿ�r����@39
��j4@P�/��!?!ԡ,hl�@�ݰtʧٿp�BUC�@$���14@d�9���!?�������@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@d[Qyi�ٿ�*�b��@ŬI5�4@�17$U�!?����@�p��y�ٿN>�S=��@�)�pV4@�D��/�!?ϒ���E�@:�;��ٿR��_p��@3 ���a4@I���!�!?�22�}�@� ϛ*�ٿ�\��@�����=4@D��7�!?��"�ۖ@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@��
�,�ٿ>�#���@��ZLR4@�>>�!?����@][���ٿ<6�_��@R���x]4@�;i/F�!?�q��^��@][���ٿ<6�_��@R���x]4@�;i/F�!?�q��^��@][���ٿ<6�_��@R���x]4@�;i/F�!?�q��^��@][���ٿ<6�_��@R���x]4@�;i/F�!?�q��^��@�L�N�ٿ"~d���@ٽH�4@����_�!?C�ʦ`�@�L�N�ٿ"~d���@ٽH�4@����_�!?C�ʦ`�@�L�N�ٿ"~d���@ٽH�4@����_�!?C�ʦ`�@�L�N�ٿ"~d���@ٽH�4@����_�!?C�ʦ`�@3 �'�ٿ�S�����@������3@��w�!?䜎����@3 �'�ٿ�S�����@������3@��w�!?䜎����@3 �'�ٿ�S�����@������3@��w�!?䜎����@U��2ٙٿ.N���<�@k�p8L�3@艏 A�!?pY:����@U��2ٙٿ.N���<�@k�p8L�3@艏 A�!?pY:����@U��2ٙٿ.N���<�@k�p8L�3@艏 A�!?pY:����@U��2ٙٿ.N���<�@k�p8L�3@艏 A�!?pY:����@U��2ٙٿ.N���<�@k�p8L�3@艏 A�!?pY:����@�Y/h�ٿ)���J��@�*��3@u��^�!?�b��v�@�q7���ٿ�炭���@����,4@���	�!?���b��@�q7���ٿ�炭���@����,4@���	�!?���b��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@ AM��ٿj.k;�@�z�%��3@L�q|g�!?|�E~��@��R���ٿড6~a�@CXh'h�3@��eؚ�!?m��i>�@ �>�ٿ)'>����@�P�4@�3C���!?��.��@ �>�ٿ)'>����@�P�4@�3C���!?��.��@ �>�ٿ)'>����@�P�4@�3C���!?��.��@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@����ٿ2]He�^�@ϡ�B4@��k��!?�r&YU�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@�����ٿn���@)#O��N4@j����!?5�`f(�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@V�Z�ڙٿ�wr'��@`�RG4@�,.�!?���#9w�@�t�b��ٿ�����@f�E��#4@&��䧐!?�n�vt�@��%��ٿF�)����@'�L�[4@��	H��!?[��J5��@��%��ٿF�)����@'�L�[4@��	H��!?[��J5��@����N�ٿ�K/�V��@ok 7�,4@���k�!?%��,�g�@����N�ٿ�K/�V��@ok 7�,4@���k�!?%��,�g�@�+��ٿt*h��@V�K�C4@�?��s�!?s���
��@�+��ٿt*h��@V�K�C4@�?��s�!?s���
��@�+��ٿt*h��@V�K�C4@�?��s�!?s���
��@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@˧��Ġٿ�ޝ���@��@Q4@�$+�!?�^`�Ǖ@��f�ٿv� 4���@g�?�}4@�Rd�!?�m4�@��f�ٿv� 4���@g�?�}4@�Rd�!?�m4�@83Qۛٿ�ߪ�c�@�D���4@�G�tv�!?�Y,A��@83Qۛٿ�ߪ�c�@�D���4@�G�tv�!?�Y,A��@83Qۛٿ�ߪ�c�@�D���4@�G�tv�!?�Y,A��@83Qۛٿ�ߪ�c�@�D���4@�G�tv�!?�Y,A��@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@�Z���ٿ�
���@X?R�a4@�)W��!?_ϭ2���@��D+�ٿ�^?�~�@�GSd4@{�axs�!?2Dp\��@��D+�ٿ�^?�~�@�GSd4@{�axs�!?2Dp\��@��D+�ٿ�^?�~�@�GSd4@{�axs�!?2Dp\��@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@�=�=�ٿO��#��@�)�4@	���!?��:0C�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@ot�"A�ٿ�6QB��@@�J�
4@\0

��!?&0�k?0�@���m�ٿ8����@���0�3@�AX`�!?��(�p"�@���m�ٿ8����@���0�3@�AX`�!?��(�p"�@���m�ٿ8����@���0�3@�AX`�!?��(�p"�@w�"P�ٿ��W;�/�@B��M�4@��[�!?�F	���@8��P�ٿH�NZK��@���4@W�w�!?.H���@8��P�ٿH�NZK��@���4@W�w�!?.H���@8��P�ٿH�NZK��@���4@W�w�!?.H���@8��P�ٿH�NZK��@���4@W�w�!?.H���@8��P�ٿH�NZK��@���4@W�w�!?.H���@_{�R�ٿ�h�v��@T��a4@^�=W�!?ܺ[���@W3�&��ٿ-s�C4!�@+,�?4@��`�͐!?�Xu|Y�@tE�W�ٿ&���,�@�R�8�3@v�݁ѐ!?��3��@��po �ٿ��F܇�@��b4@m�p�/�!?Z�v�@��po �ٿ��F܇�@��b4@m�p�/�!?Z�v�@��po �ٿ��F܇�@��b4@m�p�/�!?Z�v�@��po �ٿ��F܇�@��b4@m�p�/�!?Z�v�@Co�?a�ٿ�O�[8�@#�?�4@yč��!?��w���@Co�?a�ٿ�O�[8�@#�?�4@yč��!?��w���@Co�?a�ٿ�O�[8�@#�?�4@yč��!?��w���@Co�?a�ٿ�O�[8�@#�?�4@yč��!?��w���@탗�ٛٿ�p�W�@�Zˆֶ3@�yȞ��!?%z����@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@�Ux+�ٿ2acl#��@!�"��3@�.����!?	�]��@pV��~�ٿYu0K���@�X���3@�
9���!?���Ul��@pV��~�ٿYu0K���@�X���3@�
9���!?���Ul��@ph�ٿG�nJ��@�����3@1²�!?ۑϞ�ɕ@!0ޗt�ٿc`��'e�@ �M��3@�C��x�!?�)*X�˕@!0ޗt�ٿc`��'e�@ �M��3@�C��x�!?�)*X�˕@!0ޗt�ٿc`��'e�@ �M��3@�C��x�!?�)*X�˕@R"�U��ٿV��$>�@�����3@��D�R�!?��^˕@R"�U��ٿV��$>�@�����3@��D�R�!?��^˕@L�ǋ2�ٿ��S-o��@!a��v4@���O�!?�AX�c�@L�ǋ2�ٿ��S-o��@!a��v4@���O�!?�AX�c�@L�ǋ2�ٿ��S-o��@!a��v4@���O�!?�AX�c�@L�ǋ2�ٿ��S-o��@!a��v4@���O�!?�AX�c�@L�ǋ2�ٿ��S-o��@!a��v4@���O�!?�AX�c�@BAA1�ٿ�6�&!v�@����<4@��m�!?���}��@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@pV��~�ٿ�$�d��@�[4@�J<#�!?��'0�)�@�X���ٿV<g����@̈́�ݞ�3@6��b�!?+���o�@�X���ٿV<g����@̈́�ݞ�3@6��b�!?+���o�@�X���ٿV<g����@̈́�ݞ�3@6��b�!?+���o�@�X���ٿV<g����@̈́�ݞ�3@6��b�!?+���o�@��y��ٿ��FUzC�@��a�4@ �&7�!?���W1�@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@�&6 �ٿu����@��v�54@"�W]>�!?��@yX��ٿ���rb�@d����3@�bǄ�!?ϨyDw�@yX��ٿ���rb�@d����3@�bǄ�!?ϨyDw�@SAwr��ٿ~K
����@�3h�R4@�u��r�!?u�
����@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�xyF��ٿl\�V�@�i]�V4@���-�!?�'�iǕ@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@�����ٿ���t|^�@�߁>�4@�d%1�!?�m/�7	�@��H�ٿD�,x�@�v��3?4@�
�!?�RO�$�@%O�ʘٿsup.�@�b���3@Y�!��!?����,�@%O�ʘٿsup.�@�b���3@Y�!��!?����,�@&R�#�ٿ�[ �@��^�4@s�'*�!?�(-G��@&R�#�ٿ�[ �@��^�4@s�'*�!?�(-G��@&R�#�ٿ�[ �@��^�4@s�'*�!?�(-G��@�U�!�ٿ���O�@��q�3@�#�D�!?�5Rѕ@�U�!�ٿ���O�@��q�3@�#�D�!?�5Rѕ@h� ᄙٿ��L�g��@͌7�Q4@�����!?I��-���@h� ᄙٿ��L�g��@͌7�Q4@�����!?I��-���@j�ҙٿE%�RdO�@��<�3@��6,�!?yTm}�}�@j�ҙٿE%�RdO�@��<�3@��6,�!?yTm}�}�@j�ҙٿE%�RdO�@��<�3@��6,�!?yTm}�}�@j�ҙٿE%�RdO�@��<�3@��6,�!?yTm}�}�@I��x�ٿ��;m	��@�=�z�3@�f;�k�!?Rk(�=�@I��x�ٿ��;m	��@�=�z�3@�f;�k�!?Rk(�=�@I��x�ٿ��;m	��@�=�z�3@�f;�k�!?Rk(�=�@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@��da��ٿ�������@��L��/4@h�W$��!?,��瓕@�/��ٿ.i"��@������3@7�&�Q�!?��+!;H�@�O>C4�ٿ�����@G4��O�3@�4�x�!?�}�>C;�@Og�F�ٿ�d�K�@�D�L"4@k����!?Dy<��V�@Og�F�ٿ�d�K�@�D�L"4@k����!?Dy<��V�@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�Qvpj�ٿ��� ��@׊M�44@�����!?�t����@�GY�؛ٿ��b?��@�4��M4@�Y��!?����M��@�GY�؛ٿ��b?��@�4��M4@�Y��!?����M��@�� �ٿ�\;5���@9����3@d��F�!?��
�:Y�@�� �ٿ�\;5���@9����3@d��F�!?��
�:Y�@�� �ٿ�\;5���@9����3@d��F�!?��
�:Y�@�� �ٿ�\;5���@9����3@d��F�!?��
�:Y�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@��To�ٿ�Y��(�@�Q��3@��qy�!?FɪG�L�@9��Z��ٿ������@��@4@�f��'�!?�8^�^ߕ@9��Z��ٿ������@��@4@�f��'�!?�8^�^ߕ@pv�8�ٿ]ġF_I�@��Ch4@X���8�!?o����@v�p��ٿ����/�@�A54@�Q�ߏ!?��etz�@����ٿ{�����@~�Qf�3@��P���!?�6D���@����ٿ{�����@~�Qf�3@��P���!?�6D���@9S[S��ٿ�+����@S=�L84@���V�!?�#<���@9S[S��ٿ�+����@S=�L84@���V�!?�#<���@9S[S��ٿ�+����@S=�L84@���V�!?�#<���@9S[S��ٿ�+����@S=�L84@���V�!?�#<���@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@�T��i�ٿ6;ɴ@�@�>�J��3@�b��r�!?Ҏ�dM�@8���I�ٿG�m|�@,�/�4@���)�!?ޑ!wP��@8���I�ٿG�m|�@,�/�4@���)�!?ޑ!wP��@������ٿ�#�4��@W��M�4@����!?�_v���@������ٿ�#�4��@W��M�4@����!?�_v���@������ٿ�#�4��@W��M�4@����!?�_v���@oU	�D�ٿ(:{8���@��!�j!4@��$���!?�J��v�@�z���ٿ�m`_v)�@L��S@4@����Ӑ!?8�/�0��@�z���ٿ�m`_v)�@L��S@4@����Ӑ!?8�/�0��@,�mv��ٿm.��Q�@t
��u4@x�W��!?� JE�@,�mv��ٿm.��Q�@t
��u4@x�W��!?� JE�@,�mv��ٿm.��Q�@t
��u4@x�W��!?� JE�@,�mv��ٿm.��Q�@t
��u4@x�W��!?� JE�@,�mv��ٿm.��Q�@t
��u4@x�W��!?� JE�@���l��ٿim�m��@�Goʫ`4@˱�L��!?!8_}4D�@���l��ٿim�m��@�Goʫ`4@˱�L��!?!8_}4D�@�̹�C�ٿ��mGFN�@kM�94@GJ�	�!?>bHb�@qx4q�ٿ��"0z�@a���3@C�ֹ��!?
�Iٕ@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@aj|��ٿ<0��>��@�y����3@5�[��!?@�on�@��o�ٿ���b�C�@n�� �3@�i_�!?���+R�@��o�ٿ���b�C�@n�� �3@�i_�!?���+R�@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@I�p��ٿiߋ�#u�@��<4@d�ʒ��!?S�����@�SX�n�ٿ}��m��@SA�4@�WJ�!?���?�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@H� %�ٿϩKh@�@��1`4[4@�
�R�!?3���:�@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@"���ٿ�<_h9��@��s� 4@-�qU!�!?�3N#��@h�7�ٿ�,�hWG�@I<�H3�3@�1�9[�!?9���]�@h�7�ٿ�,�hWG�@I<�H3�3@�1�9[�!?9���]�@h�7�ٿ�,�hWG�@I<�H3�3@�1�9[�!?9���]�@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@���Mͤٿ]f�@h�9�t4@k2�Ѡ�!?W[�P��@X>��ۤٿ�<U �@����4@.�/�!?(�,�ٕ@X>��ۤٿ�<U �@����4@.�/�!?(�,�ٕ@X>��ۤٿ�<U �@����4@.�/�!?(�,�ٕ@X>��ۤٿ�<U �@����4@.�/�!?(�,�ٕ@X>��ۤٿ�<U �@����4@.�/�!?(�,�ٕ@D^���ٿ�A��\u�@�,\�3@̉�Gh�!?��m�^�@D^���ٿ�A��\u�@�,\�3@̉�Gh�!?��m�^�@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@]V��ٿ�"�%�@���0�3@Y9��l�!?$��і@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@��kA�ٿ�p�XO�@˴:��4@R�Jʐ!?�S&h&X�@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@�1�1�ٿ~ԤG�@sD�[�3@��'���!?}A�v��@n��I՛ٿX�V��'�@lT���3@�*Zz��!?�|�̕@n��I՛ٿX�V��'�@lT���3@�*Zz��!?�|�̕@n��I՛ٿX�V��'�@lT���3@�*Zz��!?�|�̕@n��I՛ٿX�V��'�@lT���3@�*Zz��!?�|�̕@n��I՛ٿX�V��'�@lT���3@�*Zz��!?�|�̕@��Lη�ٿ\D���@��N�4@mj�`ϐ!?�K���@��Lη�ٿ\D���@��N�4@mj�`ϐ!?�K���@�%Y`�ٿ����6�@L���%4@�c��!?��kf���@�%Y`�ٿ����6�@L���%4@�c��!?��kf���@m��t�ٿ���X��@�i��44@rȱ��!?� ��@m��t�ٿ���X��@�i��44@rȱ��!?� ��@m��t�ٿ���X��@�i��44@rȱ��!?� ��@m��t�ٿ���X��@�i��44@rȱ��!?� ��@m��t�ٿ���X��@�i��44@rȱ��!?� ��@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@�*�aG�ٿ
�.����@���@�4@!��p��!?�'��Е@㏮���ٿ|��X�R�@��5��3@;��!?�X����@㏮���ٿ|��X�R�@��5��3@;��!?�X����@-sr�ٿ�1Kb���@�Ag�<4@ge�5�!?O �,�#�@-sr�ٿ�1Kb���@�Ag�<4@ge�5�!?O �,�#�@�)�I�ٿ� 5���@���DH4@)P���!?�.���@�)�I�ٿ� 5���@���DH4@)P���!?�.���@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@K���u�ٿ��J���@���"4@����!?�=Y�=ޕ@&�sh��ٿK<�`<�@r��,��3@K�^�)�!?],\����@&�sh��ٿK<�`<�@r��,��3@K�^�)�!?],\����@&�sh��ٿK<�`<�@r��,��3@K�^�)�!?],\����@x��եٿf���Y��@Ы�q�-4@9�1J!�!?�5�9 ��@x��եٿf���Y��@Ы�q�-4@9�1J!�!?�5�9 ��@p�^�ٿv��Ŗ	�@�ֱ4 4@4�$ҏ!?�$3'Z5�@p�^�ٿv��Ŗ	�@�ֱ4 4@4�$ҏ!?�$3'Z5�@p�^�ٿv��Ŗ	�@�ֱ4 4@4�$ҏ!?�$3'Z5�@��K�ٿ$U���@9n���4@�K�!?R0�LRŕ@��K�ٿ$U���@9n���4@�K�!?R0�LRŕ@��K�ٿ$U���@9n���4@�K�!?R0�LRŕ@��K�ٿ$U���@9n���4@�K�!?R0�LRŕ@��K�ٿ$U���@9n���4@�K�!?R0�LRŕ@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@��]��ٿ���S��@��U�pM4@EhgJ�!?g/	���@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@<h�:ȟٿ�L?ޭ�@�ʓ�fm4@\�Z�!?���|6�@�J �ٿ�2Db��@bN��?4@sb�=8�!?j����c�@�J �ٿ�2Db��@bN��?4@sb�=8�!?j����c�@�J �ٿ�2Db��@bN��?4@sb�=8�!?j����c�@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@ŏ�(��ٿK⿋��@���^B(4@�!��(�!?2sa��@=���ٿ?3�����@��]U5+4@-��!�!?q�1�@=���ٿ?3�����@��]U5+4@-��!�!?q�1�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@]'�/�ٿT��%��@v��54@z�9ʚ�!?%[�Ru�@�$B�ٿ
x��a<�@�����04@]�e���!?�$���@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@�ô��ٿ�by�>�@�a���4@��i��!?��y@�+�@5*H�-�ٿ�h��0��@Ք�
]4@wRv�!?��U�;Օ@GB��ٿ��Z`�@ur�G�_4@/`�{�!?wƹ5���@GB��ٿ��Z`�@ur�G�_4@/`�{�!?wƹ5���@GB��ٿ��Z`�@ur�G�_4@/`�{�!?wƹ5���@GB��ٿ��Z`�@ur�G�_4@/`�{�!?wƹ5���@0,� �ٿ	x5�_��@R  ��4@�ujh�!?����$~�@0,� �ٿ	x5�_��@R  ��4@�ujh�!?����$~�@0,� �ٿ	x5�_��@R  ��4@�ujh�!?����$~�@0,� �ٿ	x5�_��@R  ��4@�ujh�!?����$~�@
e���ٿ�ع���@�X�2#�4@肋x�!?�^#��=�@
e���ٿ�ع���@�X�2#�4@肋x�!?�^#��=�@��2�ٿ�kW-��@g���r4@��`v`�!?�7��C"�@��2�ٿ�kW-��@g���r4@��`v`�!?�7��C"�@��2�ٿ�kW-��@g���r4@��`v`�!?�7��C"�@��2�ٿ�kW-��@g���r4@��`v`�!?�7��C"�@��2�ٿ�kW-��@g���r4@��`v`�!?�7��C"�@WQ���ٿ�$�����@X�A`�,4@Q\kM�!?�s���#�@WQ���ٿ�$�����@X�A`�,4@Q\kM�!?�s���#�@WQ���ٿ�$�����@X�A`�,4@Q\kM�!?�s���#�@WQ���ٿ�$�����@X�A`�,4@Q\kM�!?�s���#�@WQ���ٿ�$�����@X�A`�,4@Q\kM�!?�s���#�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@~��ݞٿ(Q�7�6�@H�z�vr4@��X��!?U%���}�@9��۳�ٿ-����@ }bг54@�4����!?D����@9��۳�ٿ-����@ }bг54@�4����!?D����@9��۳�ٿ-����@ }bг54@�4����!?D����@�C��ٿ^4轥��@)<�;��3@��œ�!?
B��2�@�C��ٿ^4轥��@)<�;��3@��œ�!?
B��2�@�C��ٿ^4轥��@)<�;��3@��œ�!?
B��2�@4��ٿ�&����@]�ʔN+4@G�X�{�!?|[	�Sp�@4��ٿ�&����@]�ʔN+4@G�X�{�!?|[	�Sp�@4��ٿ�&����@]�ʔN+4@G�X�{�!?|[	�Sp�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@��fCݟٿz��rl�@�^�<'/4@������!?���`#�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@�1;�Оٿ-��v��@�����3@�1c�J�!?f4�@J��զ�ٿ�ڈ`��@PQK
4@��E�!?�ً@�=�@J��զ�ٿ�ڈ`��@PQK
4@��E�!?�ً@�=�@J��զ�ٿ�ڈ`��@PQK
4@��E�!?�ً@�=�@�uՊ,�ٿ�s~����@��1��4@AYy��!?��L�ؕ@�uՊ,�ٿ�s~����@��1��4@AYy��!?��L�ؕ@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@	U"��ٿ��~+*��@��'\�4@"=�m"�!?��q�?��@�[?l'�ٿ�_�ޔ��@�~e�4@��#�#�!?6 ��a��@�[?l'�ٿ�_�ޔ��@�~e�4@��#�#�!?6 ��a��@�[?l'�ٿ�_�ޔ��@�~e�4@��#�#�!?6 ��a��@�[?l'�ٿ�_�ޔ��@�~e�4@��#�#�!?6 ��a��@�[?l'�ٿ�_�ޔ��@�~e�4@��#�#�!?6 ��a��@Ѩ{;!�ٿ�\<kfz�@��14@�ߛ���!?��f��_�@Ѩ{;!�ٿ�\<kfz�@��14@�ߛ���!?��f��_�@Ѩ{;!�ٿ�\<kfz�@��14@�ߛ���!?��f��_�@�G %�ٿ��qn.~�@�0I
[4@���(�!?�r�D�h�@~+�}�ٿA��
���@���5��3@*���ҏ!?��� ���@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@k�;���ٿ�P-ȑ��@��%�k�3@�X�<ݏ!?�d2K�@���C�ٿ��ۑ ��@e�$�3@��C���!?*>/i�@���C�ٿ��ۑ ��@e�$�3@��C���!?*>/i�@�6�?��ٿ�9�����@��b�4@ݔmӏ!?�1�"lq�@Z��А�ٿt&���@�_��{`4@I�ƴ%�!? .�#N�@Z��А�ٿt&���@�_��{`4@I�ƴ%�!? .�#N�@Z��А�ٿt&���@�_��{`4@I�ƴ%�!? .�#N�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@�q�<�ٿ�c>�<�@�=E�V�3@�u�!?�ʆ�E�@z�ʋ��ٿ��'��@��.���3@�����!?�S5��@z�ʋ��ٿ��'��@��.���3@�����!?�S5��@z�ʋ��ٿ��'��@��.���3@�����!?�S5��@z�ʋ��ٿ��'��@��.���3@�����!?�S5��@z�ʋ��ٿ��'��@��.���3@�����!?�S5��@�u�nL�ٿ��cR��@	���24@JmM<7�!?��r�鋕@�u�nL�ٿ��cR��@	���24@JmM<7�!?��r�鋕@�~>�ٿ�܂�T��@���]4@�Z]K�!?>1b�˕@��a��ٿ����2��@���_04@��-��!?�uWީԕ@��a��ٿ����2��@���_04@��-��!?�uWީԕ@��a��ٿ����2��@���_04@��-��!?�uWީԕ@��a��ٿ����2��@���_04@��-��!?�uWީԕ@��a��ٿ����2��@���_04@��-��!?�uWީԕ@�%~���ٿ�}���@�c��Q<4@���q�!?9`~�@�%~���ٿ�}���@�c��Q<4@���q�!?9`~�@�%~���ٿ�}���@�c��Q<4@���q�!?9`~�@n��=I�ٿ�NjI���@����)�3@����`�!?,<So�@n��=I�ٿ�NjI���@����)�3@����`�!?,<So�@n��=I�ٿ�NjI���@����)�3@����`�!?,<So�@n��=I�ٿ�NjI���@����)�3@����`�!?,<So�@n��=I�ٿ�NjI���@����)�3@����`�!?,<So�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@��O��ٿ� �,@�@��tf(4@�Ly�!?K,�S1�@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@ܞ�>��ٿ���|1��@�8aLY4@�E���!?ͼ�9��@��s�ٿ��o���@�(qd�54@K|CaJ�!?���]'�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@�>��M�ٿ�ZHP��@z u� 4@$�iO��!?c[� �
�@���VR�ٿ���g&�@1�A�R4@7�{{�!?�T�'��@���VR�ٿ���g&�@1�A�R4@7�{{�!?�T�'��@���VR�ٿ���g&�@1�A�R4@7�{{�!?�T�'��@���VR�ٿ���g&�@1�A�R4@7�{{�!?�T�'��@0�pЧ�ٿ_'�dRM�@�hS�@4@?,r�A�!?m�C�ѕ@0�pЧ�ٿ_'�dRM�@�hS�@4@?,r�A�!?m�C�ѕ@0�pЧ�ٿ_'�dRM�@�hS�@4@?,r�A�!?m�C�ѕ@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�<\�ٿcX�M��@���+74@eoe阐!?E��Y�@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@�y��ٿ��Xd���@5 	�/4@�{L�2�!?�<��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@-'��6�ٿ���}�@߆c[�-4@�3�|�!?/0\5��@/��*r�ٿ۞��}��@k]�W;�3@����%�!?��!3�@/��*r�ٿ۞��}��@k]�W;�3@����%�!?��!3�@P��e�ٿ@�$���@���4@���4�!?̃�s0J�@P��e�ٿ@�$���@���4@���4�!?̃�s0J�@P��e�ٿ@�$���@���4@���4�!?̃�s0J�@P��e�ٿ@�$���@���4@���4�!?̃�s0J�@7!p��ٿU&7\�d�@d<,���3@�AZx�!?G�aVl[�@7!p��ٿU&7\�d�@d<,���3@�AZx�!?G�aVl[�@7!p��ٿU&7\�d�@d<,���3@�AZx�!?G�aVl[�@7!p��ٿU&7\�d�@d<,���3@�AZx�!?G�aVl[�@�/�<�ٿHs����@�D��K�3@|(�G�!?G}���E�@�/�<�ٿHs����@�D��K�3@|(�G�!?G}���E�@�/�<�ٿHs����@�D��K�3@|(�G�!?G}���E�@��ܪ��ٿx_ ���@����3@���|Z�!?rL)�ǟ�@��ܪ��ٿx_ ���@����3@���|Z�!?rL)�ǟ�@��ܪ��ٿx_ ���@����3@���|Z�!?rL)�ǟ�@�6/�ٿ3�����@��=4@yD	���!?\m�v�Y�@�6/�ٿ3�����@��=4@yD	���!?\m�v�Y�@�6/�ٿ3�����@��=4@yD	���!?\m�v�Y�@�6/�ٿ3�����@��=4@yD	���!?\m�v�Y�@�6/�ٿ3�����@��=4@yD	���!?\m�v�Y�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@y��b?�ٿBa�bQ�@���
�3@��^��!?I�^�J�@BЍf��ٿ[�~�0�@�61�^�3@,m��q�!?�(_���@�sJ+�ٿd8bJ\)�@��7�4@s돨��!?d��l�r�@�sJ+�ٿd8bJ\)�@��7�4@s돨��!?d��l�r�@�R[>�ٿ�ݢb��@�y[�4@�%���!?Gt�H�@�\�yq�ٿ��ʹ��@�=*�3@��G�!?���
�H�@�\�yq�ٿ��ʹ��@�=*�3@��G�!?���
�H�@�\�yq�ٿ��ʹ��@�=*�3@��G�!?���
�H�@�\�yq�ٿ��ʹ��@�=*�3@��G�!?���
�H�@�Q�.�ٿ=�ZQH��@����3@j���|�!?��M���@Ħa��ٿ�^��(t�@�%���3@��A�!?AHA�@F�\%�ٿd�1c��@L:&� 4@�]���!?>�f���@F�\%�ٿd�1c��@L:&� 4@�]���!?>�f���@F�\%�ٿd�1c��@L:&� 4@�]���!?>�f���@F�\%�ٿd�1c��@L:&� 4@�]���!?>�f���@F�\%�ٿd�1c��@L:&� 4@�]���!?>�f���@y!?͟ٿV��ɼ�@�H��3@]跣�!?^l^��h�@y!?͟ٿV��ɼ�@�H��3@]跣�!?^l^��h�@y!?͟ٿV��ɼ�@�H��3@]跣�!?^l^��h�@1�Z��ٿǊs���@*��*�3@څ0ܨ�!?ٞ�z���@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@H���ٿ����T�@�,��H�3@������!?6�m2�ڕ@�sQ�Ϟٿ�����e�@.�P4@�}񺗐!?v�#��@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@��k莜ٿ5��v��@]�?0��3@:A��j�!?N:����@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@5�M���ٿS���3��@d�F�34@eu�4�!?��jQҕ@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@���ٿ[������@�0uaF�3@��<z+�!?���@W�E�ٿ|�����@���1(4@�@���!?�FZH��@W�E�ٿ|�����@���1(4@�@���!?�FZH��@W�E�ٿ|�����@���1(4@�@���!?�FZH��@W�E�ٿ|�����@���1(4@�@���!?�FZH��@W�E�ٿ|�����@���1(4@�@���!?�FZH��@j�T��ٿ���K��@����Y4@j����!?lh�����@j�T��ٿ���K��@����Y4@j����!?lh�����@ߐl�;�ٿ�q����@M�#�4@ɉ	�V�!?0txR�@ߐl�;�ٿ�q����@M�#�4@ɉ	�V�!?0txR�@ߐl�;�ٿ�q����@M�#�4@ɉ	�V�!?0txR�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@�Ai�ٿ[J�=���@�/��+4@�E��P�!?�Q��'�@Ë���ٿetڇƃ�@*�q�4@�F�8�!??n�c�S�@Ë���ٿetڇƃ�@*�q�4@�F�8�!??n�c�S�@��	j�ٿi�-{�@uW�[�3@j��(�!?��(�g)�@��oj�ٿa=4�\�@���S��3@���7�!?����vr�@��oj�ٿa=4�\�@���S��3@���7�!?����vr�@9j@��ٿӰ}fJ�@��)>�3@	�1@�!?�*�&)�@9j@��ٿӰ}fJ�@��)>�3@	�1@�!?�*�&)�@9j@��ٿӰ}fJ�@��)>�3@	�1@�!?�*�&)�@��v�ٿ�*g���@�h�ao4@�X��)�!?��<H��@��v�ٿ�*g���@�h�ao4@�X��)�!?��<H��@��v�ٿ�*g���@�h�ao4@�X��)�!?��<H��@'��G��ٿ�mP�@��5!�]4@i����!?._�ϕ@'��G��ٿ�mP�@��5!�]4@i����!?._�ϕ@�b6V�ٿ��3���@�O"�;4@P�V�!?q\����@�b6V�ٿ��3���@�O"�;4@P�V�!?q\����@�b6V�ٿ��3���@�O"�;4@P�V�!?q\����@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@o%FR`�ٿ��(��^�@o1���D4@dOV�!?���qf�@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@��|t�ٿkIy,�n�@�r�>4@�b�U��!?��S����@lC�N�ٿ�
n3%��@r9�`4@|&\i��!?�N6�͕@lC�N�ٿ�
n3%��@r9�`4@|&\i��!?�N6�͕@lC�N�ٿ�
n3%��@r9�`4@|&\i��!?�N6�͕@lC�N�ٿ�
n3%��@r9�`4@|&\i��!?�N6�͕@��,;��ٿ���h�@u*br4@�h��!?QQ����@���g�ٿa�HN3a�@�3L��?4@�kR{�!?e�����@���g�ٿa�HN3a�@�3L��?4@�kR{�!?e�����@���g�ٿa�HN3a�@�3L��?4@�kR{�!?e�����@tazq�ٿ���3_�@���4@����F�!?�"�2�@tazq�ٿ���3_�@���4@����F�!?�"�2�@tazq�ٿ���3_�@���4@����F�!?�"�2�@tazq�ٿ���3_�@���4@����F�!?�"�2�@tazq�ٿ���3_�@���4@����F�!?�"�2�@8�<���ٿ�#1��(�@�)�YT�3@Q�i:i�!?�պW��@8�<���ٿ�#1��(�@�)�YT�3@Q�i:i�!?�պW��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��S3��ٿ�כ�_,�@���z��3@t��<�!?��A_4��@��'4�ٿ�ə9d�@6`*L�3@���I�!?�zj�."�@��'4�ٿ�ə9d�@6`*L�3@���I�!?�zj�."�@��'4�ٿ�ə9d�@6`*L�3@���I�!?�zj�."�@Ǥ��ٿ�����@3����3@7Ձ�!?F'g&֕@H�
��ٿ��Q�! �@����4@l�L��!?"�.��o�@l��f7�ٿ ��LR�@����3@4��Ge�!?.����S�@P�o$c�ٿD����@��m:��3@t]��!?+��Ne��@P�o$c�ٿD����@��m:��3@t]��!?+��Ne��@P�o$c�ٿD����@��m:��3@t]��!?+��Ne��@��J)6�ٿ��28"��@V},IH4@��F��!?@$C~ٖ@���|�ٿ�k���@�W�.9t4@t�aTZ�!?��Fe~�@���|�ٿ�k���@�W�.9t4@t�aTZ�!?��Fe~�@���|�ٿ�k���@�W�.9t4@t�aTZ�!?��Fe~�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@����ٿ#ؽ����@{Ic��24@VϡÐ!?�|�LQ?�@��%�ٿ�����I�@ބZt�B4@h�Ð!?�.��(�@��%�ٿ�����I�@ބZt�B4@h�Ð!?�.��(�@��%�ٿ�����I�@ބZt�B4@h�Ð!?�.��(�@��@���ٿ�IW{��@���^4@6Fʬ��!?(��V�U�@M'{��ٿ~۠� �@�,8�4@����!?��QN���@�+�^��ٿ��4�@�6r:�84@�J��5�!?�
c�@�+�^��ٿ��4�@�6r:�84@�J��5�!?�
c�@6���ٿ��h1vK�@��R�34@k��S�!?��(��@6���ٿ��h1vK�@��R�34@k��S�!?��(��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�D�d�ٿ̼vs���@�h��:�3@W�9l-�!?�[�̽��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@�ԙ��ٿ�/!���@[L��H64@(M�!?�M-��@��5ԙٿ�R��s�@)���A4@'�6U,�!?j��<���@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@֟@���ٿ���g�@�r��PT4@����'�!?ê%����@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@���2f�ٿ��YOԝ�@��$�T4@��`�Q�!?I�a>eו@x�iםٿ��5
��@;Q{JV4@	����!?��M��@x�iםٿ��5
��@;Q{JV4@	����!?��M��@x�iםٿ��5
��@;Q{JV4@	����!?��M��@x�iםٿ��5
��@;Q{JV4@	����!?��M��@��ɞٿ�F�[!|�@��W4@���y�!?���q�@X�V��ٿF�O)�G�@"�A�4@�5̞�!?��W��@X�V��ٿF�O)�G�@"�A�4@�5̞�!?��W��@{����ٿ	چ�;�@�7�4@7��!?���W��@{����ٿ	چ�;�@�7�4@7��!?���W��@{����ٿ	چ�;�@�7�4@7��!?���W��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@��m�ٿ��|9��@q�Mf�4@=�S�!?fD&7��@�j�o�ٿ�w��R��@b%���4@r��+�!?�f�:g)�@�j�o�ٿ�w��R��@b%���4@r��+�!?�f�:g)�@oFW5�ٿq��֍�@&�6��3@���!?���7�@oFW5�ٿq��֍�@&�6��3@���!?���7�@R3��ٿRz�=� �@��e���3@N���!?��:O�ʖ@R3��ٿRz�=� �@��e���3@N���!?��:O�ʖ@��C�֚ٿ<MZ����@�S�a��3@����!?��ؗ�/�@��C�֚ٿ<MZ����@�S�a��3@����!?��ؗ�/�@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@1N]d��ٿ�1�P "�@'b*��4@ZV�y�!?�(ˌ ە@�x1�}�ٿ�.ĆZ�@uMm�4@Z4��!?��C��@�x1�}�ٿ�.ĆZ�@uMm�4@Z4��!?��C��@�x1�}�ٿ�.ĆZ�@uMm�4@Z4��!?��C��@�x1�}�ٿ�.ĆZ�@uMm�4@Z4��!?��C��@+�i�/�ٿ���e�9�@��;S4@8Z�#{�!?E���@+�i�/�ٿ���e�9�@��;S4@8Z�#{�!?E���@J*�/�ٿ����L��@��zѝ44@��<�c�!?��]��@J*�/�ٿ����L��@��zѝ44@��<�c�!?��]��@J*�/�ٿ����L��@��zѝ44@��<�c�!?��]��@,j�ۣ�ٿ��wv�}�@��;W�M4@d��f�!?��C���@,j�ۣ�ٿ��wv�}�@��;W�M4@d��f�!?��C���@,j�ۣ�ٿ��wv�}�@��;W�M4@d��f�!?��C���@�e���ٿ�+E����@���:4@"���e�!?}�y㜕@�e���ٿ�+E����@���:4@"���e�!?}�y㜕@�e���ٿ�+E����@���:4@"���e�!?}�y㜕@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@Z��@ �ٿ�.�D��@MJA=��3@���lY�!?Ѽ>_��@�[��:�ٿPl����@�����3@8W��)�!?�+Ck�ʕ@�[��:�ٿPl����@�����3@8W��)�!?�+Ck�ʕ@�[��:�ٿPl����@�����3@8W��)�!?�+Ck�ʕ@Z��$�ٿ<'��>�@
nXf��3@*3�?�!?���j+Ε@Z��$�ٿ<'��>�@
nXf��3@*3�?�!?���j+Ε@Z��$�ٿ<'��>�@
nXf��3@*3�?�!?���j+Ε@���H��ٿ�[���J�@#���4@r���C�!?��ch�@���H��ٿ�[���J�@#���4@r���C�!?��ch�@���=��ٿ�{�D��@�����4@���;��!?�T�Е@W�|��ٿ����!�@$��5l4@j��z�!?Ve!`�@J+q`�ٿc:�.���@�E�-Xk4@\4�{�!?�1��ޕ@�45�ٿC��fw�@</���I4@?�/셐!?�l;���@�45�ٿC��fw�@</���I4@?�/셐!?�l;���@�45�ٿC��fw�@</���I4@?�/셐!?�l;���@�45�ٿC��fw�@</���I4@?�/셐!?�l;���@�45�ٿC��fw�@</���I4@?�/셐!?�l;���@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@~��� �ٿ��> ��@�~�4@�[�AL�!?Z�����@Y3��ٿ��m_�@��b�4@E���!?�I2�V�@i�;ܤ�ٿ����Z-�@��
^54@��+�!?3Hk䆕@i�;ܤ�ٿ����Z-�@��
^54@��+�!?3Hk䆕@i�;ܤ�ٿ����Z-�@��
^54@��+�!?3Hk䆕@|��{|�ٿ&(���V�@��c494@VC�/��!?7��	)�@�f�Y!�ٿ��d��@R�c�d4@�"�L�!?�U�l�@�f�Y!�ٿ��d��@R�c�d4@�"�L�!?�U�l�@+H�^3�ٿHv��@���.4@�.	��!?!|�dΕ@+H�^3�ٿHv��@���.4@�.	��!?!|�dΕ@+H�^3�ٿHv��@���.4@�.	��!?!|�dΕ@+H�^3�ٿHv��@���.4@�.	��!?!|�dΕ@-��ʜٿ4���t�@�Z�Q��3@�[ŀ�!?YXjb@Ε@?`���ٿW�-CP��@v�H4@>o���!?,�ٔ�!�@?`���ٿW�-CP��@v�H4@>o���!?,�ٔ�!�@?`���ٿW�-CP��@v�H4@>o���!?,�ٔ�!�@?`���ٿW�-CP��@v�H4@>o���!?,�ٔ�!�@?`���ٿW�-CP��@v�H4@>o���!?,�ٔ�!�@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@��b<֖ٿ�!�2f�@�K��4@��0�E�!?�+����@�BM�6�ٿ[�t&��@��bat�3@��B�!?'��,��@�BM�6�ٿ[�t&��@��bat�3@��B�!?'��,��@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@RI�ٿ{E�Ļ�@����R�3@j&��<�!?J�şEM�@>�;՘ٿ���U�~�@Ƣӆ��3@���F�!?���&�R�@>�;՘ٿ���U�~�@Ƣӆ��3@���F�!?���&�R�@>�;՘ٿ���U�~�@Ƣӆ��3@���F�!?���&�R�@>�;՘ٿ���U�~�@Ƣӆ��3@���F�!?���&�R�@�:�gԛٿ�S���\�@�0���3@��#&�!?ϔ�$_A�@�:�gԛٿ�S���\�@�0���3@��#&�!?ϔ�$_A�@�:�gԛٿ�S���\�@�0���3@��#&�!?ϔ�$_A�@�:�gԛٿ�S���\�@�0���3@��#&�!?ϔ�$_A�@P?�E+�ٿ�dL����@��Χ��3@Z��n��!?��Fl�@P?�E+�ٿ�dL����@��Χ��3@Z��n��!?��Fl�@P?�E+�ٿ�dL����@��Χ��3@Z��n��!?��Fl�@P?�E+�ٿ�dL����@��Χ��3@Z��n��!?��Fl�@7�V��ٿ~�v����@�.�4@\h�$�!?�.!}��@7�V��ٿ~�v����@�.�4@\h�$�!?�.!}��@7�V��ٿ~�v����@�.�4@\h�$�!?�.!}��@7�V��ٿ~�v����@�.�4@\h�$�!?�.!}��@�7�z�ٿ�G��@�0�)hJ4@�2�.�!?2M��W`�@�;N���ٿ�8ݟЍ�@�2��;U4@���c7�!?�����ޕ@/�ЛٿH�+`���@t�3�0B4@���r��!?ť��@/�ЛٿH�+`���@t�3�0B4@���r��!?ť��@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@~ܖW��ٿ?��u���@���4@�r�9��!?��r%;�@)fϡܙٿ�;�'��@�p�M4@n�mA��!?k��h�@|�{�ٿ�=�Ę`�@�𿾆"4@P��d�!?��5����@|�{�ٿ�=�Ę`�@�𿾆"4@P��d�!?��5����@|�{�ٿ�=�Ę`�@�𿾆"4@P��d�!?��5����@|�{�ٿ�=�Ę`�@�𿾆"4@P��d�!?��5����@|�{�ٿ�=�Ę`�@�𿾆"4@P��d�!?��5����@e�X��ٿ�Q5wM�@ۉ�Q-4@�0�o�!?ŕ$��@e�X��ٿ�Q5wM�@ۉ�Q-4@�0�o�!?ŕ$��@e�X��ٿ�Q5wM�@ۉ�Q-4@�0�o�!?ŕ$��@e�X��ٿ�Q5wM�@ۉ�Q-4@�0�o�!?ŕ$��@��U��ٿ�D
��+�@5M��
24@��g�!?��ch��@��U��ٿ�D
��+�@5M��
24@��g�!?��ch��@��U��ٿ�D
��+�@5M��
24@��g�!?��ch��@��U��ٿ�D
��+�@5M��
24@��g�!?��ch��@��u�ٿ�1��@��H���3@Z�k�;�!?õV�7��@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�����ٿ�k>I���@��
SP4@�
SHɐ!?=sZy5�@�´�ٿ�fͧ��@��o
4@r��N�!?t6�A;,�@�]X�k�ٿV��Iu��@�����3@�RZN�!?��6��@�U4�l�ٿ��AY��@�N2w{4@z*��}�!?1�w���@�U4�l�ٿ��AY��@�N2w{4@z*��}�!?1�w���@�U4�l�ٿ��AY��@�N2w{4@z*��}�!?1�w���@�#w�Ҝٿl
t��@�{g;4@F�O���!?0�?��@�#w�Ҝٿl
t��@�{g;4@F�O���!?0�?��@�#w�Ҝٿl
t��@�{g;4@F�O���!?0�?��@�d'��ٿ`�,���@�$N	�@4@�>��!?_��+���@�d'��ٿ`�,���@�$N	�@4@�>��!?_��+���@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@NL�ޗٿ0n�����@�VS�!4@krȘ�!?G	"�I��@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@����ٿ�;��\��@y�}�wS4@��
���!?2 gDC�@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@n�z�ǜٿq]E����@��1�n:4@��F��!?�kzl�ו@5-Z{�ٿ��o�9�@âf+�3@��<8-�!?ldY@<��@5-Z{�ٿ��o�9�@âf+�3@��<8-�!?ldY@<��@5-Z{�ٿ��o�9�@âf+�3@��<8-�!?ldY@<��@J/��B�ٿL�a���@�ݺ��#4@Qpk1V�!?P�X+�@J/��B�ٿL�a���@�ݺ��#4@Qpk1V�!?P�X+�@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@W��ٜٿ������@Z����3@KV��G�!?耣^^��@��OQR�ٿO.?0��@�X�%�3@�G�D�!?��W��@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@p"��ٿR��Rs�@�	�$� 4@�𩾒�!?� x�e�@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@?��{�ٿ^��<�?�@N��J�3@�� [�!?���ޕ@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@��{粛ٿ��<�t��@#J�)P4@����!?�"6�a&�@�-�z�ٿ��d?�@��V�:	4@y��I��!?�OjNN�@'����ٿ�ء/�E�@�J�a�4@�W��!?�P��쪖@'����ٿ�ء/�E�@�J�a�4@�W��!?�P��쪖@'����ٿ�ء/�E�@�J�a�4@�W��!?�P��쪖@'����ٿ�ء/�E�@�J�a�4@�W��!?�P��쪖@'����ٿ�ء/�E�@�J�a�4@�W��!?�P��쪖@.Z�32�ٿ��d�@~��&4@��`Y�!?yk�����@.Z�32�ٿ��d�@~��&4@��`Y�!?yk�����@�g,��ٿ�bR�#�@#چ-9"4@"\/z_�!?$�~־��@�g,��ٿ�bR�#�@#چ-9"4@"\/z_�!?$�~־��@�g,��ٿ�bR�#�@#چ-9"4@"\/z_�!?$�~־��@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@1��'�ٿ��n���@ϻ�|�Y4@�B.P�!?c��6D�@�`���ٿ�X����@td�6�3@�8���!?��1���@�`���ٿ�X����@td�6�3@�8���!?��1���@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@_s�]�ٿA��YU�@��g\t�3@h��C�!?M�<X��@V�oj�ٿ�n��@-�@8	2�4@�?�=�!?��@૊�@V�oj�ٿ�n��@-�@8	2�4@�?�=�!?��@૊�@V�oj�ٿ�n��@-�@8	2�4@�?�=�!?��@૊�@V�oj�ٿ�n��@-�@8	2�4@�?�=�!?��@૊�@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@������ٿ �i�(�@v�+�~"4@�+&�I�!?ϒ��9ʕ@�����ٿ�Ȳ�.m�@��2΍4@�ZR>�!?��}��@�����ٿ�Ȳ�.m�@��2΍4@�ZR>�!?��}��@��P��ٿM�����@�"�4@Ξ�Fy�!?�)؆��@`CW�ٿOxQ�&>�@$k�:%4@�i�(5�!?=��yOp�@`CW�ٿOxQ�&>�@$k�:%4@�i�(5�!?=��yOp�@�Ͷ���ٿ$��`�@�S�D4@��4���!?�|(�^�@�Ͷ���ٿ$��`�@�S�D4@��4���!?�|(�^�@�Ͷ���ٿ$��`�@�S�D4@��4���!?�|(�^�@�Ͷ���ٿ$��`�@�S�D4@��4���!?�|(�^�@�RdΧٿ�B�Ev'�@�7V�::4@P�t�x�!?��o�k�@�RdΧٿ�B�Ev'�@�7V�::4@P�t�x�!?��o�k�@���Ϟٿ�{����@ϲ�Dw4@����k�!?>�e�Е@���Ϟٿ�{����@ϲ�Dw4@����k�!?>�e�Е@���Ϟٿ�{����@ϲ�Dw4@����k�!?>�e�Е@����ٿ�mI���@R�d�{�4@�$�|��!?Ի�W"��@����ٿ�mI���@R�d�{�4@�$�|��!?Ի�W"��@����ٿ�mI���@R�d�{�4@�$�|��!?Ի�W"��@�,Z�ڦٿ�>�F��@�5GA�b4@�i;J��!?�
��Kݕ@�~a5�ٿ�I�ɬ�@R��E�-4@�O�e�!?�β��ە@�~a5�ٿ�I�ɬ�@R��E�-4@�O�e�!?�β��ە@���Ξٿ�uh#3�@��ؠY84@QlV�!?n�oc0�@���Ξٿ�uh#3�@��ؠY84@QlV�!?n�oc0�@���Ξٿ�uh#3�@��ؠY84@QlV�!?n�oc0�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@7�O�ٿ�)����@+C4�44@$�`��!?�pS�U)�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@��毻�ٿ��7]Ⱥ�@����'4@E�r��!?W'�U�$�@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�7 ���ٿ84A�s�@D�6��*4@�oltl�!?��A���@�¨m�ٿ�5��@�	�G*44@-Q���!?3���0��@�¨m�ٿ�5��@�	�G*44@-Q���!?3���0��@�¨m�ٿ�5��@�	�G*44@-Q���!?3���0��@0t8
#�ٿc��ee�@��u�4@��$�W�!??f)���@0t8
#�ٿc��ee�@��u�4@��$�W�!??f)���@�7��ٿO�h�k�@|"��84@:2�m�!?�Bf���@�9��ٿ�13Yk��@h�I�=4@U�:�!?w�t0р�@�9��ٿ�13Yk��@h�I�=4@U�:�!?w�t0р�@>^wH�ٿf��{^ �@+�u�-)4@4�j�,�!?��C��@a�mu��ٿs��.���@`�Lg4@(P_�!?�&��@a�mu��ٿs��.���@`�Lg4@(P_�!?�&��@a�mu��ٿs��.���@`�Lg4@(P_�!?�&��@-��3��ٿ���_ɡ�@
��*4@�Z�`$�!?.{>�2u�@���F�ٿ\<q1��@���KR�3@yǴ�!?}ߌN��@���F�ٿ\<q1��@���KR�3@yǴ�!?}ߌN��@U?	j��ٿu[����@`&:�K�3@��o+�!?Z�v [Ǖ@U?	j��ٿu[����@`&:�K�3@��o+�!?Z�v [Ǖ@�]xL�ٿ��o��~�@I��-�3@ך��[�!?1��Y��@�]xL�ٿ��o��~�@I��-�3@ך��[�!?1��Y��@�]xL�ٿ��o��~�@I��-�3@ך��[�!?1��Y��@�]xL�ٿ��o��~�@I��-�3@ך��[�!?1��Y��@�]xL�ٿ��o��~�@I��-�3@ך��[�!?1��Y��@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@���z�ٿD�����@-	Z]�3@��@P�!?2 a��k�@�2��W�ٿK�z�p�@}��Ŭ4@�B���!?���6䦕@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@���/�ٿ4x�F�@�~I�3@@6��T�!?z]�iҕ@��|Y̠ٿ(-���@e/��4@	7�Z�!?Y
m��(�@�E����ٿ+ncj��@��x� 4@�"u2�!?5\$��U�@�E����ٿ+ncj��@��x� 4@�"u2�!?5\$��U�@�E����ٿ+ncj��@��x� 4@�"u2�!?5\$��U�@�E����ٿ+ncj��@��x� 4@�"u2�!?5\$��U�@e³�ٿ������@^m_ /�3@����K�!?_�>v�@e³�ٿ������@^m_ /�3@����K�!?_�>v�@e³�ٿ������@^m_ /�3@����K�!?_�>v�@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@���V��ٿ���Ǌ��@�WJ�#\4@�D�!?������@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�NĂ�ٿ�y$��@Ԫ��On4@��/�#�!?T>���@�	�ʞٿڌl̃,�@?�IoH4@E�E"�!?{ͣ3v�@��"&s�ٿt�!�@k�J8J4@����N�!?�V��쮕@��"&s�ٿt�!�@k�J8J4@����N�!?�V��쮕@B.����ٿH3����@��ɩ4@��s�}�!?�F��0��@B.����ٿH3����@��ɩ4@��s�}�!?�F��0��@B.����ٿH3����@��ɩ4@��s�}�!?�F��0��@B.����ٿH3����@��ɩ4@��s�}�!?�F��0��@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@h��}v�ٿs"�jE�@<�)�-)4@�H4��!?�̬wi_�@|A�O��ٿ<0�,�M�@�q�4@��6,��!?����RЕ@|A�O��ٿ<0�,�M�@�q�4@��6,��!?����RЕ@9V\潞ٿ���)���@�����3@�2�89�!?go�@9V\潞ٿ���)���@�����3@�2�89�!?go�@�QNR��ٿu��"�@��4��3@>Y���!?!��	�@�QNR��ٿu��"�@��4��3@>Y���!?!��	�@���ƛ�ٿ<7n<�@���=��3@p�.-�!?~����@���ƛ�ٿ<7n<�@���=��3@p�.-�!?~����@���ƛ�ٿ<7n<�@���=��3@p�.-�!?~����@Kv�O��ٿ!�rx���@��]��3@�Tu�z�!?#gDЭ�@Kv�O��ٿ!�rx���@��]��3@�Tu�z�!?#gDЭ�@Kv�O��ٿ!�rx���@��]��3@�Tu�z�!?#gDЭ�@Kv�O��ٿ!�rx���@��]��3@�Tu�z�!?#gDЭ�@&�p4:�ٿ$�j��@A׳���3@��p�E�!?X�x�N��@�Q�ٿ�Z.9S��@Y	_W�4@�s��5�!?c78E��@�Q�ٿ�Z.9S��@Y	_W�4@�s��5�!?c78E��@#-�t��ٿ�hy��w�@\��%4@&~E\4�!?�.��o[�@#-�t��ٿ�hy��w�@\��%4@&~E\4�!?�.��o[�@�����ٿ��z��@�|]��4@U@N/�!?A�%��˕@���tǝٿ���*��@�39�7^4@1���!?�̜���@���tǝٿ���*��@�39�7^4@1���!?�̜���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@���2��ٿCb��@�@]0Q4@��7�!?�RM+���@�K_��ٿ��Dp�:�@�}L�v4@l�H���!?���T�d�@�K_��ٿ��Dp�:�@�}L�v4@l�H���!?���T�d�@�K_��ٿ��Dp�:�@�}L�v4@l�H���!?���T�d�@�K_��ٿ��Dp�:�@�}L�v4@l�H���!?���T�d�@����؜ٿ��s����@���_P4@���!?W��+�}�@����؜ٿ��s����@���_P4@���!?W��+�}�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@��%勝ٿ�!<��B�@S�h�w4@��r��!?K�!�g�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@6�
Fa�ٿz�*���@y�pP�s4@ML(�!?��~B�@��K��ٿ3&#���@�9D�4@�JzY�!?#~�X&�@ Zr���ٿ\�����@�D���3@7��@r�!?<e�@ Zr���ٿ\�����@�D���3@7��@r�!?<e�@ Zr���ٿ\�����@�D���3@7��@r�!?<e�@ Zr���ٿ\�����@�D���3@7��@r�!?<e�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@QZO�@�ٿ����2C�@w�V4@n P�.�!?����W�@Y  �ٿ?�����@~K`�3@��u#m�!?7��y�ӕ@Y  �ٿ?�����@~K`�3@��u#m�!?7��y�ӕ@Y  �ٿ?�����@~K`�3@��u#m�!?7��y�ӕ@Y  �ٿ?�����@~K`�3@��u#m�!?7��y�ӕ@MkR���ٿ�����@>��E4@ ޑ�.�!?"d@�X��@MkR���ٿ�����@>��E4@ ޑ�.�!?"d@�X��@MkR���ٿ�����@>��E4@ ޑ�.�!?"d@�X��@ø���ٿXr�0]�@(g��a#4@�Պz<�!?��LI�A�@ø���ٿXr�0]�@(g��a#4@�Պz<�!?��LI�A�@ø���ٿXr�0]�@(g��a#4@�Պz<�!?��LI�A�@t;��G�ٿ��f���@®tV
4@���:�!?�� I���@t;��G�ٿ��f���@®tV
4@���:�!?�� I���@t;��G�ٿ��f���@®tV
4@���:�!?�� I���@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@0	7yF�ٿw�� �A�@:}�/S4@��i���!?T����C�@,b\֚ٿG�X4U�@Z��4@cϑK^�!?#c��쩕@,b\֚ٿG�X4U�@Z��4@cϑK^�!?#c��쩕@,b\֚ٿG�X4U�@Z��4@cϑK^�!?#c��쩕@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@\먐��ٿ�o>���@"7N/4@xYl�k�!?SPx@�@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@��F�}�ٿr��Zwl�@��/c4@�a�F��!?�x6���@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@p��ٿ1?���B�@��@�P4@�}�`h�!?8�+�ƕ@ߖ�:3�ٿ����~�@0�E	�C4@�F��!?���d��@ߖ�:3�ٿ����~�@0�E	�C4@�F��!?���d��@ߖ�:3�ٿ����~�@0�E	�C4@�F��!?���d��@ߖ�:3�ٿ����~�@0�E	�C4@�F��!?���d��@��eе�ٿ�{߽��@�?̆B�3@/|!?����1�@��eе�ٿ�{߽��@�?̆B�3@/|!?����1�@��eе�ٿ�{߽��@�?̆B�3@/|!?����1�@Ԑ:�Y�ٿK_��/�@���@%4@Ȓ��0�!?�aGK:��@a�~��ٿҥ}��R�@$��T-4@Bsg�*�!?�/\41��@a�~��ٿҥ}��R�@$��T-4@Bsg�*�!?�/\41��@a�~��ٿҥ}��R�@$��T-4@Bsg�*�!?�/\41��@a�~��ٿҥ}��R�@$��T-4@Bsg�*�!?�/\41��@a�~��ٿҥ}��R�@$��T-4@Bsg�*�!?�/\41��@���d�ٿ|����@�nt�WU4@D�|��!?�e��4�@���d�ٿ|����@�nt�WU4@D�|��!?�e��4�@���d�ٿ|����@�nt�WU4@D�|��!?�e��4�@�lbաٿ�OP�-�@4y�s�n4@���Ų�!?��@�lbաٿ�OP�-�@4y�s�n4@���Ų�!?��@�lbաٿ�OP�-�@4y�s�n4@���Ų�!?��@�lbաٿ�OP�-�@4y�s�n4@���Ų�!?��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@q:�h�ٿ��ʢ=��@ozf��{4@��Ϗ!?t�ٿ��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@E��K�ٿvp�9�@? y��t4@}��a�!?��P�A��@e8�ߠٿ�j�g{�@ y�HAV4@�"`{�!?��K5u�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@%�Xޟٿ��$zs�@i��BK4@:,�V�!?�RV�tC�@b�z�K�ٿ��h��@v��{34@�!�b��!?�krh^�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@�VW�-�ٿ*�~���@V�e�	4@�7U氐!? �h�4�@���h��ٿ��V�v!�@���,c@4@��i#��!?VB�B��@���h��ٿ��V�v!�@���,c@4@��i#��!?VB�B��@���h��ٿ��V�v!�@���,c@4@��i#��!?VB�B��@����X�ٿ��HH��@����#4@���)Y�!?	�Y����@����X�ٿ��HH��@����#4@���)Y�!?	�Y����@����X�ٿ��HH��@����#4@���)Y�!?	�Y����@����X�ٿ��HH��@����#4@���)Y�!?	�Y����@g����ٿ�Zj��a�@^�mG�(4@��1A�!?��G�Q�@g����ٿ�Zj��a�@^�mG�(4@��1A�!?��G�Q�@g����ٿ�Zj��a�@^�mG�(4@��1A�!?��G�Q�@g����ٿ�Zj��a�@^�mG�(4@��1A�!?��G�Q�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@���Y�ٿ��up�8�@��3ox14@��x�L�!?�oᦷt�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@%ǁ�{�ٿ����@c��p*f4@�3�!?F���֦�@��J�ٿy����e�@��ۅU4@�����!?ȲN-��@��J�ٿy����e�@��ۅU4@�����!?ȲN-��@��J�ٿy����e�@��ۅU4@�����!?ȲN-��@��J�ٿy����e�@��ۅU4@�����!?ȲN-��@_W��ٿ4��|��@��T��3@���\:�!?����¿�@_W��ٿ4��|��@��T��3@���\:�!?����¿�@_W��ٿ4��|��@��T��3@���\:�!?����¿�@_W��ٿ4��|��@��T��3@���\:�!?����¿�@_W��ٿ4��|��@��T��3@���\:�!?����¿�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@�ԁ�}�ٿ��q"��@E�TB��3@i�ҷ��!?/u��E�@zhR�ٿ����@�nX�a14@bk�3�!?��4[7�@zhR�ٿ����@�nX�a14@bk�3�!?��4[7�@���D�ٿ$���SY�@��<4@c�U{�!?��1��@���D�ٿ$���SY�@��<4@c�U{�!?��1��@Q�_�ٿGC&��@��f��3@s�V�!?�F;fF�@Q�_�ٿGC&��@��f��3@s�V�!?�F;fF�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@�C0��ٿ��Z����@�?74@X+��H�!?q|�UK�@мN��ٿ��{����@�O�4@�t���!?�G^�QJ�@мN��ٿ��{����@�O�4@�t���!?�G^�QJ�@мN��ٿ��{����@�O�4@�t���!?�G^�QJ�@мN��ٿ��{����@�O�4@�t���!?�G^�QJ�@Lw�rޞٿ�UE���@��mh4@0e=�\�!?؎m�H}�@Lw�rޞٿ�UE���@��mh4@0e=�\�!?؎m�H}�@Lw�rޞٿ�UE���@��mh4@0e=�\�!?؎m�H}�@Lw�rޞٿ�UE���@��mh4@0e=�\�!?؎m�H}�@Lw�rޞٿ�UE���@��mh4@0e=�\�!?؎m�H}�@�5|	�ٿΞ����@4��F%4@�omv�!?[1���#�@�5|	�ٿΞ����@4��F%4@�omv�!?[1���#�@�5|	�ٿΞ����@4��F%4@�omv�!?[1���#�@�5|	�ٿΞ����@4��F%4@�omv�!?[1���#�@�5|	�ٿΞ����@4��F%4@�omv�!?[1���#�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@r����ٿe���c�@�A�	4@��iOH�!?s��b�@˄o_՝ٿ��WB�e�@���^�3@+n��>�!?*l�
�"�@��뀛ٿ�BX���@E���3@RTr=,�!?d�*�%�@��뀛ٿ�BX���@E���3@RTr=,�!?d�*�%�@��뀛ٿ�BX���@E���3@RTr=,�!?d�*�%�@��뀛ٿ�BX���@E���3@RTr=,�!?d�*�%�@��뀛ٿ�BX���@E���3@RTr=,�!?d�*�%�@OD�Yg�ٿ�OK��3�@���`�3@9�y�*�!?��d�!�@OD�Yg�ٿ�OK��3�@���`�3@9�y�*�!?��d�!�@OD�Yg�ٿ�OK��3�@���`�3@9�y�*�!?��d�!�@ݦ�6e�ٿ�%��@�� |e�3@O�)Z]�!?���V��@����~�ٿ���p�@`��k
4@�é�=�!?mkz��@����~�ٿ���p�@`��k
4@�é�=�!?mkz��@����~�ٿ���p�@`��k
4@�é�=�!?mkz��@����~�ٿ���p�@`��k
4@�é�=�!?mkz��@�=X��ٿȮ��� �@���� 4@>�@�G�!?-}�5:�@��=�ٿ����@o��*4@>21�!?��Z��@��=�ٿ����@o��*4@>21�!?��Z��@��=�ٿ����@o��*4@>21�!?��Z��@Ej����ٿH��e��@���S"4@LL�%�!?
O�� �@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@�\�U�ٿ#6Kړ��@q�.���3@n���]�!?C�1$v��@��+e�ٿ@�@�@�P��m"4@"�O�!?�r�XM��@��+e�ٿ@�@�@�P��m"4@"�O�!?�r�XM��@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@���ϟٿ�R���@�i!/��3@���ě�!?��Q�e̕@Y!
c]�ٿ~[���D�@ޝ�y(4@-�{���!?�Y�H��@Y!
c]�ٿ~[���D�@ޝ�y(4@-�{���!?�Y�H��@Y!
c]�ٿ~[���D�@ޝ�y(4@-�{���!?�Y�H��@Y!
c]�ٿ~[���D�@ޝ�y(4@-�{���!?�Y�H��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@��A��ٿJlT2�@��]�3@����v�!?S޺S��@p��ٿ`㚧���@pW���=4@��!?���Cy�@p��ٿ`㚧���@pW���=4@��!?���Cy�@p��ٿ`㚧���@pW���=4@��!?���Cy�@p��ٿ`㚧���@pW���=4@��!?���Cy�@ͺK���ٿ�v>uZ�@A���.4@�ŷ�H�!?�����@ͺK���ٿ�v>uZ�@A���.4@�ŷ�H�!?�����@ͺK���ٿ�v>uZ�@A���.4@�ŷ�H�!?�����@7U$�&�ٿ��d��-�@��X2{�3@�a� 6�!?*���㩖@WZO��ٿ
�rA�@�9۞4@��� �!?���|Rc�@WZO��ٿ
�rA�@�9۞4@��� �!?���|Rc�@WZO��ٿ
�rA�@�9۞4@��� �!?���|Rc�@�T1���ٿ6�Ba�U�@5`\m�3@�f�~��!?�oy��@�t����ٿ[R���U�@8=K�(4@��'R��!?��hV���@�t����ٿ[R���U�@8=K�(4@��'R��!?��hV���@�L�8�ٿ��_P�4�@|㕭�4@E�̐!?<�o,wF�@o�X��ٿ�������@䆼ѹ4@�6m���!?EJr�� �@o�X��ٿ�������@䆼ѹ4@�6m���!?EJr�� �@��
���ٿS���@�JG�=4@����,�!?��ە@��
���ٿS���@�JG�=4@����,�!?��ە@6�J�Q�ٿ|��b��@�1�6u\4@Y�uQJ�!?v�1� ��@6�J�Q�ٿ|��b��@�1�6u\4@Y�uQJ�!?v�1� ��@f��X�ٿtl�]��@] �B�L4@=�tJ�!?���Õ@n��ʝٿS�SR��@;4K�}94@���|�!?z��~��@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@N �j�ٿ�"�`�-�@]0�C�4@�
9�W�!?$!-��y�@:�*g��ٿ^����[�@��!�3@��tXK�!?@}rYi�@�h��ٿٺE(��@ʋylP�3@��.�\�!?���rB-�@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@ �t�H�ٿF7����@0�y�"4@�h�7\�!?��(��@	x�ٿ	�uw��@��Tr	4@)"���!?jSJ�[�@	x�ٿ	�uw��@��Tr	4@)"���!?jSJ�[�@�����ٿ��J�Z\�@��̈́�3@
��q�!?�)�5��@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@C+��ٿ�
ֵI��@!�Ӷ�4@�2�3�!?a�6�7�@\�!��ٿr�)�E��@�nM4@�Vp_t�!?��vW͕@\�!��ٿr�)�E��@�nM4@�Vp_t�!?��vW͕@<g����ٿJ���05�@3g�#�@4@Z?�&�!?��ۢ��@��x��ٿrpVAN�@�d�5\4@Рݏ!?l��J4�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�H�x�ٿw�(V��@.�6+14@�G�$�!?�C+�iE�@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@�5���ٿ\�Y!Y��@���Z� 4@�3�fv�!?�P>���@6�+�ٿ�ϧ����@(�%�		4@�C%Z�!?�~|Hc�@6�+�ٿ�ϧ����@(�%�		4@�C%Z�!?�~|Hc�@p�@�-�ٿ���v��@�{�5�3@��T��!?[�k��@�P�0z�ٿ	��r2�@�ӍX�3@3��|��!?܉;�ɕ@�P�0z�ٿ	��r2�@�ӍX�3@3��|��!?܉;�ɕ@�P�0z�ٿ	��r2�@�ӍX�3@3��|��!?܉;�ɕ@�P�0z�ٿ	��r2�@�ӍX�3@3��|��!?܉;�ɕ@���ͤ�ٿ��{��P�@>߹��24@^�����!?Op;H��@�$��k�ٿ�p�E�@�����4@Zq�4i�!?�

�<�@����ٿ�ʟ�4�@�C��|4@UIk�^�!?	�l�@����ٿ�ʟ�4�@�C��|4@UIk�^�!?	�l�@xh���ٿ����@�c�4�3@���(��!?<�V���@xh���ٿ����@�c�4�3@���(��!?<�V���@xh���ٿ����@�c�4�3@���(��!?<�V���@xh���ٿ����@�c�4�3@���(��!?<�V���@"v>�ٿc�ݫ��@ ��'`(4@� ġ��!?�\ �@�.9�T�ٿӉ	|�@;O�?��3@%w�6��!?�Z]�n;�@�.9�T�ٿӉ	|�@;O�?��3@%w�6��!?�Z]�n;�@�.9�T�ٿӉ	|�@;O�?��3@%w�6��!?�Z]�n;�@)��^�ٿ������@�D#�3@<�\�!?�U��H�@�u���ٿ�`u��@������3@�P�9�!?/f�ڷ=�@�u���ٿ�`u��@������3@�P�9�!?/f�ڷ=�@�u���ٿ�`u��@������3@�P�9�!?/f�ڷ=�@�u���ٿ�`u��@������3@�P�9�!?/f�ڷ=�@�u���ٿ�`u��@������3@�P�9�!?/f�ڷ=�@]I���ٿtv��^��@�uU��3@��h�W�!?��ݘ�@D�4J>�ٿ����3�@��F�3@�9��!?��MZ1'�@D�4J>�ٿ����3�@��F�3@�9��!?��MZ1'�@����ٿ"�� y�@��Η:�3@%�nh�!?�{a���@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@�J��g�ٿg��yf�@�1��E4@�^�I'�!?�eҰ�Ε@'�Ǯ�ٿB���}
�@sH`&Q4@1�]�!?Q�UL
�@'�Ǯ�ٿB���}
�@sH`&Q4@1�]�!?Q�UL
�@B����ٿ�yz����@�dv�U4@s�@|E�!?lAKTݕ@,t!�՟ٿ"(8\�f�@���E/4@��JN�!?�H��ߕ@,t!�՟ٿ"(8\�f�@���E/4@��JN�!?�H��ߕ@���Z�ٿi�:F�@�;�4@����E�!?x��4��@���Z�ٿi�:F�@�;�4@����E�!?x��4��@���Z�ٿi�:F�@�;�4@����E�!?x��4��@�;�Q�ٿ�U�W�@�V�G�O4@6?�pn�!?�J���@���n5�ٿ��%�O��@3��	�4@���cZ�!?���	ݕ@��v&�ٿQ�
(�6�@?��CcP4@k����!?�^ٴ��@��v&�ٿQ�
(�6�@?��CcP4@k����!?�^ٴ��@��v&�ٿQ�
(�6�@?��CcP4@k����!?�^ٴ��@��v&�ٿQ�
(�6�@?��CcP4@k����!?�^ٴ��@��v&�ٿQ�
(�6�@?��CcP4@k����!?�^ٴ��@*׹�Ιٿ�J2���@Ц�]94@�ց��!?/�yLw��@0�ߤ�ٿ�Ӯ���@b -��4@9U/��!?Dd\���@0�ߤ�ٿ�Ӯ���@b -��4@9U/��!?Dd\���@0�ߤ�ٿ�Ӯ���@b -��4@9U/��!?Dd\���@0�ߤ�ٿ�Ӯ���@b -��4@9U/��!?Dd\���@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@/ĺ:Ȗٿ�#K)J�@R3�+4@лQ.��!?�)�}��@s�K�J�ٿ��ZlX��@\�&�L@4@����d�!?�.��9�@s�K�J�ٿ��ZlX��@\�&�L@4@����d�!?�.��9�@s�K�J�ٿ��ZlX��@\�&�L@4@����d�!?�.��9�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@rI�PʚٿKoC���@�帤f4@����!?���� #�@J�ՒL�ٿ]Ԗ�;��@�.c0�4@0���h�!?.�6D1�@Q֡�ٿ��F�@Z"}P-P4@}H&��!?2�PV��@Q֡�ٿ��F�@Z"}P-P4@}H&��!?2�PV��@Q֡�ٿ��F�@Z"}P-P4@}H&��!?2�PV��@t�o`�ٿ��2Z��@�xeB�+4@lll�r�!?ɶ �ŕ@����F�ٿ�j詤<�@3��� 4@�(�xː!?��G9��@����F�ٿ�j詤<�@3��� 4@�(�xː!?��G9��@����F�ٿ�j詤<�@3��� 4@�(�xː!?��G9��@����F�ٿ�j詤<�@3��� 4@�(�xː!?��G9��@�����ٿ�~/HX��@�H,��.4@�b�-s�!?!O�nՕ@�����ٿ�~/HX��@�H,��.4@�b�-s�!?!O�nՕ@&Q�SH�ٿ.�wh��@sQ�{A4@a�g�7�!??���$�@&Q�SH�ٿ.�wh��@sQ�{A4@a�g�7�!??���$�@&Q�SH�ٿ.�wh��@sQ�{A4@a�g�7�!??���$�@&Q�SH�ٿ.�wh��@sQ�{A4@a�g�7�!??���$�@&Q�SH�ٿ.�wh��@sQ�{A4@a�g�7�!??���$�@
)��ٿ"Y�o2M�@��Ց�:4@<��̊�!?�LQR�@
)��ٿ"Y�o2M�@��Ց�:4@<��̊�!?�LQR�@
)��ٿ"Y�o2M�@��Ց�:4@<��̊�!?�LQR�@
)��ٿ"Y�o2M�@��Ց�:4@<��̊�!?�LQR�@
)��ٿ"Y�o2M�@��Ց�:4@<��̊�!?�LQR�@�J�֜ٿ��
L��@l_���(4@�'��w�!?����?�@�J�֜ٿ��
L��@l_���(4@�'��w�!?����?�@�J�֜ٿ��
L��@l_���(4@�'��w�!?����?�@��S\�ٿ#$�(��@'���84@
7��^�!?F�)n!�@��S\�ٿ#$�(��@'���84@
7��^�!?F�)n!�@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@l�u��ٿ�CY^��@�m�m&F4@�saB�!?�]&^��@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@p�ɅR�ٿ6���y��@%�w4
4@T�h��!?�K�{�@0o���ٿ�u#��@[��V�K4@��f�H�!?��f�v�@0o���ٿ�u#��@[��V�K4@��f�H�!?��f�v�@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@%o��ٿ�_��@	3�j4@��m^�!?`�4ז@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@~��|�ٿV��Ĺ[�@�?\��4@ 0�Dr�!?�mbk��@���ܮ�ٿ�/���@��j�3@	�H>H�!?Mh4��@���ܮ�ٿ�/���@��j�3@	�H>H�!?Mh4��@A$j��ٿ0�r����@�D] _�3@� �q�!?�~HL��@A$j��ٿ0�r����@�D] _�3@� �q�!?�~HL��@A$j��ٿ0�r����@�D] _�3@� �q�!?�~HL��@A$j��ٿ0�r����@�D] _�3@� �q�!?�~HL��@A$j��ٿ0�r����@�D] _�3@� �q�!?�~HL��@�O�_��ٿ��/v��@� ��4@պ����!?r�[du��@�O�_��ٿ��/v��@� ��4@պ����!?r�[du��@}�QTßٿ�?��F��@��xa(4@��<-�!?#z"ɩ��@}�QTßٿ�?��F��@��xa(4@��<-�!?#z"ɩ��@}�QTßٿ�?��F��@��xa(4@��<-�!?#z"ɩ��@}�QTßٿ�?��F��@��xa(4@��<-�!?#z"ɩ��@}�QTßٿ�?��F��@��xa(4@��<-�!?#z"ɩ��@�rƲ��ٿ�LMQ��@��b��4@��:���!?K�M����@���מٿ:D)r��@2 ��.4@��TsH�!?f�=�ȕ@���מٿ:D)r��@2 ��.4@��TsH�!?f�=�ȕ@���מٿ:D)r��@2 ��.4@��TsH�!?f�=�ȕ@%��S�ٿ��\���@�=��j94@�J��`�!?���ŵ�@%��S�ٿ��\���@�=��j94@�J��`�!?���ŵ�@%��S�ٿ��\���@�=��j94@�J��`�!?���ŵ�@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@)�1.7�ٿ �)a���@L}�%��3@�ި�]�!?"�}b�ӕ@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@���+�ٿ�p:^|��@���L<4@PQ�#�!?� UR`�@��pA�ٿv`E����@c6!��3@5(}�x�!?z(�p鮕@�b���ٿ�����u�@nO���3@.�M�!?#��X#�@�b���ٿ�����u�@nO���3@.�M�!?#��X#�@�b���ٿ�����u�@nO���3@.�M�!?#��X#�@�b���ٿ�����u�@nO���3@.�M�!?#��X#�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@�	FX��ٿ��x%���@}ʄlg4@ �&�W�!?a���A�@Ǭ{㨜ٿ��/$,��@T�ek��3@6-;�j�!?HswD&��@Ǭ{㨜ٿ��/$,��@T�ek��3@6-;�j�!?HswD&��@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@��"g֟ٿ�d�"��@�"<�l�3@�}�6x�!?K8B"�	�@�rǢA�ٿ(4屘s�@���Z4@5-����!?F����@�rǢA�ٿ(4屘s�@���Z4@5-����!?F����@I�O�ٿ�_�R�@	+m��L4@K�L�J�!?�ڋ��8�@I�O�ٿ�_�R�@	+m��L4@K�L�J�!?�ڋ��8�@I�O�ٿ�_�R�@	+m��L4@K�L�J�!?�ڋ��8�@�ŉ���ٿ �G���@�L#%714@�S9�`�!? N��Е@
,#�=�ٿ-ߟ����@- �204@۔9w8�!?p�ܠ��@�I塤�ٿti��1�@͕�8�4@ŷ��\�!?]�(`k�@�I塤�ٿti��1�@͕�8�4@ŷ��\�!?]�(`k�@�I塤�ٿti��1�@͕�8�4@ŷ��\�!?]�(`k�@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@Hr�e�ٿp��A�V�@n�%�4@[�o_M�!?N�4�L��@�n$�ٿ߻m�rU�@�i��5I4@`{L��!?b-_�\W�@��b���ٿ�(�J�@��|Y�#4@�P���!?qO�<���@��b���ٿ�(�J�@��|Y�#4@�P���!?qO�<���@��b���ٿ�(�J�@��|Y�#4@�P���!?qO�<���@��b���ٿ�(�J�@��|Y�#4@�P���!?qO�<���@�zdd�ٿ���X!�@�dj�U34@���`�!?9�]�B�@�zdd�ٿ���X!�@�dj�U34@���`�!?9�]�B�@��o�ٿ��@D:��@��:Z-�3@�)���!?����&ߕ@��o�ٿ��@D:��@��:Z-�3@�)���!?����&ߕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@7ϰ�ٿ��v� ��@$�U��4@:R�,�!?���gƕ@퇴Şٿ�\=zyT�@��P�4@�Q�h�!?<=�E˕@�7���ٿ���#r�@�% V�'4@�״_�!?����A�@�����ٿ���Bc��@V�X�@4@�2�A�!?��?�̕@����ٿT�3RFX�@�=�\G4@�ۃ�!?f��=\#�@����ٿT�3RFX�@�=�\G4@�ۃ�!?f��=\#�@����ٿT�3RFX�@�=�\G4@�ۃ�!?f��=\#�@_��~�ٿ&�M���@�T��DD4@W~�'��!?�u\�WΖ@_��~�ٿ&�M���@�T��DD4@W~�'��!?�u\�WΖ@8۱���ٿKUZ]�w�@xj �ut4@A{^�!?e��%?�@8۱���ٿKUZ]�w�@xj �ut4@A{^�!?e��%?�@8۱���ٿKUZ]�w�@xj �ut4@A{^�!?e��%?�@8۱���ٿKUZ]�w�@xj �ut4@A{^�!?e��%?�@�V_E�ٿ'��D�@���E�a4@�l._��!? [m�ĕ@�V_E�ٿ'��D�@���E�a4@�l._��!? [m�ĕ@�V_E�ٿ'��D�@���E�a4@�l._��!? [m�ĕ@ib`�2�ٿ�h)~�@;���p�3@��Q�!?�~�N~�@ib`�2�ٿ�h)~�@;���p�3@��Q�!?�~�N~�@ib`�2�ٿ�h)~�@;���p�3@��Q�!?�~�N~�@ib`�2�ٿ�h)~�@;���p�3@��Q�!?�~�N~�@ib`�2�ٿ�h)~�@;���p�3@��Q�!?�~�N~�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@���`�ٿO�Ȁ�\�@��J�3@dS��k�!?m�0�|�@�ò �ٿ����"�@!�l4a�3@��<|6�!?i 3���@�ò �ٿ����"�@!�l4a�3@��<|6�!?i 3���@�ò �ٿ����"�@!�l4a�3@��<|6�!?i 3���@����>�ٿ�g�����@�H��3@�%��!?��� ��@6M�s��ٿ����}��@�K)�6�3@�@�y�!?)�6)�b�@6M�s��ٿ����}��@�K)�6�3@�@�y�!?)�6)�b�@��D�ٿJT��@��-���3@�ƕ��!?_��&�@~ǿ5�ٿ菳j�5�@OG��4@x-M��!?�T���C�@~ǿ5�ٿ菳j�5�@OG��4@x-M��!?�T���C�@m�O�ٿ��+���@/����4@�$(Ð!?�R6.M	�@m�O�ٿ��+���@/����4@�$(Ð!?�R6.M	�@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@��bI��ٿ��|/�@�o�]
4@~ �X�!?ag Y6͕@e�I��ٿ�o���@~
��4@�S(��!?�Z;ৰ�@e�I��ٿ�o���@~
��4@�S(��!?�Z;ৰ�@���, �ٿ�-g�@��9�4@mD��R�!?������@��he�ٿ̝����@{U04@�0��!?T@;���@��he�ٿ̝����@{U04@�0��!?T@;���@��he�ٿ̝����@{U04@�0��!?T@;���@�Ⱥ_�ٿwh��P�@��]e�$4@�}�l�!?�e"�
+�@�Ⱥ_�ٿwh��P�@��]e�$4@�}�l�!?�e"�
+�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@ˍ�[�ٿa$+�h��@�q	��3@�Q�!?4��_]�@`�R�'�ٿ,2�bMl�@A\
'4@����!?��Qqx�@`�R�'�ٿ,2�bMl�@A\
'4@����!?��Qqx�@`�R�'�ٿ,2�bMl�@A\
'4@����!?��Qqx�@ ��+g�ٿ��"���@yQ��3�3@ S��!?#��;���@�#7g��ٿ��(>un�@�g���4@��EǏ!?V���@�#7g��ٿ��(>un�@�g���4@��EǏ!?V���@�#7g��ٿ��(>un�@�g���4@��EǏ!?V���@�!�c�ٿ"�KӾ{�@�Tow�3@ç��ď!?��C\��@�!�c�ٿ"�KӾ{�@�Tow�3@ç��ď!?��C\��@�X*Иٿ1g͉D�@�i���3@�7�3#�!?Ũ�X�X�@�X*Иٿ1g͉D�@�i���3@�7�3#�!?Ũ�X�X�@�X*Иٿ1g͉D�@�i���3@�7�3#�!?Ũ�X�X�@�X*Иٿ1g͉D�@�i���3@�7�3#�!?Ũ�X�X�@�X*Иٿ1g͉D�@�i���3@�7�3#�!?Ũ�X�X�@�l]Q�ٿ�\�?D��@����p4@�n���!?oK�r�@�l]Q�ٿ�\�?D��@����p4@�n���!?oK�r�@�l]Q�ٿ�\�?D��@����p4@�n���!?oK�r�@�l]Q�ٿ�\�?D��@����p4@�n���!?oK�r�@��N֛ٿ�2%#+�@	
"\�@4@9N�@��!?2���P��@��N֛ٿ�2%#+�@	
"\�@4@9N�@��!?2���P��@�=�Y�ٿ�'?���@����F4@p �>k�!?Z�ӝ���@�=�Y�ٿ�'?���@����F4@p �>k�!?Z�ӝ���@�� �ٿ����kY�@��b4@yK�*��!?<=$�L�@�� �ٿ����kY�@��b4@yK�*��!?<=$�L�@A}L#"�ٿS��8��@NqBW4@9��*ʐ!?��V%�L�@A}L#"�ٿS��8��@NqBW4@9��*ʐ!?��V%�L�@A}L#"�ٿS��8��@NqBW4@9��*ʐ!?��V%�L�@>��ٿ�N@fZ��@����?4@�2nz�!?yE&�{7�@sY$�?�ٿ�o��"�@^+��O4@-�:b�!?�'2���@sY$�?�ٿ�o��"�@^+��O4@-�:b�!?�'2���@sY$�?�ٿ�o��"�@^+��O4@-�:b�!?�'2���@;by�[�ٿ�����@n��QE4@�|=L�!?�ڤs��@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�;��ٿ߯2��_�@n��"�L4@@6�_�!?g��M�@�
�p�ٿ��HKn�@v�8��'4@Ҋ'W��!?g=��p�@�"`��ٿ* ���@)����3@�@Q=�!?�G����@}�"ħٿ�$����@��-8O4@�c�i�!?��xIM�@}�"ħٿ�$����@��-8O4@�c�i�!?��xIM�@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@|B�3�ٿ����@6,�-X4@_��j�!?��_e�ƕ@���̧�ٿ��	�g)�@g�-�]4@Jv��o�!?q�#g�@���̧�ٿ��	�g)�@g�-�]4@Jv��o�!?q�#g�@���̧�ٿ��	�g)�@g�-�]4@Jv��o�!?q�#g�@���̧�ٿ��	�g)�@g�-�]4@Jv��o�!?q�#g�@���̧�ٿ��	�g)�@g�-�]4@Jv��o�!?q�#g�@|[K���ٿ^������@sv�,�=4@���XH�!?tX�VL�@|[K���ٿ^������@sv�,�=4@���XH�!?tX�VL�@|[K���ٿ^������@sv�,�=4@���XH�!?tX�VL�@|[K���ٿ^������@sv�,�=4@���XH�!?tX�VL�@|[K���ٿ^������@sv�,�=4@���XH�!?tX�VL�@����ٿ
�`g"�@�J�(T4@|f���!?P��	"�@����ٿ
�`g"�@�J�(T4@|f���!?P��	"�@����ٿ
�`g"�@�J�(T4@|f���!?P��	"�@����ٿ
�`g"�@�J�(T4@|f���!?P��	"�@���kѢٿ������@�.
�'4@��,;N�!?�r9��@���kѢٿ������@�.
�'4@��,;N�!?�r9��@���kѢٿ������@�.
�'4@��,;N�!?�r9��@���kѢٿ������@�.
�'4@��,;N�!?�r9��@���kѢٿ������@�.
�'4@��,;N�!?�r9��@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@9�F�ٿk�S�6�@�ŕQ^4@����{�!?��<g���@�����ٿB@�<��@�k�%4@r�'뒐!?Ur�t���@\�QmB�ٿ��M����@����?4@3�����!?v"��O��@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@���S�ٿ�W�o��@��aa4@�6�z��!?�D�,-X�@x6Ӥ�ٿ�ѿ.�@&���=4@����H�!?9��^���@x6Ӥ�ٿ�ѿ.�@&���=4@����H�!?9��^���@x6Ӥ�ٿ�ѿ.�@&���=4@����H�!?9��^���@x6Ӥ�ٿ�ѿ.�@&���=4@����H�!?9��^���@���z�ٿxz��w��@O�2�A4@��(ΐ!?���Ŋ�@?�A�b�ٿs�҉B�@���JN44@Q�_IE�!??�Yr�$�@?�A�b�ٿs�҉B�@���JN44@Q�_IE�!??�Yr�$�@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@֩rv�ٿ
5�5�@>~u`��3@xab�5�!?�i }⫕@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@��J�ٿ�t�~��@<~~�0�3@�D�.�!?���ܕ@�ZE֞ٿ�rZ�W�@�V��0�3@W�5�!?�:6,�y�@�ZE֞ٿ�rZ�W�@�V��0�3@W�5�!?�:6,�y�@�2C^��ٿ�l8����@l�C 4@n�?ή�!?�/Q�B�@�2C^��ٿ�l8����@l�C 4@n�?ή�!?�/Q�B�@�2C^��ٿ�l8����@l�C 4@n�?ή�!?�/Q�B�@�2C^��ٿ�l8����@l�C 4@n�?ή�!?�/Q�B�@`'�3E�ٿ��#>+��@���Y�,4@Sĝ�6�!?@�_	�@`'�3E�ٿ��#>+��@���Y�,4@Sĝ�6�!?@�_	�@�|�<�ٿ<�>0��@̃�ԁL4@���4N�!?JJG�'��@�|�<�ٿ<�>0��@̃�ԁL4@���4N�!?JJG�'��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@k�f^�ٿ�^��y��@��J4@��x�!?Ly�@��@9��sC�ٿ$̌���@�'�U4@�1J}�!?MIE�c�@��̉�ٿJ�k(��@����<4@�S`B?�!?bYl�'��@��̉�ٿJ�k(��@����<4@�S`B?�!?bYl�'��@��̉�ٿJ�k(��@����<4@�S`B?�!?bYl�'��@��̉�ٿJ�k(��@����<4@�S`B?�!?bYl�'��@�ME�ٿ���(���@�8�Z�#4@��<�~�!?��ٕ@�ME�ٿ���(���@�8�Z�#4@��<�~�!?��ٕ@�ME�ٿ���(���@�8�Z�#4@��<�~�!?��ٕ@�ME�ٿ���(���@�8�Z�#4@��<�~�!?��ٕ@�ME�ٿ���(���@�8�Z�#4@��<�~�!?��ٕ@���Țٿ���3�@g��R�	4@���Ð!?���@�� 
�ٿ��`[���@�A�o4@��۬^�!?��Mb���@VċE��ٿ&ȶ[!*�@N]���!4@>،;�!?�����@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�g��Ԟٿ;)u��@�S7�-	4@��ڔ�!?�N�I ��@�nm���ٿ��yN6/�@N`L�K4@=l<��!?�M]�Qѕ@�nm���ٿ��yN6/�@N`L�K4@=l<��!?�M]�Qѕ@�nm���ٿ��yN6/�@N`L�K4@=l<��!?�M]�Qѕ@�*��X�ٿH������@�e'��'4@�ȣq�!?��9�O�@�*��X�ٿH������@�e'��'4@�ȣq�!?��9�O�@�*��X�ٿH������@�e'��'4@�ȣq�!?��9�O�@�*��X�ٿH������@�e'��'4@�ȣq�!?��9�O�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@��4�ٿ7������@�t�c*4@i>iݱ�!?#���f9�@w���ٿ�5����@��-�344@��;��!?��}g�	�@w���ٿ�5����@��-�344@��;��!?��}g�	�@w���ٿ�5����@��-�344@��;��!?��}g�	�@����Ξٿ�Z<���@�vv�A4@�enV�!?�c��p��@����Ξٿ�Z<���@�vv�A4@�enV�!?�c��p��@����Ξٿ�Z<���@�vv�A4@�enV�!?�c��p��@����Ξٿ�Z<���@�vv�A4@�enV�!?�c��p��@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@�ZC��ٿ,��%�C�@S�s�
4@��5C�!?��ݼy�@D�����ٿ����~�@�1��W�3@���X5�!?x%ˋ~.�@D�����ٿ����~�@�1��W�3@���X5�!?x%ˋ~.�@D�����ٿ����~�@�1��W�3@���X5�!?x%ˋ~.�@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@����ʠٿPO�����@����3@gN㊐!?� �� �@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@���v�ٿ�բ�K�@ ��{�.4@�`F�H�!?}�ͩ)�@�1��ٿ�Nh4�=�@�RL��b4@@cr�B�!?p���I�@~�f+�ٿ8�1��@s�ƍQ4@x(5��!?ظ_tT�@~�f+�ٿ8�1��@s�ƍQ4@x(5��!?ظ_tT�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@fU^���ٿlKՒn��@޶o�jB4@��/<u�!?���<V�@H%��J�ٿئ�]��@�Mh��64@u�@�d�!?Bε-E�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@7��ٿ/�����@�� ��3@:v�T�!?:�m�9�@;�R�-�ٿtP�g���@ R�3@��s��!?�z:?EЕ@;�R�-�ٿtP�g���@ R�3@��s��!?�z:?EЕ@;�R�-�ٿtP�g���@ R�3@��s��!?�z:?EЕ@;�R�-�ٿtP�g���@ R�3@��s��!?�z:?EЕ@;�R�-�ٿtP�g���@ R�3@��s��!?�z:?EЕ@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@@�"��ٿ���Q�@�9����3@DH̩;�!?\��(�@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@Ƴ���ٿm#�4��@��v�4@��=S�!?� X��@�'U���ٿn:P��@�[�(14@ź�hw�!?�zX��
�@�'U���ٿn:P��@�[�(14@ź�hw�!?�zX��
�@�hnw�ٿ��
*<�@zK��4@C�q�!?�k��&�@%��oZ�ٿ�����@3B���3@`���T�!?�Fl<D�@%��oZ�ٿ�����@3B���3@`���T�!?�Fl<D�@%��oZ�ٿ�����@3B���3@`���T�!?�Fl<D�@m��>�ٿ�(,ϟ$�@���3@�@�}Z�!?P��`n�@m��>�ٿ�(,ϟ$�@���3@�@�}Z�!?P��`n�@E��ID�ٿ��"���@�Vߌ��3@:�!Ў�!?���]���@E��ID�ٿ��"���@�Vߌ��3@:�!Ў�!?���]���@E��ID�ٿ��"���@�Vߌ��3@:�!Ў�!?���]���@E��ID�ٿ��"���@�Vߌ��3@:�!Ў�!?���]���@�~ٿ�M�2���@؛~Z��3@��	�!?\w*�@�~ٿ�M�2���@؛~Z��3@��	�!?\w*�@�~ٿ�M�2���@؛~Z��3@��	�!?\w*�@�~ٿ�M�2���@؛~Z��3@��	�!?\w*�@ �)*�ٿJ���p�@)g���3@ O)�!?�@��!�@ �)*�ٿJ���p�@)g���3@ O)�!?�@��!�@0#b�m�ٿ칇 ��@��3�
4@^Qό�!?qF=��ܕ@� �@�ٿz�ѓ���@jb{��3@�rU�!?ժ��U�@��#�ٿ�D�7�@�l�Q�3@��Rd�!?�e-���@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@����Ęٿ�Rt�e��@�0��4@�A�;�!?�mZ"i��@�?%R�ٿ�<�w#��@�غM>4@��&$A�!?���8ݕ@�?%R�ٿ�<�w#��@�غM>4@��&$A�!?���8ݕ@����ٿ��r�@A�'.4@X_L߇�!?����Bݕ@�+�k�ٿ�1�v��@���
4@��ߋ�!?5�&��@�+�k�ٿ�1�v��@���
4@��ߋ�!?5�&��@�ŏΉ�ٿWe�!���@��)r4@�C>�!?�	�F#h�@�ŏΉ�ٿWe�!���@��)r4@�C>�!?�	�F#h�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@�����ٿV�L��C�@ҳQ4@0�:���!?�l���X�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@>�|��ٿQ�v�x/�@K ��N)4@��z��!?L4Ѐb�@�y��^�ٿ@__B��@�Z��3@����d�!?/��e�ܕ@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@Ҙ �ٿ���Û��@�#a7��3@����:�!?�({�:�@�$�Z��ٿҌ?L�@�v�G�3@a��64�!?����?�@��⁺�ٿ}҈�"��@ܣ��3@@�B�!?��{�u�@��⁺�ٿ}҈�"��@ܣ��3@@�B�!?��{�u�@�4��ٿC��m}i�@�A�,E�3@��!H�!?�A[�(��@�4��ٿC��m}i�@�A�,E�3@��!H�!?�A[�(��@�4��ٿC��m}i�@�A�,E�3@��!H�!?�A[�(��@�a<)P�ٿ�A�-9�@:�a<��3@��bJ�!?�̿�c��@�a<)P�ٿ�A�-9�@:�a<��3@��bJ�!?�̿�c��@u rs�ٿ������@6��8N�3@�/�6F�!?�0�Z6z�@u rs�ٿ������@6��8N�3@�/�6F�!?�0�Z6z�@u rs�ٿ������@6��8N�3@�/�6F�!?�0�Z6z�@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@>*�ٿ�������@0[թ�3@�SKY2�!?x�V����@?.#�ٿ���	�@F�#x��3@�0STi�!?6�1��ӕ@?.#�ٿ���	�@F�#x��3@�0STi�!?6�1��ӕ@?.#�ٿ���	�@F�#x��3@�0STi�!?6�1��ӕ@?.#�ٿ���	�@F�#x��3@�0STi�!?6�1��ӕ@?.#�ٿ���	�@F�#x��3@�0STi�!?6�1��ӕ@�-��ٿ�=ѩR�@rPP��3@�+	;�!?��m��x�@8��!ԙٿ��./>��@�����3@4���!?O8�;/��@8��!ԙٿ��./>��@�����3@4���!?O8�;/��@8��!ԙٿ��./>��@�����3@4���!?O8�;/��@8��!ԙٿ��./>��@�����3@4���!?O8�;/��@8��!ԙٿ��./>��@�����3@4���!?O8�;/��@-EX�ٿŷ���@�(�/�>4@��W�!?%��ᦕ@-EX�ٿŷ���@�(�/�>4@��W�!?%��ᦕ@�:6��ٿ��c�'��@.�*�C4@�&��O�!?��| �?�@�:6��ٿ��c�'��@.�*�C4@�&��O�!?��| �?�@�:6��ٿ��c�'��@.�*�C4@�&��O�!?��| �?�@TC��G�ٿy��0�^�@!Y/��S4@XY�lY�!?+H����@TC��G�ٿy��0�^�@!Y/��S4@XY�lY�!?+H����@TC��G�ٿy��0�^�@!Y/��S4@XY�lY�!?+H����@���
�ٿ1�QoM�@M�`�P4@������!?3�c��@���
�ٿ1�QoM�@M�`�P4@������!?3�c��@���
�ٿ1�QoM�@M�`�P4@������!?3�c��@���
�ٿ1�QoM�@M�`�P4@������!?3�c��@+UT�ٿ	 ۏ��@!��0%4@谵���!?i��Ӊ��@]����ٿ�pm�&�@6��.�"4@xP���!?��$����@]����ٿ�pm�&�@6��.�"4@xP���!?��$����@]����ٿ�pm�&�@6��.�"4@xP���!?��$����@,_c��ٿճY��1�@U5 غ3@P�AH��!?�����ϕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@Mk���ٿN S��@�� A�3@Ȼ����!?zv��ȕ@J�ǅ�ٿ��[��@#է���3@s�v_�!?����6�@J�ǅ�ٿ��[��@#է���3@s�v_�!?����6�@J�ǅ�ٿ��[��@#է���3@s�v_�!?����6�@�[̎��ٿ3�:wy�@����3@į=�k�!?�Zz�/]�@�ʹ��ٿ���Z�@�cq�h�3@w��I.�!?�Q�N�6�@��M�=�ٿ8�k ���@��%|/�3@6]�Q�!?����@��M�=�ٿ8�k ���@��%|/�3@6]�Q�!?����@��M�=�ٿ8�k ���@��%|/�3@6]�Q�!?����@��M�=�ٿ8�k ���@��%|/�3@6]�Q�!?����@��M�=�ٿ8�k ���@��%|/�3@6]�Q�!?����@��dm�ٿβ�"j��@�OEY .4@��bv�!?�3}����@��dm�ٿβ�"j��@�OEY .4@��bv�!?�3}����@��dm�ٿβ�"j��@�OEY .4@��bv�!?�3}����@�}_��ٿg�k][#�@�D�@';4@����!?�E\��C�@c���ٿ�9�yQ�@�C�i��3@�צ���!?W3� 
֕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@'��ʜ�ٿ�R?�׸�@ެw ��3@������!?�c��᱕@m:�A��ٿ�Hq0��@��E4@� 	0��!?��{t�@�7���ٿ��W8A��@᫹�k4@�X§�!?gm�K�@�7���ٿ��W8A��@᫹�k4@�X§�!?gm�K�@�7���ٿ��W8A��@᫹�k4@�X§�!?gm�K�@�7���ٿ��W8A��@᫹�k4@�X§�!?gm�K�@u9�*��ٿ������@�H���3@�YqL��!?�� �Օ@u9�*��ٿ������@�H���3@�YqL��!?�� �Օ@u9�*��ٿ������@�H���3@�YqL��!?�� �Օ@����Q�ٿ/!XN�@����3@��ٱ�!?fG�.7,�@����Q�ٿ/!XN�@����3@��ٱ�!?fG�.7,�@����Q�ٿ/!XN�@����3@��ٱ�!?fG�.7,�@�:Q�ٿ)}��@�O�U;4@?e8 ��!?Ρp�9��@�.�i��ٿ���M�a�@y�%�=P4@�1o��!??�ť��@�.�i��ٿ���M�a�@y�%�=P4@�1o��!??�ť��@�ikȿ�ٿl�h��@ٕ��=4@!]-\��!?e����^�@�ikȿ�ٿl�h��@ٕ��=4@!]-\��!?e����^�@�ikȿ�ٿl�h��@ٕ��=4@!]-\��!?e����^�@�W�ٱ�ٿ�e4di��@�%� 4@4�m���!?��s�5�@�W�ٱ�ٿ�e4di��@�%� 4@4�m���!?��s�5�@oJ��˗ٿ"��Ȕ��@"�*��A4@b}l��!?ΧOh�.�@oJ��˗ٿ"��Ȕ��@"�*��A4@b}l��!?ΧOh�.�@
�P�4�ٿ����L�@<)�C�14@��ɒ�!?�O���6�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@��"�ٿ��EJ0�@��L��'4@E5�i�!?�y�d�,�@@�A�ԝٿ~IO�f�@ش9�Y�3@@�{r�!?!��J�ҕ@@�A�ԝٿ~IO�f�@ش9�Y�3@@�{r�!?!��J�ҕ@@�A�ԝٿ~IO�f�@ش9�Y�3@@�{r�!?!��J�ҕ@@�A�ԝٿ~IO�f�@ش9�Y�3@@�{r�!?!��J�ҕ@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@���Șٿ$�s�@���=Q&4@Y��`�!?v=K<� �@��kq�ٿ�.�����@��\F4@�0��F�!?�w�����@��kq�ٿ�.�����@��\F4@�0��F�!?�w�����@��kq�ٿ�.�����@��\F4@�0��F�!?�w�����@��kq�ٿ�.�����@��\F4@�0��F�!?�w�����@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@UW�v̗ٿE�蹦�@>f�(��3@f�)l��!?̥T�g�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@HM�șٿ�Y.B���@��K�4@{tx�!? T��w�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�R��X�ٿ\g!0�)�@Pf�v�74@��F>r�!?<�8s"�@�V!^�ٿ�=�9R�@@*P�4@݈�졐!?�ɝ�`�@�V!^�ٿ�=�9R�@@*P�4@݈�졐!?�ɝ�`�@���ס�ٿs��5^�@!ԒM��3@l�=Z��!?�����@���ס�ٿs��5^�@!ԒM��3@l�=Z��!?�����@���ס�ٿs��5^�@!ԒM��3@l�=Z��!?�����@���ס�ٿs��5^�@!ԒM��3@l�=Z��!?�����@���ס�ٿs��5^�@!ԒM��3@l�=Z��!?�����@_<Fc}�ٿ)��G�K�@g ���3@�c��!?6#d�l��@_<Fc}�ٿ)��G�K�@g ���3@�c��!?6#d�l��@_<Fc}�ٿ)��G�K�@g ���3@�c��!?6#d�l��@�!6���ٿ�*މ���@+s��5�3@,,�*��!?�����@�!6���ٿ�*މ���@+s��5�3@,,�*��!?�����@�!6���ٿ�*މ���@+s��5�3@,,�*��!?�����@�!6���ٿ�*މ���@+s��5�3@,,�*��!?�����@6��b#�ٿ��Ycb �@0�EW�3@	��͐!?��
9�3�@6��b#�ٿ��Ycb �@0�EW�3@	��͐!?��
9�3�@6��b#�ٿ��Ycb �@0�EW�3@	��͐!?��
9�3�@�E�iОٿDJ(jv��@�40R+�3@���Գ�!?��e��@Nf���ٿ�ĈRx�@��884@!f���!?LM�O���@Nf���ٿ�ĈRx�@��884@!f���!?LM�O���@Nf���ٿ�ĈRx�@��884@!f���!?LM�O���@Nf���ٿ�ĈRx�@��884@!f���!?LM�O���@�^r���ٿ>#���@���1,�3@ᙵF��!?	t�K�@�^r���ٿ>#���@���1,�3@ᙵF��!?	t�K�@�^r���ٿ>#���@���1,�3@ᙵF��!?	t�K�@�^r���ٿ>#���@���1,�3@ᙵF��!?	t�K�@~va��ٿح�����@�H��4@�� �!?)���#��@�)��%�ٿ�����@@���4@.�M��!?��R��l�@�)��%�ٿ�����@@���4@.�M��!?��R��l�@�H��1�ٿ=۔�,n�@���Y4@eF�G�!?����@�H��1�ٿ=۔�,n�@���Y4@eF�G�!?����@�H��1�ٿ=۔�,n�@���Y4@eF�G�!?����@W���ٿژ��6�@��h@Ds4@� ��}�!?QAk���@W���ٿژ��6�@��h@Ds4@� ��}�!?QAk���@!���D�ٿx%I���@k�u�="4@`�ID�!?�P+@�Օ@��u-��ٿA�@<�@��(O�#4@�<�#�!?
��ir�@ֵAǚٿc��f{��@N���3@2 ��!?G����@/k���ٿ6h�8,�@9v��3@V��j�!?�)�r�@/k���ٿ6h�8,�@9v��3@V��j�!?�)�r�@/k���ٿ6h�8,�@9v��3@V��j�!?�)�r�@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@n�G�ٿ�cO��*�@���7�3@|	,�z�!?��a����@h�u�ٿ������@��F�4@VVD�A�!?Ԥ+o���@h�u�ٿ������@��F�4@VVD�A�!?Ԥ+o���@h�u�ٿ������@��F�4@VVD�A�!?Ԥ+o���@�����ٿ�W�G���@�6���=4@��%��!?jҟҊ\�@�����ٿ�W�G���@�6���=4@��%��!?jҟҊ\�@�����ٿ�W�G���@�6���=4@��%��!?jҟҊ\�@�����ٿ�W�G���@�6���=4@��%��!?jҟҊ\�@H
����ٿ��}���@/�U��+4@��L�X�!?���'�`�@&ܕ�>�ٿ�Aՙ0�@�u tA4@�-ùV�!?jzrON�@&ܕ�>�ٿ�Aՙ0�@�u tA4@�-ùV�!?jzrON�@&ܕ�>�ٿ�Aՙ0�@�u tA4@�-ùV�!?jzrON�@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��bp�ٿ\8 8!��@/B�ńY4@��.
��!?v7P���@��#��ٿ�i��@�d�[4@��랐!??Z�V}�@��#��ٿ�i��@�d�[4@��랐!??Z�V}�@��#��ٿ�i��@�d�[4@��랐!??Z�V}�@��#��ٿ�i��@�d�[4@��랐!??Z�V}�@�E>��ٿ\ڷ3���@u �*=4@���u�!?ʴ�OZ�@�E>��ٿ\ڷ3���@u �*=4@���u�!?ʴ�OZ�@�E>��ٿ\ڷ3���@u �*=4@���u�!?ʴ�OZ�@�E>��ٿ\ڷ3���@u �*=4@���u�!?ʴ�OZ�@�,���ٿ?��� ��@�+>4�3@��b#�!?ɋ��@)f�ȿ�ٿνY�o�@��[`"�3@���&��!?W?�s�@Ƨ��x�ٿ��#�@��Pm�=4@�'Ĝ��!?')/	�{�@Ƨ��x�ٿ��#�@��Pm�=4@�'Ĝ��!?')/	�{�@l)�=k�ٿQ��oZg�@��u�04@r#�Ґ!?��}Z<��@l)�=k�ٿQ��oZg�@��u�04@r#�Ґ!?��}Z<��@���ef�ٿ̏��Ǡ�@
�Ǣ4@fi�o�!?�o"6��@���ef�ٿ̏��Ǡ�@
�Ǣ4@fi�o�!?�o"6��@V�="�ٿ������@z�h��(4@�4�4U�!?O��]s̕@V�="�ٿ������@z�h��(4@�4�4U�!?O��]s̕@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@�˜�ٿ=��	6�@ླྀE4@�4@�6�!?�����@M\?'��ٿq�wRb��@5���3@V��u�!?���^(��@M\?'��ٿq�wRb��@5���3@V��u�!?���^(��@S��&�ٿ�u���@_O̼&4@�U����!?)?�It�@S��&�ٿ�u���@_O̼&4@�U����!?)?�It�@S��&�ٿ�u���@_O̼&4@�U����!?)?�It�@S��&�ٿ�u���@_O̼&4@�U����!?)?�It�@�K�4�ٿ~����@T�g�3@){����!?��dޕ@�K�4�ٿ~����@T�g�3@){����!?��dޕ@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@lo�(�ٿ�|SW�@�����3@��]�!?=�����@����f�ٿz�r����@te�(P4@蜍n�!?-"u${�@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@,Ns���ٿ`�����@��ir�'4@+��%��!?�dH��@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@=A�h��ٿ�����@�T�{:4@�����!?�%�ߔƕ@�RޫO�ٿ�N2���@�$��84@"E�׫�!?�f֑i�@�RޫO�ٿ�N2���@�$��84@"E�׫�!?�f֑i�@�RޫO�ٿ�N2���@�$��84@"E�׫�!?�f֑i�@J� %Y�ٿ�_j��@���_C4@7��8b�!?�2cÕ@J� %Y�ٿ�_j��@���_C4@7��8b�!?�2cÕ@J� %Y�ٿ�_j��@���_C4@7��8b�!?�2cÕ@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@bw���ٿ�w`����@����)04@�_��!?0�_�w��@xh�֬�ٿ~�2��@�@'�9k34@�����!?��g�ʕ@3h��T�ٿ�R:S1�@�v�#`%4@��K�f�!?���le��@3h��T�ٿ�R:S1�@�v�#`%4@��K�f�!?���le��@3h��T�ٿ�R:S1�@�v�#`%4@��K�f�!?���le��@3h��T�ٿ�R:S1�@�v�#`%4@��K�f�!?���le��@3h��T�ٿ�R:S1�@�v�#`%4@��K�f�!?���le��@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@C�D蛘ٿ�����@�{{�3@������!?6��<���@'�H���ٿ��后��@�+ņ�Z4@������!?�u?a��@'�H���ٿ��后��@�+ņ�Z4@������!?�u?a��@�g`���ٿ`�<t��@A �-"4@�
X�d�!?|%��[�@�g`���ٿ`�<t��@A �-"4@�
X�d�!?|%��[�@�g`���ٿ`�<t��@A �-"4@�
X�d�!?|%��[�@�Lܙ��ٿ:�d�_0�@�W�5�3@2���2�!?���̕@�Lܙ��ٿ:�d�_0�@�W�5�3@2���2�!?���̕@�e��ٿ(yQB!�@J�V���3@��ߗ@�!?6F�����@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�٪f�ٿJ�|�	��@kw��]-4@���k�!?ybI-��@�PZɟٿf�Ӹԑ�@���sD4@���o�!?*�@ݕ@�PZɟٿf�Ӹԑ�@���sD4@���o�!?*�@ݕ@�PZɟٿf�Ӹԑ�@���sD4@���o�!?*�@ݕ@�PZɟٿf�Ӹԑ�@���sD4@���o�!?*�@ݕ@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@~���ٿ_����@�WI-4@�ɘ(_�!?&�-R8�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@���`�ٿ�0��?�@����w�3@"ނ�=�!?`�#	`9�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@E:�7�ٿ�������@M�����3@3��qc�!?��o�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@�K��ٿB�� ��@#W�+4@GT!4�!?\yy�H�@ZL��ٿ�Â���@L�u�b	4@F��!?�4YH�+�@��3K�ٿ�7T���@�YYdO$4@�����!?nf���@�/�Cٜٿ�����@��k�>4@P*���!?n�ֿ�ĕ@��p��ٿ�Yő���@�z��0:4@�y)��!?B��/o!�@��p��ٿ�Yő���@�z��0:4@�y)��!?B��/o!�@��p��ٿ�Yő���@�z��0:4@�y)��!?B��/o!�@��p��ٿ�Yő���@�z��0:4@�y)��!?B��/o!�@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@; ���ٿ>�ʁtT�@�߮Y�_4@<���G�!?fp�Nڕ@�&֟ٿ��Ic���@;_�|54@�k�HQ�!?|DK2.�@�&֟ٿ��Ic���@;_�|54@�k�HQ�!?|DK2.�@�&֟ٿ��Ic���@;_�|54@�k�HQ�!?|DK2.�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@��*'G�ٿ����n�@����f4@6�Ac�!?TrX�2:�@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@�^-��ٿ�-÷�b�@�>�LrQ4@���g�!?=U�k���@L�:�ٿ�~r��@�͚�_4@;v��`�!?s�P��@L�:�ٿ�~r��@�͚�_4@;v��`�!?s�P��@L�:�ٿ�~r��@�͚�_4@;v��`�!?s�P��@���ٿ4�%��@.j(�E4@D0M�x�!?�J�XJ��@���ٿ4�%��@.j(�E4@D0M�x�!?�J�XJ��@ÀJ�1�ٿQ�ס=��@�@��/4@C�6N�!?w/���@ÀJ�1�ٿQ�ס=��@�@��/4@C�6N�!?w/���@C3��s�ٿ>���>��@wLΐ�4@og�!?d��:��@C3��s�ٿ>���>��@wLΐ�4@og�!?d��:��@I��� �ٿ��@2���@��j�/34@(��#�!?�0���@I��� �ٿ��@2���@��j�/34@(��#�!?�0���@I��� �ٿ��@2���@��j�/34@(��#�!?�0���@73p4іٿ���A�*�@���1(G4@�v=Q�!?~[hyq�@73p4іٿ���A�*�@���1(G4@�v=Q�!?~[hyq�@p�(��ٿPj#,�@M��B�n4@��(�!?�]��3�@p�(��ٿPj#,�@M��B�n4@��(�!?�]��3�@gt��ٿ���A�{�@�]�9Z4@��{i�!?�1%vDЕ@gt��ٿ���A�{�@�]�9Z4@��{i�!?�1%vDЕ@gt��ٿ���A�{�@�]�9Z4@��{i�!?�1%vDЕ@gt��ٿ���A�{�@�]�9Z4@��{i�!?�1%vDЕ@gt��ٿ���A�{�@�]�9Z4@��{i�!?�1%vDЕ@��1�ٿE����@o/��4@)M;~*�!?��?�e�@��1�ٿE����@o/��4@)M;~*�!?��?�e�@z�^d��ٿh"6��@䘥,4@Y�У-�!?_�8��@z�^d��ٿh"6��@䘥,4@Y�У-�!?_�8��@�|���ٿ�.�����@�m�[�3@X�q�4�!?M;��̗�@�|���ٿ�.�����@�m�[�3@X�q�4�!?M;��̗�@�|���ٿ�.�����@�m�[�3@X�q�4�!?M;��̗�@ʭ� �ٿo��1J�@X �g4@�U��@�!?.e�2�v�@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@��ٿ��"�@OYu��>4@ ���h�!?j���@�����ٿW��b�@xD��4@2Yjv�!?Q��̕@4�x���ٿ�Y��V;�@�����D4@�H1X�!?�8m�2��@4�x���ٿ�Y��V;�@�����D4@�H1X�!?�8m�2��@4�x���ٿ�Y��V;�@�����D4@�H1X�!?�8m�2��@4�x���ٿ�Y��V;�@�����D4@�H1X�!?�8m�2��@4�x���ٿ�Y��V;�@�����D4@�H1X�!?�8m�2��@�����ٿr�B��@Z�Wy�O4@
i6^�!?��A*���@�����ٿr�B��@Z�Wy�O4@
i6^�!?��A*���@�����ٿr�B��@Z�Wy�O4@
i6^�!?��A*���@�����ٿr�B��@Z�Wy�O4@
i6^�!?��A*���@�����ٿr�B��@Z�Wy�O4@
i6^�!?��A*���@$>�)��ٿ������@	���04@�6�m�!?N�'��@$>�)��ٿ������@	���04@�6�m�!?N�'��@�%�v��ٿ�إ/J��@��cz�4@��F��!?+�.���@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@>�Bɝٿgn����@�#��4@���P��!?�f�0;�@���I�ٿ�ZIc t�@��8�
�3@���*~�!?��P�l��@���I�ٿ�ZIc t�@��8�
�3@���*~�!?��P�l��@���I�ٿ�ZIc t�@��8�
�3@���*~�!?��P�l��@�����ٿ���,�@G'�'��3@u)"�Z�!?�qN�N��@����Ԣٿ�����"�@o��vm�3@�B�I�!?>���ؕ@����Ԣٿ�����"�@o��vm�3@�B�I�!?>���ؕ@����Ԣٿ�����"�@o��vm�3@�B�I�!?>���ؕ@����Ԣٿ�����"�@o��vm�3@�B�I�!?>���ؕ@����Ԣٿ�����"�@o��vm�3@�B�I�!?>���ؕ@wb[:ˡٿB7R����@����o4@�5�)g�!?��n���@wb[:ˡٿB7R����@����o4@�5�)g�!?��n���@wb[:ˡٿB7R����@����o4@�5�)g�!?��n���@wb[:ˡٿB7R����@����o4@�5�)g�!?��n���@\&�^�ٿ���G��@8���$4@x �L&�!?8zc(� �@\&�^�ٿ���G��@8���$4@x �L&�!?8zc(� �@��UiW�ٿsP	y��@6��~4@!CZ~1�!?���=��@��UiW�ٿsP	y��@6��~4@!CZ~1�!?���=��@��UiW�ٿsP	y��@6��~4@!CZ~1�!?���=��@��UiW�ٿsP	y��@6��~4@!CZ~1�!?���=��@b$��ǡٿI����@����(4@�f�yh�!?G�(93Օ@[|��o�ٿ���f���@]_��W4@
�N��!?h�E}Ǖ@v�ѝ�ٿ��y���@{�u��(4@c	r�[�!?�w�U^�@v�ѝ�ٿ��y���@{�u��(4@c	r�[�!?�w�U^�@v�ѝ�ٿ��y���@{�u��(4@c	r�[�!?�w�U^�@v�ѝ�ٿ��y���@{�u��(4@c	r�[�!?�w�U^�@v�ѝ�ٿ��y���@{�u��(4@c	r�[�!?�w�U^�@�?��ɟٿ���K>�@����64@h[ڨ*�!?�d�)�ȕ@�?��ɟٿ���K>�@����64@h[ڨ*�!?�d�)�ȕ@�?��ɟٿ���K>�@����64@h[ڨ*�!?�d�)�ȕ@�?��ɟٿ���K>�@����64@h[ڨ*�!?�d�)�ȕ@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@�v�ٿ�ʣ9�@N�I�-
4@f�{<�!?XE�DP��@?��֚ٿ�K��@>���z�3@VbP�+�!?���zM	�@|ތ+�ٿ��I�l�@��+��
4@�bp6W�!?�����@���ҕ�ٿ�,�j��@R����3@�Ft�!?J�u63�@���ҕ�ٿ�,�j��@R����3@�Ft�!?J�u63�@���ҕ�ٿ�,�j��@R����3@�Ft�!?J�u63�@,m��;�ٿ7���,��@�ԼV�4@��[��!?�і�@,m��;�ٿ7���,��@�ԼV�4@��[��!?�і�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@_����ٿİT�eS�@���P�"4@KE���!?�Y�(�@a�f�ٿ��	c�8�@��zJ��3@�͌g�!?* t'�2�@[��Q��ٿ&M���A�@�R���3@	_ CV�!?p���AE�@[��Q��ٿ&M���A�@�R���3@	_ CV�!?p���AE�@?��l�ٿ[��8(��@�]y��3@����!?zk�O-f�@?��l�ٿ[��8(��@�]y��3@����!?zk�O-f�@���:äٿtİN)�@ȹ<Q�3@H]5L�!?&<2QQ��@���:äٿtİN)�@ȹ<Q�3@H]5L�!?&<2QQ��@u��aK�ٿ�KB�T�@�Xr,��3@:%�.�!?`LC�.�@u��aK�ٿ�KB�T�@�Xr,��3@:%�.�!?`LC�.�@�$eO��ٿ9��J�@��CP�N4@6�
T�!?��3��G�@�$eO��ٿ9��J�@��CP�N4@6�
T�!?��3��G�@�$eO��ٿ9��J�@��CP�N4@6�
T�!?��3��G�@�$eO��ٿ9��J�@��CP�N4@6�
T�!?��3��G�@�$eO��ٿ9��J�@��CP�N4@6�
T�!?��3��G�@#�μ��ٿ[{�����@�B�M4@�o{��!?�s���@#�μ��ٿ[{�����@�B�M4@�o{��!?�s���@�$��ٿiI����@��6��.4@YSU�!?�،��@���ٿ*����@� �v�94@�����!?����@���ٿ*����@� �v�94@�����!?����@���ٿ*����@� �v�94@�����!?����@Rn�ܞٿu[̇��@E�U~��3@�tk��!?U����@Rn�ܞٿu[̇��@E�U~��3@�tk��!?U����@Rn�ܞٿu[̇��@E�U~��3@�tk��!?U����@Rn�ܞٿu[̇��@E�U~��3@�tk��!?U����@Rn�ܞٿu[̇��@E�U~��3@�tk��!?U����@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@Xs��ٿcM��8��@�%N�3@�H��!?�j�&|�@�@5�T�ٿ���be�@��s�D�3@}h���!?�X����@�@5�T�ٿ���be�@��s�D�3@}h���!?�X����@�@5�T�ٿ���be�@��s�D�3@}h���!?�X����@�@5�T�ٿ���be�@��s�D�3@}h���!?�X����@�@5�T�ٿ���be�@��s�D�3@}h���!?�X����@��,�ٿ�1�ԡ�@饱T84@A��ܐ!?Ō��<�@��E��ٿ��� H��@b�N�4@e�`*�!?S�"I��@#��+�ٿ�;��P�@�
h��3@��ŗ/�!?�VP�
�@#��+�ٿ�;��P�@�
h��3@��ŗ/�!?�VP�
�@#��+�ٿ�;��P�@�
h��3@��ŗ/�!?�VP�
�@#��+�ٿ�;��P�@�
h��3@��ŗ/�!?�VP�
�@�$���ٿ@�����@�a�k��3@�`	��!?o�	 #<�@�$���ٿ@�����@�a�k��3@�`	��!?o�	 #<�@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@J0zv�ٿ�8�Zj�@�h�Ny�3@��\�ҏ!?8N��@�hq�g�ٿ�ޱ|.�@K_��:,4@�Q��!?�%��@�hq�g�ٿ�ޱ|.�@K_��:,4@�Q��!?�%��@�hq�g�ٿ�ޱ|.�@K_��:,4@�Q��!?�%��@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@���t�ٿ��'���@�0!ʉ4@-k�d�!?�i �o<�@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�s)k0�ٿ�-�C4�@���b4@U�xb�!?�j(��@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@�]�R�ٿ2�"�-�@0����4@���d��!?;�\`y�@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@ LD��ٿ�]R��	�@<��(R4@��"�{�!?�Ĩ�b��@={&Ԝٿ܍��rV�@gKЁ��3@atq�1�!?Pl�l���@={&Ԝٿ܍��rV�@gKЁ��3@atq�1�!?Pl�l���@={&Ԝٿ܍��rV�@gKЁ��3@atq�1�!?Pl�l���@q���ٿ����X��@ڱ��G�3@[k��!?�O<̉+�@���ٿ9j��x��@�:᫄3@��HH�!?�� eՕ@���ٿ9j��x��@�:᫄3@��HH�!?�� eՕ@*�͒?�ٿ������@�:
�3@i�=�e�!?sQ�4֮�@*�͒?�ٿ������@�:
�3@i�=�e�!?sQ�4֮�@�bM+�ٿ@������@���E�3@?x��q�!?"���[��@�bM+�ٿ@������@���E�3@?x��q�!?"���[��@�����ٿ�[�X��@���4@�RУy�!?��q���@�����ٿ�[�X��@���4@�RУy�!?��q���@�����ٿ�[�X��@���4@�RУy�!?��q���@�����ٿ�[�X��@���4@�RУy�!?��q���@�����ٿ�[�X��@���4@�RУy�!?��q���@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@�_�?_�ٿ��o-�@�.�d�3@�JA�!?fKh�A��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@4c�f�ٿ]����h�@E���4@��U;>�!?O�Mek��@���᎛ٿu�L��s�@��_�4@����d�!?��I�ڕ@���
��ٿ�/Ӆ7;�@�GHEZ4@��/v�!?,w��~)�@���
��ٿ�/Ӆ7;�@�GHEZ4@��/v�!?,w��~)�@���
��ٿ�/Ӆ7;�@�GHEZ4@��/v�!?,w��~)�@�GM�ٿ����@͸���!4@���c��!?����)�@�GM�ٿ����@͸���!4@���c��!?����)�@�GM�ٿ����@͸���!4@���c��!?����)�@�GM�ٿ����@͸���!4@���c��!?����)�@�GM�ٿ����@͸���!4@���c��!?����)�@�GM�ٿ����@͸���!4@���c��!?����)�@�^���ٿ����bd�@��N�@4@Ra��א!?�qU���@�^���ٿ����bd�@��N�@4@Ra��א!?�qU���@�^���ٿ����bd�@��N�@4@Ra��א!?�qU���@�^���ٿ����bd�@��N�@4@Ra��א!?�qU���@��ܖ��ٿ��sOHw�@����3@�]�i��!?�`���@��ܖ��ٿ��sOHw�@����3@�]�i��!?�`���@��ܖ��ٿ��sOHw�@����3@�]�i��!?�`���@��ܖ��ٿ��sOHw�@����3@�]�i��!?�`���@��ܖ��ٿ��sOHw�@����3@�]�i��!?�`���@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@ j �N�ٿ�_x�O��@)GF���3@�`XN�!?���|�2�@��1c��ٿ����W �@��V�3@  @փ�!?����; �@��1c��ٿ����W �@��V�3@  @փ�!?����; �@��1c��ٿ����W �@��V�3@  @փ�!?����; �@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@��_~ʚٿ�)8!c�@]�B�4@���-��!?�97r��@
���C�ٿ�����@fu��C04@�;p�!?������@
���C�ٿ�����@fu��C04@�;p�!?������@
���C�ٿ�����@fu��C04@�;p�!?������@
���C�ٿ�����@fu��C04@�;p�!?������@
���C�ٿ�����@fu��C04@�;p�!?������@
���C�ٿ�����@fu��C04@�;p�!?������@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�/ڹx�ٿ��D����@�;m�4@J�MdJ�!?0��'7ߕ@�eFS�ٿ��^
�@��{�h4@)���'�!?D���@�eFS�ٿ��^
�@��{�h4@)���'�!?D���@�eFS�ٿ��^
�@��{�h4@)���'�!?D���@�eFS�ٿ��^
�@��{�h4@)���'�!?D���@�e��ٿ�((�O��@��4@-�,y�!?�LY�ɕ@�e��ٿ�((�O��@��4@-�,y�!?�LY�ɕ@�e��ٿ�((�O��@��4@-�,y�!?�LY�ɕ@�e��ٿ�((�O��@��4@-�,y�!?�LY�ɕ@բ�]�ٿ���@���	4@�d�l�!?������@բ�]�ٿ���@���	4@�d�l�!?������@^\��ٿ�G�+�o�@�V��4@��VK�!?]^┬��@��&&��ٿ�jWw���@&x�SP4@�m)�l�!?��akꖕ@�� Č�ٿ8����@��%�D4@�Dc�p�!?�(�|��@�� Č�ٿ8����@��%�D4@�Dc�p�!?�(�|��@�� Č�ٿ8����@��%�D4@�Dc�p�!?�(�|��@V�]�ٿ�����@e��*�>4@�[��!?�o���ݕ@V�]�ٿ�����@e��*�>4@�[��!?�o���ݕ@�Z�6�ٿs��(���@f%���R4@�m,0�!?g)�u�$�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@��u�s�ٿ�dd��@��@�N4@�!��{�!?���jh�@�����ٿ�����@��ꆏ4@d��J��!?
/��8��@sD◚ٿ4m����@.��R4@�Lo�!?�̓�T]�@sD◚ٿ4m����@.��R4@�Lo�!?�̓�T]�@Hg˚ٿ�J��Z`�@b4tm�D4@�qGя�!?bO2�VI�@�H���ٿ����k�@�{�kz4@��@h�!?Ħz���@�H���ٿ����k�@�{�kz4@��@h�!?Ħz���@=��ٿ�6�����@�i��4@&�?C �!?�sډ�ە@=��ٿ�6�����@�i��4@&�?C �!?�sډ�ە@=��ٿ�6�����@�i��4@&�?C �!?�sډ�ە@�DAN��ٿ1bJ?�$�@k�p�Q4@�[x���!?��ځq�@P�R���ٿ����-��@�Uߥb4@�|A3�!?r8I����@8����ٿ��b��@����o4@��7�!?�ߍ�2��@8����ٿ��b��@����o4@��7�!?�ߍ�2��@8����ٿ��b��@����o4@��7�!?�ߍ�2��@8����ٿ��b��@����o4@��7�!?�ߍ�2��@8����ٿ��b��@����o4@��7�!?�ߍ�2��@7�!�Ԙٿ9u����@��zr4@
�Xa�!?�K�-��@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@���`�ٿ����j�@Vx�M=4@��x?�!?o:����@�����ٿ� ���@!dQw�4@b�!?��i�ӕ@&rWQ�ٿ6��K�h�@�EQ��3@����P�!?��W"R�@&rWQ�ٿ6��K�h�@�EQ��3@����P�!?��W"R�@ �>AO�ٿY�5��@����s�3@:�-�w�!?�@�#�@ �>AO�ٿY�5��@����s�3@:�-�w�!?�@�#�@ �>AO�ٿY�5��@����s�3@:�-�w�!?�@�#�@ �>AO�ٿY�5��@����s�3@:�-�w�!?�@�#�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@cp�D��ٿ(�/f��@������3@�LCc�!?���_�@Mi�d�ٿ��� �@B��,��3@Z���f�!?nۆ�kO�@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@�T��ٿ�VT�F0�@���	4@��_�!?�<~֕@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@���5v�ٿW���@``3.4@ip�t!�!?]����@�7o+)�ٿ#������@���MD4@���Z�!?f����Е@�7o+)�ٿ#������@���MD4@���Z�!?f����Е@�7o+)�ٿ#������@���MD4@���Z�!?f����Е@b��Wܜٿ%��_b��@��}��4@���i�!?��B썕@b��Wܜٿ%��_b��@��}��4@���i�!?��B썕@b��Wܜٿ%��_b��@��}��4@���i�!?��B썕@b��Wܜٿ%��_b��@��}��4@���i�!?��B썕@b��Wܜٿ%��_b��@��}��4@���i�!?��B썕@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@��:͊�ٿ�G`a�`�@�o�4@���O �!?�FOV@ƕ@g��y0�ٿJ��n��@E��.4@�
�!?�1��@g��y0�ٿJ��n��@E��.4@�
�!?�1��@g��y0�ٿJ��n��@E��.4@�
�!?�1��@g��y0�ٿJ��n��@E��.4@�
�!?�1��@��^�_�ٿ��cJXm�@7Fΐ�4@A.�rF�!?5뚱<�@��^�_�ٿ��cJXm�@7Fΐ�4@A.�rF�!?5뚱<�@��^�_�ٿ��cJXm�@7Fΐ�4@A.�rF�!?5뚱<�@�M�ɹ�ٿ:��1#�@�����3@�J��!?&����@�i�}9�ٿ��Ԧ�@�(��U�3@�C��r�!?�3q�ɕ@�i�}9�ٿ��Ԧ�@�(��U�3@�C��r�!?�3q�ɕ@�i�}9�ٿ��Ԧ�@�(��U�3@�C��r�!?�3q�ɕ@�i�}9�ٿ��Ԧ�@�(��U�3@�C��r�!?�3q�ɕ@U�	%,�ٿ����u�@	��#4@�=��y�!?a�j:�@U�	%,�ٿ����u�@	��#4@�=��y�!?a�j:�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@�-ޞw�ٿH�'����@]��@4@�/�?�!?�C�
�@eE�Z�ٿ�9Ā&�@��.��+4@�[��]�!?���b8"�@eE�Z�ٿ�9Ā&�@��.��+4@�[��]�!?���b8"�@eE�Z�ٿ�9Ā&�@��.��+4@�[��]�!?���b8"�@�F����ٿB~(�B^�@�xH4@x,U�!?�1��F�@�F����ٿB~(�B^�@�xH4@x,U�!?�1��F�@�F����ٿB~(�B^�@�xH4@x,U�!?�1��F�@rx*D�ٿ�w��@�v���4@�u;6�!?D�[��$�@KoT͚ٿy�h�qp�@��<�k4@gC�!?!�|���@KoT͚ٿy�h�qp�@��<�k4@gC�!?!�|���@KoT͚ٿy�h�qp�@��<�k4@gC�!?!�|���@KoT͚ٿy�h�qp�@��<�k4@gC�!?!�|���@KoT͚ٿy�h�qp�@��<�k4@gC�!?!�|���@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@��빖ٿbE��o��@���m<4@�T 5�!?F�3H�M�@���"ߗٿZш����@�R���3@YQ�!?���)6�@��AL�ٿ롣�T��@z��5:4@%Wаt�!?ɭ��LN�@��AL�ٿ롣�T��@z��5:4@%Wаt�!?ɭ��LN�@��AL�ٿ롣�T��@z��5:4@%Wаt�!?ɭ��LN�@��AL�ٿ롣�T��@z��5:4@%Wаt�!?ɭ��LN�@��,�ٿ�P�Y,�@0R-�U_4@A�F�!?�\��Q�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@ta���ٿ�����@T2&�>4@�%�+Y�!?v3hG�(�@"�Lɥ�ٿ$�n����@f-�|�#4@l���m�!?�3���@"�Lɥ�ٿ$�n����@f-�|�#4@l���m�!?�3���@/�=w5�ٿ��/��`�@�:9Z��3@�6�Od�!?�I���@/�=w5�ٿ��/��`�@�:9Z��3@�6�Od�!?�I���@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@��-�N�ٿ�鲴��@�����3@Y�YT�!?���}�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@���:N�ٿ�@����@Ն��624@��J�m�!?)#ϳ�@�Ͱ��ٿ�ф�T�@5+�4@�����!?E���ȕ@�Ͱ��ٿ�ф�T�@5+�4@�����!?E���ȕ@�Ͱ��ٿ�ф�T�@5+�4@�����!?E���ȕ@^G��ɗٿ�ᜳJ�@�Gd,4@�4Ň�!?�ˆ2�@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@V�(˝ٿ�J
�@�ΜU�3@�x��!?�g�� ��@R��ߘٿ�3V�<�@	M5J24@����h�!?m'@k�_�@R��ߘٿ�3V�<�@	M5J24@����h�!?m'@k�_�@R��ߘٿ�3V�<�@	M5J24@����h�!?m'@k�_�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��WY�ٿc��?���@�o6�:4@Fcd�!?#-y�a�@��C��ٿ(�:���@�k��n-4@Vދɐ!?;���@��C��ٿ(�:���@�k��n-4@Vދɐ!?;���@�����ٿ�$�n�@�|�qD4@k��z��!?-�^���@�����ٿ�$�n�@�|�qD4@k��z��!?-�^���@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@M�Sn��ٿ��QEk�@�m�wD4@���i��!? %�]�:�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@�n(�ٿ'�����@�n74@Ό�'��!?��8ik�@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@{-�m�ٿ��.��@��[��-4@�t^HT�!?`��}��@�:��	�ٿZl�j���@�^p\�4@�s"^\�!?~&p�)M�@��L�ٿ3����	�@C����4@�+�a��!?M�kW��@>B�h�ٿ���WF�@���H4@�U>�)�!?��ӥ���@��4N��ٿ+��`y{�@�A4@	��>�!?�Ձ�1�@��4N��ٿ+��`y{�@�A4@	��>�!?�Ձ�1�@��4N��ٿ+��`y{�@�A4@	��>�!?�Ձ�1�@�祼��ٿ��rѭ�@Q�*}��3@v�4O8�!? ��B��@���ןٿ��0�5��@�ԡ84@[�	�w�!?�%/��@���ןٿ��0�5��@�ԡ84@[�	�w�!?�%/��@���ןٿ��0�5��@�ԡ84@[�	�w�!?�%/��@nR��ٿ#�U#I��@���I��3@t�ƣe�!?GnM
���@nR��ٿ#�U#I��@���I��3@t�ƣe�!?GnM
���@nR��ٿ#�U#I��@���I��3@t�ƣe�!?GnM
���@nR��ٿ#�U#I��@���I��3@t�ƣe�!?GnM
���@7�G�O�ٿ?��:<{�@�b�&�3@��c~E�!?jx����@7�G�O�ٿ?��:<{�@�b�&�3@��c~E�!?jx����@�n�r�ٿ��X�Lj�@\+k74@��G?�!?������@�n�r�ٿ��X�Lj�@\+k74@��G?�!?������@XS�l�ٿ��zyE��@S�q�IC4@w{�9��!?VD��@XS�l�ٿ��zyE��@S�q�IC4@w{�9��!?VD��@XS�l�ٿ��zyE��@S�q�IC4@w{�9��!?VD��@XS�l�ٿ��zyE��@S�q�IC4@w{�9��!?VD��@���/�ٿxM�:��@��6��"4@�qɜ�!?��L���@���/�ٿxM�:��@��6��"4@�qɜ�!?��L���@!)�8G�ٿ"��sr�@�u�� 4@t	z�i�!?T﹁YY�@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@Ӧ^�ٿ\B�?A��@�y6.4@���zv�!?��G�d��@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@�Y}w��ٿ}�h&^��@p �>4@;m�(k�!?����@'��{��ٿ
ט� �@� ��Sj4@��N�*�!?aqI��@�nj?�ٿ��$r���@h�In,4@�%�&�!?�	��#~�@�nj?�ٿ��$r���@h�In,4@�%�&�!?�	��#~�@�nj?�ٿ��$r���@h�In,4@�%�&�!?�	��#~�@t��B�ٿ����@�[d�+�3@)�B��!?۪��ޕ@t��B�ٿ����@�[d�+�3@)�B��!?۪��ޕ@t��B�ٿ����@�[d�+�3@)�B��!?۪��ޕ@t��B�ٿ����@�[d�+�3@)�B��!?۪��ޕ@��޸�ٿ��'�f �@|�!��4@:�"��!?�B�)�@��޸�ٿ��'�f �@|�!��4@:�"��!?�B�)�@��~�ԣٿ�#_����@^��ɹ�3@[Pۙ��!?|� 
x�@��~�ԣٿ�#_����@^��ɹ�3@[Pۙ��!?|� 
x�@��~�ԣٿ�#_����@^��ɹ�3@[Pۙ��!?|� 
x�@��bO�ٿ�cJ�+��@6�u�3@�d;S��!?��|��@��bO�ٿ�cJ�+��@6�u�3@�d;S��!?��|��@��bO�ٿ�cJ�+��@6�u�3@�d;S��!?��|��@���>�ٿH��Ƈ��@���3@���!?�=��@&MpW�ٿHo��@_��
4@*��K?�!?�{��@&MpW�ٿHo��@_��
4@*��K?�!?�{��@&MpW�ٿHo��@_��
4@*��K?�!?�{��@&MpW�ٿHo��@_��
4@*��K?�!?�{��@Q�;f.�ٿ�ҋ,\�@�ّl�3@�q�l�!?��#��@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@��n��ٿ�����@L��ȕ�3@�@��L�!?������@�\� ��ٿ����0��@rm7�A4@`km�!?l=�*ի�@�\� ��ٿ����0��@rm7�A4@`km�!?l=�*ի�@����T�ٿ�zfԧ��@tr�G�4@�lO��!? V�R�@����T�ٿ�zfԧ��@tr�G�4@�lO��!? V�R�@[@	��ٿ��h��o�@,~�Iu4@�!��ݐ!?*�"��I�@[@	��ٿ��h��o�@,~�Iu4@�!��ݐ!?*�"��I�@[@	��ٿ��h��o�@,~�Iu4@�!��ݐ!?*�"��I�@[@	��ٿ��h��o�@,~�Iu4@�!��ݐ!?*�"��I�@�RTYΜٿ�����@^?���!4@��X࿐!?�mw=�@Ҷ76�ٿ�+�"�@��ifd4@�~ՓŐ!?��mk�@Ҷ76�ٿ�+�"�@��ifd4@�~ՓŐ!?��mk�@U{� �ٿ�	D���@%_�4@�!�֢�!?۞�x�@U{� �ٿ�	D���@%_�4@�!�֢�!?۞�x�@��C&�ٿLS��-x�@����&4@z�<���!?�sJ��@�6��ٿ�1p�L�@o�\y�L4@G��5�!?��@�g:�t�ٿ!����Y�@Q�?�)4@�,2.�!?+[˗~��@�g:�t�ٿ!����Y�@Q�?�)4@�,2.�!?+[˗~��@�g:�t�ٿ!����Y�@Q�?�)4@�,2.�!?+[˗~��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�6E��ٿ�I����@,����f4@E��u�!?�RiL��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�"�q�ٿ@�?:��@����^4@���c�!?V��%E��@�m���ٿ��}�3�@4�0�{4@��^���!?cc~��@�m���ٿ��}�3�@4�0�{4@��^���!?cc~��@�m���ٿ��}�3�@4�0�{4@��^���!?cc~��@�m���ٿ��}�3�@4�0�{4@��^���!?cc~��@�m���ٿ��}�3�@4�0�{4@��^���!?cc~��@	�ς��ٿe����g�@W/E4@u���;�!?PW9����@	�ς��ٿe����g�@W/E4@u���;�!?PW9����@	�ς��ٿe����g�@W/E4@u���;�!?PW9����@���1)�ٿ�Ht@�b�@[\�~"4@(TPk�!?�;����@���1)�ٿ�Ht@�b�@[\�~"4@(TPk�!?�;����@���1)�ٿ�Ht@�b�@[\�~"4@(TPk�!?�;����@���1)�ٿ�Ht@�b�@[\�~"4@(TPk�!?�;����@2��9�ٿ���EO�@W��$4@1C!fP�!?͓��K�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@�1��ٿu�L�y�@'��(4@Fe�	y�!?�0�@�@}��#��ٿz�G9��@��}�04@h�;ً�!?���"@?q�y;�ٿn�<b>�@ɭ�j�P4@��N�9�!?wJ\wp�@��I�ٿ�85�m��@V�)a"4@�~R�8�!?��t����@���i/�ٿ�� P4�@`���y4@��J�9�!?m�𜣕@���i/�ٿ�� P4�@`���y4@��J�9�!?m�𜣕@���i/�ٿ�� P4�@`���y4@��J�9�!?m�𜣕@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@�t_)E�ٿO��Ǫ7�@���ܔ
4@��U�v�!?W����ƕ@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@P(�� �ٿ��'����@~��84@c��h<�!??��-�P�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@�Q[	]�ٿ=ɞ��@&�iY��3@�}���!?#��J�@Z��Ѣ�ٿ��Wf��@ƣ��N4@j"x�{�!?����@��[i��ٿ�<9���@��"��=4@�$M틐!?,Z(��@��[i��ٿ�<9���@��"��=4@�$M틐!?,Z(��@��[i��ٿ�<9���@��"��=4@�$M틐!?,Z(��@R��\��ٿs�V��@_�D�� 4@��^i�!?g?��Z��@R��\��ٿs�V��@_�D�� 4@��^i�!?g?��Z��@R��\��ٿs�V��@_�D�� 4@��^i�!?g?��Z��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@;!�&��ٿ'���c��@,�*�%4@�9J(�!?
%f>��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@��N�ٿ�d�ِ�@������3@m��U�!?��Ǵ��@
R��n�ٿ��tb�@�l�E��3@<:$j�!?�����@
R��n�ٿ��tb�@�l�E��3@<:$j�!?�����@
R��n�ٿ��tb�@�l�E��3@<:$j�!?�����@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@	%��ٿ!�LfO��@=�Ƹ4@"�o1��!?k���@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@���d�ٿY�y��@t@��4@� �<d�!?"����ٕ@�,��j�ٿR��ܙ��@��i$�Z4@�ִ���!?8�X�$�@5@�aޛٿ8�����@�n� 4@�o���!?�-r!ܶ�@5@�aޛٿ8�����@�n� 4@�o���!?�-r!ܶ�@0Zč�ٿ��+�O��@!o�"4@QO󲀐!?�>��@0Zč�ٿ��+�O��@!o�"4@QO󲀐!?�>��@"(^��ٿ~����@Q�(CEG4@r��x�!?w.A���@"(^��ٿ~����@Q�(CEG4@r��x�!?w.A���@"(^��ٿ~����@Q�(CEG4@r��x�!?w.A���@F���ٿĚɦ���@���c�4@�&F�C�!?E����@F���ٿĚɦ���@���c�4@�&F�C�!?E����@F���ٿĚɦ���@���c�4@�&F�C�!?E����@�}>J�ٿ ��o�9�@��?s�3@@C�Z(�!?��L[a�@�}>J�ٿ ��o�9�@��?s�3@@C�Z(�!?��L[a�@�)\3�ٿP{�:r�@��犹4@o��F�!?�a�a��@�)\3�ٿP{�:r�@��犹4@o��F�!?�a�a��@��Z`��ٿao����@���P�Y4@!?0��!?�('n�@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@��9t��ٿ�m����@w,��Hw4@���3Ɛ!?"� ���@�T���ٿ���{�C�@�K$Ej�4@��w�!?U@��@�T���ٿ���{�C�@�K$Ej�4@��w�!?U@��@�T���ٿ���{�C�@�K$Ej�4@��w�!?U@��@�T���ٿ���{�C�@�K$Ej�4@��w�!?U@��@��H��ٿ<O�N��@|�a�-X4@�?���!?-d����@�O#��ٿ7��f�!�@��փG44@T�Vb�!?��w�=Z�@��f6�ٿS����@�S����3@q3*�!?tԾK�@kƈ��ٿ��)��K�@�XC���3@����!?��,��@kƈ��ٿ��)��K�@�XC���3@����!?��,��@?�Q�ˣٿ��|�*�@J����3@V�{�!?t�� >��@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@Qp�=��ٿy/T���@�H��x�3@Ƕ-ߏ!?D�L�@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@m+�gٿ �Z]8y�@�$}��4@�!�oC�!?�e��@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@��I	�ٿ�Z� ��@0���"&4@��>�}�!?o)!k:Е@*'�Ά�ٿ���S6��@��iy,+4@�a� -�!?"~� ���@*'�Ά�ٿ���S6��@��iy,+4@�a� -�!?"~� ���@*'�Ά�ٿ���S6��@��iy,+4@�a� -�!?"~� ���@�Ï��ٿ�L_�K@�@!,�G)4@��ϽC�!?q/!e�f�@�R*�ٿ�����_�@�>�"'4@��"3�!?5o�A���@�R*�ٿ�����_�@�>�"'4@��"3�!?5o�A���@�R*�ٿ�����_�@�>�"'4@��"3�!?5o�A���@�R*�ٿ�����_�@�>�"'4@��"3�!?5o�A���@p�̝ٿ�&���@�4U-4@C�f���!?�*q��@p�̝ٿ�&���@�4U-4@C�f���!?�*q��@��{�ڟٿ{3���@/@�T�4@J�$$�!?�����7�@�%�/D�ٿ����@�|�ҏ=4@3����!?��fu�,�@�%�/D�ٿ����@�|�ҏ=4@3����!?��fu�,�@
2P!��ٿ29c)���@� }�4@ecp���!?Դ3Ee�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@��m�Νٿ���_��@��xN4@65d�W�!?�dx��s�@�^��Νٿ,��=_�@�xo�M4@�����!?�j㤏�@�^��Νٿ,��=_�@�xo�M4@�����!?�j㤏�@���#�ٿ�T�0��@�cw^4@��� ��!?&�P�8�@���#�ٿ�T�0��@�cw^4@��� ��!?&�P�8�@F}�ٿ�gU(�@�B#wU4@����m�!?H�Adٕ@F}�ٿ�gU(�@�B#wU4@����m�!?H�Adٕ@F}�ٿ�gU(�@�B#wU4@����m�!?H�Adٕ@F}�ٿ�gU(�@�B#wU4@����m�!?H�Adٕ@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@�x�.�ٿ�)K��@b�:4@i�3C�!?��u��@��CK�ٿ�2O<{��@��/�iC4@ʓ���!?�����@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@:"֛�ٿ83�7d��@2�;".4@�� �!?/rv�Ε@={��D�ٿ�'�1|��@�tԽi04@Hc=j|�!?哸�滕@~��x��ٿ��c��@���4@����!?˖�0;�@~��x��ٿ��c��@���4@����!?˖�0;�@~��x��ٿ��c��@���4@����!?˖�0;�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@t�8/�ٿ;L_�@o�3��3@�!�
�!?!&� -�@�����ٿԀ��"��@��4*:(4@�E�͵�!?��r��@�����ٿԀ��"��@��4*:(4@�E�͵�!?��r��@�����ٿԀ��"��@��4*:(4@�E�͵�!?��r��@�����ٿԀ��"��@��4*:(4@�E�͵�!?��r��@�����ٿԀ��"��@��4*:(4@�E�͵�!?��r��@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�J�R��ٿ�J����@�E���.4@D����!?���V�ؕ@�����ٿz	JHX�@�1b�=�3@`�W3�!?< ����@�����ٿz	JHX�@�1b�=�3@`�W3�!?< ����@Q�X�<�ٿ��Fv04�@��`[��3@y�4��!?�5��ǵ�@Q�X�<�ٿ��Fv04�@��`[��3@y�4��!?�5��ǵ�@
WX\�ٿv�eUj�@0L�!\�3@©��@�!?{��;^0�@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@z���ٿ��TQ��@�J�3��3@��|�U�!?94>=ߕ@�n� Ϛٿ��jd-�@T��N��3@Xs��!?�KdP�ƕ@�n� Ϛٿ��jd-�@T��N��3@Xs��!?�KdP�ƕ@�>��ٿ��jȘ�@��2�3@�N��!?�!0�ו@#_`��ٿU�vWG��@mN�d4@b��e�!?�J��d�@#_`��ٿU�vWG��@mN�d4@b��e�!?�J��d�@i�(*�ٿ=`s����@{�>���3@Z�ѰE�!?��5ɫ@i�(*�ٿ=`s����@{�>���3@Z�ѰE�!?��5ɫ@i�(*�ٿ=`s����@{�>���3@Z�ѰE�!?��5ɫ@�'ͪ��ٿ��u�t�@E�1���3@ފFm9�!?)�C3��@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@Tq��ٿ�=�����@�����4@�㪼�!?6iK�DЕ@D&�a�ٿ���S���@���:4@{�����!?�S8��@:S���ٿl��f�i�@+-�lp4@���!?ɾ:�5�@:S���ٿl��f�i�@+-�lp4@���!?ɾ:�5�@� �7�ٿ�6��K�@y�ok�94@ mv(��!?,�?��ŕ@� �7�ٿ�6��K�@y�ok�94@ mv(��!?,�?��ŕ@� �7�ٿ�6��K�@y�ok�94@ mv(��!?,�?��ŕ@� �7�ٿ�6��K�@y�ok�94@ mv(��!?,�?��ŕ@� �7�ٿ�6��K�@y�ok�94@ mv(��!?,�?��ŕ@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�M���ٿУ;2@��@�H϶O14@M�1��!?�ۈr֕@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@�ie�ٿ�.��&��@��-ł4@+y�!?E�s��@EM��ݖٿ��@�NZ�@2�D��4@	��A9�!?�'�YPՕ@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@BE��
�ٿ���m̗�@'�D�3@��]~�!?JcY�L�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@����S�ٿ^����@�gR�w)4@���Ő!?��-nW�@b?�a�ٿ��QX��@%u�"4@�Ox=�!?�0��bR�@b?�a�ٿ��QX��@%u�"4@�Ox=�!?�0��bR�@b?�a�ٿ��QX��@%u�"4@�Ox=�!?�0��bR�@b?�a�ٿ��QX��@%u�"4@�Ox=�!?�0��bR�@�8s�ٿn�����@!�F.4@nU��!?b�6VY%�@5�0l��ٿ%�s��@��⧆4@X-r��!?���y�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�v�	�ٿ�{N����@�x�4@�sĐ!?��=�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@�I?�ќٿ�TXԾy�@�N��64@_��=�!?W~��N+�@y$bL؜ٿ>��P@��@�>.�4@����!?"�F��@��v6�ٿ��q��@�u%x��3@ׯ��!?��Ѫ�ٕ@�w�0�ٿ���u���@�����3@��N�>�!?�����@���P�ٿ�a�)��@Y�c�64@��2M�!?e���@���P�ٿ�a�)��@Y�c�64@��2M�!?e���@���P�ٿ�a�)��@Y�c�64@��2M�!?e���@���P�ٿ�a�)��@Y�c�64@��2M�!?e���@����y�ٿ"����@�]�e�4@�N5X�!?$�d[�5�@����y�ٿ"����@�]�e�4@�N5X�!?$�d[�5�@����y�ٿ"����@�]�e�4@�N5X�!?$�d[�5�@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@��ҟٿ'lf�@�{oZ�4@"��5�!?�N]�ؕ@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@(iG�ٿ��2��3�@p����3@M.��v�!?�+��J3�@T=k���ٿTv!�b�@V�V���3@�����!?@	��k�@T=k���ٿTv!�b�@V�V���3@�����!?@	��k�@T=k���ٿTv!�b�@V�V���3@�����!?@	��k�@̄˕ٿ �t=�|�@�΁�a�3@2<9뤐!?4~<��;�@̄˕ٿ �t=�|�@�΁�a�3@2<9뤐!?4~<��;�@̄˕ٿ �t=�|�@�΁�a�3@2<9뤐!?4~<��;�@̄˕ٿ �t=�|�@�΁�a�3@2<9뤐!?4~<��;�@̄˕ٿ �t=�|�@�΁�a�3@2<9뤐!?4~<��;�@~����ٿ��A\��@�瓘�3@�J]]ː!?_�?1��@~����ٿ��A\��@�瓘�3@�J]]ː!?_�?1��@~����ٿ��A\��@�瓘�3@�J]]ː!?_�?1��@~����ٿ��A\��@�瓘�3@�J]]ː!?_�?1��@~����ٿ��A\��@�瓘�3@�J]]ː!?_�?1��@�L�^�ٿO��,��@�G>m��3@أm��!?�'��Y��@�L�^�ٿO��,��@�G>m��3@أm��!?�'��Y��@�L�^�ٿO��,��@�G>m��3@أm��!?�'��Y��@�L�^�ٿO��,��@�G>m��3@أm��!?�'��Y��@��0�/�ٿ�T�t|��@J�6ĸ3@��5fƐ!?8�Jޕ@��0�/�ٿ�T�t|��@J�6ĸ3@��5fƐ!?8�Jޕ@��0�/�ٿ�T�t|��@J�6ĸ3@��5fƐ!?8�Jޕ@��0�/�ٿ�T�t|��@J�6ĸ3@��5fƐ!?8�Jޕ@ ����ٿ���ݥ�@���8C�3@�G�C�!?b��5Τ�@ ����ٿ���ݥ�@���8C�3@�G�C�!?b��5Τ�@ ����ٿ���ݥ�@���8C�3@�G�C�!?b��5Τ�@ ����ٿ���ݥ�@���8C�3@�G�C�!?b��5Τ�@��k��ٿ����@�^�3@���eO�!?F;2�h֕@9�' �ٿS��0�@������3@��R�!?�9�����@9�' �ٿS��0�@������3@��R�!?�9�����@
Q^�'�ٿf/�wh��@;t�9��3@)���Đ!?�Xk��@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�J�ʚٿ���1��@��b�
4@tZ?��!?!��QlՕ@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@�{S��ٿ��a���@���7�4@ފA!��!?�j?�@eq�y�ٿ<M;���@��gڷ�3@����!?�e9����@`Z֓h�ٿr�J���@(�dU;.4@vQ�F9�!?:�3�(��@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@M4�)_�ٿ��G%�@�YL6�3@��?U�!?����@���ٿ�ߛ9)�@�d�4@ę�c<�!?�l���@���ٿ�ߛ9)�@�d�4@ę�c<�!?�l���@�GF*9�ٿ��B��@#\ߧiV4@t\���!?oQn�ܕ@�GF*9�ٿ��B��@#\ߧiV4@t\���!?oQn�ܕ@��f(�ٿ.��\ ��@��=4@<��7g�!?08�n�ĕ@��f(�ٿ.��\ ��@��=4@<��7g�!?08�n�ĕ@��f(�ٿ.��\ ��@��=4@<��7g�!?08�n�ĕ@��f(�ٿ.��\ ��@��=4@<��7g�!?08�n�ĕ@��f(�ٿ.��\ ��@��=4@<��7g�!?08�n�ĕ@�^ʇa�ٿ�gB���@Sܲ�4@q�B���!?����Z�@�T�?�ٿ"�����@Iv?�4@R�j��!?�.��H�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@Y�RI�ٿ�0<2ک�@��<�G4@]G����!?鉜�t�@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@�j|��ٿ�x*���@�����3@�~�!?ѩ ���@Nq���ٿ�p��+�@+u�u<4@{��#q�!?�[Z�@Nq���ٿ�p��+�@+u�u<4@{��#q�!?�[Z�@Nq���ٿ�p��+�@+u�u<4@{��#q�!?�[Z�@�.1~�ٿ�p�=�@���G4@["ԍҐ!?i'���ʕ@�.1~�ٿ�p�=�@���G4@["ԍҐ!?i'���ʕ@������ٿ.�#/��@����4@0fB�!?ڵ�����@ǰ"�ٿG#�����@m��E+4@eLa�3�!?�Gx�@ǰ"�ٿG#�����@m��E+4@eLa�3�!?�Gx�@ǰ"�ٿG#�����@m��E+4@eLa�3�!?�Gx�@ǰ"�ٿG#�����@m��E+4@eLa�3�!?�Gx�@��"�ٿ#{|=�
�@~�I��@4@4�r�!?O��ĩ͕@��"�ٿ#{|=�
�@~�I��@4@4�r�!?O��ĩ͕@��"�ٿ#{|=�
�@~�I��@4@4�r�!?O��ĩ͕@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@ē,WV�ٿ�@��@^����I4@��	�6�!?+�f���@����n�ٿp��81�@��"��4@]����!?]^�&��@� h�p�ٿ�r���E�@;�][�3@o�Lp�!?
�ʐ/�@�?�֞ٿ;�kP,��@�%�iU4@�0�T�!?��/o0�@�?�֞ٿ;�kP,��@�%�iU4@�0�T�!?��/o0�@�?�֞ٿ;�kP,��@�%�iU4@�0�T�!?��/o0�@�?�֞ٿ;�kP,��@�%�iU4@�0�T�!?��/o0�@��ѥ�ٿWD5;�@9�\��3@�{��L�!?��?�r�@��ѥ�ٿWD5;�@9�\��3@�{��L�!?��?�r�@��ѥ�ٿWD5;�@9�\��3@�{��L�!?��?�r�@��ځ9�ٿtܥ���@����G-4@\��0�!?�)st��@��ځ9�ٿtܥ���@����G-4@\��0�!?�)st��@��ځ9�ٿtܥ���@����G-4@\��0�!?�)st��@��3��ٿ�X�4�@��j�W"4@j�m
�!?���m��@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@)u�Z"�ٿ�ݟ���@8�ܯ�4@?q�4;�!?��G�4�@�堛ٿxr�Q���@H�c��4@ﭻ��!?��2dQӕ@�堛ٿxr�Q���@H�c��4@ﭻ��!?��2dQӕ@�堛ٿxr�Q���@H�c��4@ﭻ��!?��2dQӕ@��`]�ٿY�-�/�@�j(���3@����1�!?T[��{��@��`]�ٿY�-�/�@�j(���3@����1�!?T[��{��@���i��ٿ��V��@����3@6��e�!?m'r5�@���i��ٿ��V��@����3@6��e�!?m'r5�@���i��ٿ��V��@����3@6��e�!?m'r5�@���i��ٿ��V��@����3@6��e�!?m'r5�@���i��ٿ��V��@����3@6��e�!?m'r5�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@���9��ٿbB
��@P�o'4@a�CB�!?a!߰!>�@oh��K�ٿ�Wm��@�����4@r��!�!?	a��7�@oh��K�ٿ�Wm��@�����4@r��!�!?	a��7�@oh��K�ٿ�Wm��@�����4@r��!�!?	a��7�@oh��K�ٿ�Wm��@�����4@r��!�!?	a��7�@D͋���ٿ��%��@�9��4@�����!?��F~�@��n��ٿ�� s�@M�4�14@_��dߏ!?|��9���@��H�!�ٿ8E2B�/�@nHF%p/4@�md��!?ӵ)���@��H�!�ٿ8E2B�/�@nHF%p/4@�md��!?ӵ)���@��H�!�ٿ8E2B�/�@nHF%p/4@�md��!?ӵ)���@��= ��ٿDe�Ο�@��4@ �-�܏!?	��L���@��= ��ٿDe�Ο�@��4@ �-�܏!?	��L���@��= ��ٿDe�Ο�@��4@ �-�܏!?	��L���@��= ��ٿDe�Ο�@��4@ �-�܏!?	��L���@��= ��ٿDe�Ο�@��4@ �-�܏!?	��L���@Q��;�ٿL@���@�� �3[4@���@�!?�~����@Q��;�ٿL@���@�� �3[4@���@�!?�~����@Q��;�ٿL@���@�� �3[4@���@�!?�~����@Q��;�ٿL@���@�� �3[4@���@�!?�~����@Q��;�ٿL@���@�� �3[4@���@�!?�~����@��t�ٿ�lZ�5�@�k�W{4@��uv#�!?����j4�@��t�ٿ�lZ�5�@�k�W{4@��uv#�!?����j4�@G���W�ٿ)�(>�@2���й4@LE�4�!?{'\�*�@G���W�ٿ)�(>�@2���й4@LE�4�!?{'\�*�@G���W�ٿ)�(>�@2���й4@LE�4�!?{'\�*�@G���W�ٿ)�(>�@2���й4@LE�4�!?{'\�*�@G���W�ٿ)�(>�@2���й4@LE�4�!?{'\�*�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@��g8�ٿk_ƀ�s�@w��V%4@M���"�!?��v�B"�@���X�ٿ�z�!�&�@��1~�4@��?�!?Oȝ���@�u�U�ٿY����@TV����3@V�}�Y�!?��fC�@ꠌkQ�ٿ.�K���@��	��3@���֐!?U���,�@ꠌkQ�ٿ.�K���@��	��3@���֐!?U���,�@ꠌkQ�ٿ.�K���@��	��3@���֐!?U���,�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@S�"���ٿ�jw�r4�@0��r�3@?5���!?�*�të�@���ߕٿ:�@��t�@�
r��74@P���y�!?�MiI��@���ߕٿ:�@��t�@�
r��74@P���y�!?�MiI��@�ͪӛٿ�S��@��EA�I4@ui'��!?���a�@�����ٿ���:[�@R.<��M4@ݻDPH�!?�j��E/�@�����ٿ���:[�@R.<��M4@ݻDPH�!?�j��E/�@�����ٿ���:[�@R.<��M4@ݻDPH�!?�j��E/�@�����ٿ���:[�@R.<��M4@ݻDPH�!?�j��E/�@煖8�ٿ�@D����@g��=L4@���"b�!?B��ոh�@煖8�ٿ�@D����@g��=L4@���"b�!?B��ոh�@煖8�ٿ�@D����@g��=L4@���"b�!?B��ոh�@煖8�ٿ�@D����@g��=L4@���"b�!?B��ոh�@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@g�!j��ٿ���(�@{U��,4@��cg�!?J������@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@ʻr���ٿ	�0iN��@���L;4@�ƹ���!?�o�t֕@j��0�ٿ�{E����@�2�N4@c�q�!?}x6k�˕@j��0�ٿ�{E����@�2�N4@c�q�!?}x6k�˕@j��0�ٿ�{E����@�2�N4@c�q�!?}x6k�˕@�X��!�ٿ�Q4 ���@@�A
4@�=�M&�!?��ȕ@��w-�ٿlH5h+$�@�lK�W4@�b/�0�!?��O\롕@��w-�ٿlH5h+$�@�lK�W4@�b/�0�!?��O\롕@�x����ٿb��WP�@�or�e4@P�]w�!?J=�+���@�x����ٿb��WP�@�or�e4@P�]w�!?J=�+���@�x����ٿb��WP�@�or�e4@P�]w�!?J=�+���@�x����ٿb��WP�@�or�e4@P�]w�!?J=�+���@ Y��p�ٿ̜�.y��@|��a�X4@8N��2�!?�*��Q͕@ Y��p�ٿ̜�.y��@|��a�X4@8N��2�!?�*��Q͕@ Y��p�ٿ̜�.y��@|��a�X4@8N��2�!?�*��Q͕@3=̥ޟٿ��w��(�@����@4@����ʏ!?G��@��e$n�ٿ�u�����@����,4@.䍆�!?�ᩤH�@��e$n�ٿ�u�����@����,4@.䍆�!?�ᩤH�@ۓ���ٿ��V��4�@�碩�4@���Dҏ!?_/*�@ۓ���ٿ��V��4�@�碩�4@���Dҏ!?_/*�@ۓ���ٿ��V��4�@�碩�4@���Dҏ!?_/*�@ۓ���ٿ��V��4�@�碩�4@���Dҏ!?_/*�@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@��� ��ٿ+�ʸ�@�X�S�i4@E��/�!?������@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@=f��H�ٿ^T*��@�73 4@��K��!?�O_Ԇ�@d����ٿj��uJ��@�+�9g;4@OFw`�!?36�4ӻ�@����ٿ66]7Rp�@�� �4@Fn��!?/=�R�|�@����ٿ66]7Rp�@�� �4@Fn��!?/=�R�|�@����ٿ66]7Rp�@�� �4@Fn��!?/=�R�|�@����ٿ66]7Rp�@�� �4@Fn��!?/=�R�|�@8���2�ٿWs}'�
�@��!	%4@�gȄe�!?�1���1�@8���2�ٿWs}'�
�@��!	%4@�gȄe�!?�1���1�@8���2�ٿWs}'�
�@��!	%4@�gȄe�!?�1���1�@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@��J]q�ٿ&R}���@�x�t\#4@�ڦ�D�!?��D��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@{�XS��ٿqVD���@[Qr��14@���M�!?��cD��@s�k��ٿN�A^���@Aiq>4@�ȶn��!?��.�4�@s�k��ٿN�A^���@Aiq>4@�ȶn��!?��.�4�@s�k��ٿN�A^���@Aiq>4@�ȶn��!?��.�4�@s�k��ٿN�A^���@Aiq>4@�ȶn��!?��.�4�@��|M�ٿ�.HhM�@��?�4	4@�g�B�!?����4(�@�X/3��ٿ�P�T�@�x��#4@�R@�E�!?�z㒝��@�X/3��ٿ�P�T�@�x��#4@�R@�E�!?�z㒝��@�X/3��ٿ�P�T�@�x��#4@�R@�E�!?�z㒝��@�mx�Śٿ��"�@}��4@&Nt�D�!?9+e���@�mx�Śٿ��"�@}��4@&Nt�D�!?9+e���@`��ٿ�$]����@���� 4@`�{u�!?��z��@`��ٿ�$]����@���� 4@`�{u�!?��z��@������ٿ7�g�3��@<���3@#���h�!?�a �F��@������ٿ7�g�3��@<���3@#���h�!?�a �F��@������ٿ7�g�3��@<���3@#���h�!?�a �F��@������ٿ7�g�3��@<���3@#���h�!?�a �F��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@�#[-�ٿ��C�� �@*u��4@��b^�!?k�h4��@ԋ����ٿ2r43M��@~d���4@���!?D9,��@ԋ����ٿ2r43M��@~d���4@���!?D9,��@ԋ����ٿ2r43M��@~d���4@���!?D9,��@ԋ����ٿ2r43M��@~d���4@���!?D9,��@�ÙzϜٿ��Q�_�@CQ�4@�_mw��!?ᴭ�@/ۣ��ٿ{��F��@p�:$4@>��#�!?vQ�#)�@/ۣ��ٿ{��F��@p�:$4@>��#�!?vQ�#)�@/ۣ��ٿ{��F��@p�:$4@>��#�!?vQ�#)�@^;SÜٿaju#&�@3��*4@a�E���!?N�mr(�@^;SÜٿaju#&�@3��*4@a�E���!?N�mr(�@^;SÜٿaju#&�@3��*4@a�E���!?N�mr(�@^;SÜٿaju#&�@3��*4@a�E���!?N�mr(�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@YW^��ٿQ0�-3S�@ʠ� y4@�܏5|�!?L�kx	�@�Π��ٿ�D����@F�W84@g�LT�!?Ò�$��@�Π��ٿ�D����@F�W84@g�LT�!?Ò�$��@�Π��ٿ�D����@F�W84@g�LT�!?Ò�$��@#���,�ٿha�Bc��@�Xu�714@r�*"�!?@$Ŀb'�@#���,�ٿha�Bc��@�Xu�714@r�*"�!?@$Ŀb'�@#���,�ٿha�Bc��@�Xu�714@r�*"�!?@$Ŀb'�@#���,�ٿha�Bc��@�Xu�714@r�*"�!?@$Ŀb'�@��&�ٿ��!��@)���4@_Ot�!?{�Fmt>�@G�3�u�ٿlR#���@CoI�J4@�L�)��!?��`	ĕ@G�3�u�ٿlR#���@CoI�J4@�L�)��!?��`	ĕ@׽WYy�ٿaF,���@OE�s��3@0a���!?!�ϱ��@׽WYy�ٿaF,���@OE�s��3@0a���!?!�ϱ��@׽WYy�ٿaF,���@OE�s��3@0a���!?!�ϱ��@׽WYy�ٿaF,���@OE�s��3@0a���!?!�ϱ��@׽WYy�ٿaF,���@OE�s��3@0a���!?!�ϱ��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@G~-0!�ٿ7`=Z&�@�L��4@ K�V�!?w��{��@������ٿ#f��f�@\Z,��4@�'aO+�!?Д|�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@�d_��ٿ,��K��@Z�+�6�3@��Sr�!?ڲ�Ze�@C����ٿ�Q+z�3�@��@j 4@|�0c�!?Z��N�@C����ٿ�Q+z�3�@��@j 4@|�0c�!?Z��N�@C����ٿ�Q+z�3�@��@j 4@|�0c�!?Z��N�@C����ٿ�Q+z�3�@��@j 4@|�0c�!?Z��N�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@o�&=J�ٿ��g��b�@��c���3@��Y(�!?!{O�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@U�Ɏ��ٿ[�Pe��@� �A$�3@J�N�!?c�M�
�@��i���ٿ�fI����@"���/84@z튡��!?����5��@��i���ٿ�fI����@"���/84@z튡��!?����5��@����u�ٿ�~����@���]�4@L�?D]�!?��Y��@����u�ٿ�~����@���]�4@L�?D]�!?��Y��@����u�ٿ�~����@���]�4@L�?D]�!?��Y��@����u�ٿ�~����@���]�4@L�?D]�!?��Y��@����u�ٿ�~����@���]�4@L�?D]�!?��Y��@��7K8�ٿxuJ�~�@���O�@4@U넝�!?�:S ���@��7K8�ٿxuJ�~�@���O�@4@U넝�!?�:S ���@��7K8�ٿxuJ�~�@���O�@4@U넝�!?�:S ���@��7K8�ٿxuJ�~�@���O�@4@U넝�!?�:S ���@qx�C�ٿ�?�G@��@�2)04@�@�u<�!?s*Z��@qx�C�ٿ�?�G@��@�2)04@�@�u<�!?s*Z��@qx�C�ٿ�?�G@��@�2)04@�@�u<�!?s*Z��@�䢔�ٿ��QF�@�Q��2	4@��Uf�!?9�-�?s�@�䢔�ٿ��QF�@�Q��2	4@��Uf�!?9�-�?s�@�Z�Ƅ�ٿ�5((^�@=�;�3@��ҟs�!?0���=l�@�Z�Ƅ�ٿ�5((^�@=�;�3@��ҟs�!?0���=l�@�Z�Ƅ�ٿ�5((^�@=�;�3@��ҟs�!?0���=l�@)�r!<�ٿH�����@(��*�3@��,�!?^�.�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@O��bG�ٿ����Pq�@_jǉY44@���<p�!?�5F�@H�|2��ٿ�'��x�@����!4@�� ��!?�@�ܼ�@H�|2��ٿ�'��x�@����!4@�� ��!?�@�ܼ�@H�|2��ٿ�'��x�@����!4@�� ��!?�@�ܼ�@H�|2��ٿ�'��x�@����!4@�� ��!?�@�ܼ�@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@9r���ٿ�r�pX��@��/��4@�[D�!?7衛ڕ@��vC�ٿb�TBU��@_��v*4@A-!�!?��o�r�@s2}Y�ٿO�ס��@�JG`+>4@���{F�!?|�Y�F�@s2}Y�ٿO�ס��@�JG`+>4@���{F�!?|�Y�F�@s2}Y�ٿO�ס��@�JG`+>4@���{F�!?|�Y�F�@s2}Y�ٿO�ס��@�JG`+>4@���{F�!?|�Y�F�@�j�{�ٿ�����@B$\�/4@�����!?%(\�@]�@�j�{�ٿ�����@B$\�/4@�����!?%(\�@]�@�j�{�ٿ�����@B$\�/4@�����!?%(\�@]�@�j�{�ٿ�����@B$\�/4@�����!?%(\�@]�@�~.���ٿ.u߂���@����$4@��ز�!?,J%�a�@�~.���ٿ.u߂���@����$4@��ز�!?,J%�a�@�~.���ٿ.u߂���@����$4@��ز�!?,J%�a�@�~.���ٿ.u߂���@����$4@��ز�!?,J%�a�@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@޾�pB�ٿBn PQ��@+�F��3@�4�ȏ!?f����@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@k󯹖ٿFQG��%�@���K�3@}/B�.�!?�k@C֕@�2�x�ٿ��VVH�@B�uQ4@��Vn�!?�E��D�@�2�x�ٿ��VVH�@B�uQ4@��Vn�!?�E��D�@Pg
�ٿ�	a%�@�!2�4@$�Eʈ�!?���9^^�@Pg
�ٿ�	a%�@�!2�4@$�Eʈ�!?���9^^�@?�j�ٿu��w��@��bC� 4@��A�!?���-�@?�j�ٿu��w��@��bC� 4@��A�!?���-�@?�j�ٿu��w��@��bC� 4@��A�!?���-�@p_}�y�ٿѡ�I�$�@�v�l9*4@��i<;�!?M�p"Q*�@p_}�y�ٿѡ�I�$�@�v�l9*4@��i<;�!?M�p"Q*�@p_}�y�ٿѡ�I�$�@�v�l9*4@��i<;�!?M�p"Q*�@{�A��ٿ���d}q�@w�64@(�W%��!?o$5`�ؕ@{�A��ٿ���d}q�@w�64@(�W%��!?o$5`�ؕ@{�A��ٿ���d}q�@w�64@(�W%��!?o$5`�ؕ@{�A��ٿ���d}q�@w�64@(�W%��!?o$5`�ؕ@��ٿ��C���@&��N�"4@�{���!?|u��ɕ@��ٿ��C���@&��N�"4@�{���!?|u��ɕ@��ٿ��C���@&��N�"4@�{���!?|u��ɕ@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@t1@��ٿ�o*M�0�@XK�lP4@��`�!?w`Q`�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@[��k��ٿkL�$y%�@����F4@d�m�!?2�6�%�@�G��ٿY ���.�@����)4@�簁#�!? �ع>-�@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�*��m�ٿR���Gl�@��Հ�.4@�?�A�!?e1�ؕ@�1��ٿ><�m��@����4@h#,�!?��VÕ@�1��ٿ><�m��@����4@h#,�!?��VÕ@�Ѽ�ٿ%s	���@r���K4@Uj�&�!?ݐ�O��@iJ��ٿ�_��@��W��m4@g����!?���y�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@��_F�ٿ�ᐓ@2�@1F{d4@�7[:�!?�]EK�@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@�%t�O�ٿ��2�@���}��3@.X��&�!?���T��@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@��ͭ�ٿ%(U;&��@��(Ή�3@��)�G�!?�[����@8=�(�ٿE,9,l�@�
t= 4@��oX�!?XvX{Ӹ�@8=�(�ٿE,9,l�@�
t= 4@��oX�!?XvX{Ӹ�@8=�(�ٿE,9,l�@�
t= 4@��oX�!?XvX{Ӹ�@8=�(�ٿE,9,l�@�
t= 4@��oX�!?XvX{Ӹ�@8=�(�ٿE,9,l�@�
t= 4@��oX�!?XvX{Ӹ�@f=�|�ٿtB����@`���'4@>m2 N�!?��3+�%�@f=�|�ٿtB����@`���'4@>m2 N�!?��3+�%�@f=�|�ٿtB����@`���'4@>m2 N�!?��3+�%�@f=�|�ٿtB����@`���'4@>m2 N�!?��3+�%�@|_���ٿ�w�`�@���G4@B3�}�!?E^1�#f�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@�� '�ٿO0����@Բ�Z'4@��?���!?g���9�@p�oƟٿl7'u�*�@Հ�O;4@s�R�!?uG�?${�@p�oƟٿl7'u�*�@Հ�O;4@s�R�!?uG�?${�@p�oƟٿl7'u�*�@Հ�O;4@s�R�!?uG�?${�@p�oƟٿl7'u�*�@Հ�O;4@s�R�!?uG�?${�@;��k�ٿ��0�b�@'�U�+4@����0�!?"8��3[�@;��k�ٿ��0�b�@'�U�+4@����0�!?"8��3[�@;��k�ٿ��0�b�@'�U�+4@����0�!?"8��3[�@;��k�ٿ��0�b�@'�U�+4@����0�!?"8��3[�@?_W�*�ٿ^��k��@��C{�:4@���a�!?��x�N�@?_W�*�ٿ^��k��@��C{�:4@���a�!?��x�N�@?_W�*�ٿ^��k��@��C{�:4@���a�!?��x�N�@?_W�*�ٿ^��k��@��C{�:4@���a�!?��x�N�@?_W�*�ٿ^��k��@��C{�:4@���a�!?��x�N�@k���ٿC�:<��@헌"�4@w8���!?�rc��@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@w*�@�ٿ[���6�@Qr��4@�v<�!?=Ϳ:�@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@�&ҝp�ٿ>��*��@<؈�'4@���z�!?��$�$��@7�ID[�ٿ�$~�¨�@d
�N>�3@������!?hN��[��@�cء��ٿ#D�j�@�%L1�3@;�og��!?H���zE�@�cء��ٿ#D�j�@�%L1�3@;�og��!?H���zE�@�cء��ٿ#D�j�@�%L1�3@;�og��!?H���zE�@�cء��ٿ#D�j�@�%L1�3@;�og��!?H���zE�@�cء��ٿ#D�j�@�%L1�3@;�og��!?H���zE�@M�gؘٿ�d�1��@�l%LK�3@2)� ��!?�B�N�"�@M�gؘٿ�d�1��@�l%LK�3@2)� ��!?�B�N�"�@n���ƚٿ��[�A��@����G�3@g#��c�!?/�F�ɕ@# u��ٿNos��@�����3@�*��t�!?�����,�@# u��ٿNos��@�����3@�*��t�!?�����,�@������ٿ�C:�=��@$]�
^
4@S�c�V�!?>FC8 ��@������ٿ�C:�=��@$]�
^
4@S�c�V�!?>FC8 ��@c5�'��ٿ���y���@q_�";�3@��&W=�!?�b��/c�@�f�.��ٿ�S�[�@-q}3�3@�&��!?��u�@��6�ѝٿ��V���@���	4@�X��(�!?��n9d�@�Sۜ�ٿ/����@���Ė4@lQ�[�!?�q}�x�@���D�ٿ��D����@J��i4@����z�!?��ˇq��@���D�ٿ��D����@J��i4@����z�!?��ˇq��@���D�ٿ��D����@J��i4@����z�!?��ˇq��@���D�ٿ��D����@J��i4@����z�!?��ˇq��@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@(��:ݝٿ� �I��@%q�ފ�3@�9��z�!?Y���ޕ@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@��E��ٿ8���*�@*_�8��3@Z�)Ő!?,I���@�o�� �ٿ��KXb�@����U?4@��Z���!?�&���@�o�� �ٿ��KXb�@����U?4@��Z���!?�&���@�o�� �ٿ��KXb�@����U?4@��Z���!?�&���@�o�� �ٿ��KXb�@����U?4@��Z���!?�&���@���`�ٿH�}����@_w�� 4@��U��!?܊���'�@���`�ٿH�}����@_w�� 4@��U��!?܊���'�@�񺾌�ٿ��>�nJ�@�b�yD4@Tcv�!? 9��ԕ@�񺾌�ٿ��>�nJ�@�b�yD4@Tcv�!? 9��ԕ@���\��ٿ;@��kj�@Z��`/4@<c��Đ!?�3��oߕ@��.�ٿ{p�'.z�@ƽ��{4@C +�!?SLƶ��@�QH?��ٿ܂�[���@���_P4@j%�ې!?2�$7���@�QH?��ٿ܂�[���@���_P4@j%�ې!?2�$7���@�QH?��ٿ܂�[���@���_P4@j%�ې!?2�$7���@�X���ٿ�ش����@�_�G4@�W*a��!?�\��e��@J��)�ٿ�o�[� �@�?�/4@�qf�!?���1|��@J��)�ٿ�o�[� �@�?�/4@�qf�!?���1|��@J��)�ٿ�o�[� �@�?�/4@�qf�!?���1|��@J��)�ٿ�o�[� �@�?�/4@�qf�!?���1|��@+y���ٿJZ��[�@���k/4@W~|-\�!?0��,l�@+y���ٿJZ��[�@���k/4@W~|-\�!?0��,l�@+y���ٿJZ��[�@���k/4@W~|-\�!?0��,l�@�H���ٿ�zh��8�@1�8E4@���l�!?z[�3ɕ@�H���ٿ�zh��8�@1�8E4@���l�!?z[�3ɕ@���h�ٿda��B^�@�+	1��3@yYn�M�!?��,��&�@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@;!Ӳ�ٿ��:���@�+H��4@���!?L�7<��@���T�ٿ��ҿ�@7�6��3@@���!?8���@���T�ٿ��ҿ�@7�6��3@@���!?8���@�:���ٿ�.G<$L�@ۡ��L�3@�ߊ��!?E{Y ��@�:���ٿ�.G<$L�@ۡ��L�3@�ߊ��!?E{Y ��@!� ��ٿTz�Ӄ�@��R��3@��k �!?+�.[jĕ@y�m\5�ٿ����"�@������3@e0+��!?���&u�@y�m\5�ٿ����"�@������3@e0+��!?���&u�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@v	��ٿX�1|�@�o���3@]I���!?߇�sg�@��]i�ٿ���H��@����K4@Y�
���!?31.���@�/F嘚ٿ�3N�%	�@iL��4@��Ҟ�!?BG���;�@���_ �ٿ���f��@-���2�3@���L&�!?U�� 7�@���_ �ٿ���f��@-���2�3@���L&�!?U�� 7�@�I��!�ٿ��ܿ�v�@ra�s�3@y�A��!?Ր�_D�@�I��!�ٿ��ܿ�v�@ra�s�3@y�A��!?Ր�_D�@�I��!�ٿ��ܿ�v�@ra�s�3@y�A��!?Ր�_D�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@9b��ٿ<�"�f?�@��<un�3@��ԟ��!?�j*y�4�@Or���ٿJ��u�<�@�$��0�3@�ft��!?�d&t���@Or���ٿJ��u�<�@�$��0�3@�ft��!?�d&t���@����Y�ٿ%ƆIN��@��,:4@��Df�!?E�n�ڕ@����Y�ٿ%ƆIN��@��,:4@��Df�!?E�n�ڕ@����Y�ٿ%ƆIN��@��,:4@��Df�!?E�n�ڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@N_x0��ٿ O#��@@C�+'4@M 컐!?��ؘڕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@� �l�ٿ�k�P�@�MfD�.4@�G,��!?P�2sĕ@DL�t!�ٿ7��ܟ7�@|��e,�3@����!?]o�3�@DL�t!�ٿ7��ܟ7�@|��e,�3@����!?]o�3�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@�?�hL�ٿ�Gr��	�@Q�S14@�2N�!?�T4�F�@װ���ٿ��Y���@D�T=�3@p���Ϗ!?��Q�@װ���ٿ��Y���@D�T=�3@p���Ϗ!?��Q�@װ���ٿ��Y���@D�T=�3@p���Ϗ!?��Q�@�ܔĤٿ����Й�@��'+4@���Ǐ!?z!��6��@�ܔĤٿ����Й�@��'+4@���Ǐ!?z!��6��@�ܔĤٿ����Й�@��'+4@���Ǐ!?z!��6��@�ܔĤٿ����Й�@��'+4@���Ǐ!?z!��6��@�6Z��ٿ��eqm%�@[��T4@w�B�]�!?�ʜ�	�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@8�(?��ٿ�`		��@��9�4@���6�!?4�_�"?�@�R�	�ٿ�h��O��@� L$�M4@�j�8�!?� Èݕ@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@=� ���ٿJ��,���@��.�[4@R3�䱐!?)���oU�@�1���ٿ��AW��@s6�~�f4@)�K���!?F�=�$�@�1���ٿ��AW��@s6�~�f4@)�K���!?F�=�$�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�X�=��ٿ����@jmIlN4@��;S��!?u��!�@�D�EX�ٿ�8e�0�@�崙&4@4Yh�t�!?��iF��@�D�EX�ٿ�8e�0�@�崙&4@4Yh�t�!?��iF��@�D�EX�ٿ�8e�0�@�崙&4@4Yh�t�!?��iF��@�D�EX�ٿ�8e�0�@�崙&4@4Yh�t�!?��iF��@�D�EX�ٿ�8e�0�@�崙&4@4Yh�t�!?��iF��@�)�i��ٿ��#'�Y�@�O'Xa�3@$c �!?K͇��ĕ@�)�i��ٿ��#'�Y�@�O'Xa�3@$c �!?K͇��ĕ@Ô�K%�ٿ�TD iS�@uπV��3@>ƙ<ҏ!?6�"ߕ@Ô�K%�ٿ�TD iS�@uπV��3@>ƙ<ҏ!?6�"ߕ@Ô�K%�ٿ�TD iS�@uπV��3@>ƙ<ҏ!?6�"ߕ@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@�f6�ؠٿ֜vH���@���f�4@�^��>�!?��=�@Ņ�2��ٿwY �@�8�E��3@��M9�!?�\�**ݕ@Ņ�2��ٿwY �@�8�E��3@��M9�!?�\�**ݕ@Ņ�2��ٿwY �@�8�E��3@��M9�!?�\�**ݕ@��P�̗ٿ�VO���@�����3@�Oc���!?���In��@��P�̗ٿ�VO���@�����3@�Oc���!?���In��@��P�̗ٿ�VO���@�����3@�Oc���!?���In��@��P�̗ٿ�VO���@�����3@�Oc���!?���In��@��P�̗ٿ�VO���@�����3@�Oc���!?���In��@����k�ٿ��s����@)s-Dr�3@>�r�+�!?�����+�@����k�ٿ��s����@)s-Dr�3@>�r�+�!?�����+�@����k�ٿ��s����@)s-Dr�3@>�r�+�!?�����+�@&��ٿ�H�SWU�@�W���3@���s�!?0mV6!0�@;U,�ٿT�=����@�0_##4@�M�{�!?�S���@�����ٿI*ˡU�@���x24@�ʒ�E�!?`d�ڕ@�����ٿI*ˡU�@���x24@�ʒ�E�!?`d�ڕ@�����ٿI*ˡU�@���x24@�ʒ�E�!?`d�ڕ@�����ٿI*ˡU�@���x24@�ʒ�E�!?`d�ڕ@�����ٿI*ˡU�@���x24@�ʒ�E�!?`d�ڕ@���"��ٿpP��@��	���3@�M��!?w��{���@���"��ٿpP��@��	���3@�M��!?w��{���@���"��ٿpP��@��	���3@�M��!?w��{���@���"��ٿpP��@��	���3@�M��!?w��{���@���"��ٿpP��@��	���3@�M��!?w��{���@���"��ٿpP��@��	���3@�M��!?w��{���@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@o��聜ٿsl��'�@����3@����Z�!?�((����@
�d�יٿ���;L�@����� 4@��ʏ!?m+��Q�@
�d�יٿ���;L�@����� 4@��ʏ!?m+��Q�@
�d�יٿ���;L�@����� 4@��ʏ!?m+��Q�@
!�7�ٿ��p2b��@��$�A4@Y�}^�!?i���@
!�7�ٿ��p2b��@��$�A4@Y�}^�!?i���@
!�7�ٿ��p2b��@��$�A4@Y�}^�!?i���@
!�7�ٿ��p2b��@��$�A4@Y�}^�!?i���@
!�7�ٿ��p2b��@��$�A4@Y�}^�!?i���@��{���ٿiv�fE�@�ʏ�E4@3P�%1�!?�;�0�@��{���ٿiv�fE�@�ʏ�E4@3P�%1�!?�;�0�@��{���ٿiv�fE�@�ʏ�E4@3P�%1�!?�;�0�@��{���ٿiv�fE�@�ʏ�E4@3P�%1�!?�;�0�@��{���ٿiv�fE�@�ʏ�E4@3P�%1�!?�;�0�@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@\�c��ٿ�c[1�M�@����2�3@y�����!? �D����@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@Eڃ}��ٿ�%_���@�oF%�3@����!?~*b��@MPh�5�ٿ���3�@�u#4@l3
��!?&$b@��@MPh�5�ٿ���3�@�u#4@l3
��!?&$b@��@MPh�5�ٿ���3�@�u#4@l3
��!?&$b@��@MPh�5�ٿ���3�@�u#4@l3
��!?&$b@��@MPh�5�ٿ���3�@�u#4@l3
��!?&$b@��@�����ٿ�u���y�@�FY�5 4@X��`�!?��Fõ�@�����ٿ�u���y�@�FY�5 4@X��`�!?��Fõ�@�����ٿ�u���y�@�FY�5 4@X��`�!?��Fõ�@�����ٿ�u���y�@�FY�5 4@X��`�!?��Fõ�@�����ٿ�u���y�@�FY�5 4@X��`�!?��Fõ�@8��G�ٿ�	�/J�@踩��4@�*�n�!?l�אK��@�>�<�ٿy�cd�@4gy�|=4@)�~x�!?�z���d�@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�O��'�ٿ��4a��@ᾷ��4@�d���!?յ�����@�.f2��ٿ���4��@&���� 4@�=-��!?	Ѭ��@�.f2��ٿ���4��@&���� 4@�=-��!?	Ѭ��@�.f2��ٿ���4��@&���� 4@�=-��!?	Ѭ��@��:��ٿ��N�K�@Z��;y4@�����!?��mA�Е@��:��ٿ��N�K�@Z��;y4@�����!?��mA�Е@��:��ٿ��N�K�@Z��;y4@�����!?��mA�Е@��:��ٿ��N�K�@Z��;y4@�����!?��mA�Е@��,�ٿ܌���@��s4@�FMg��!?�B&K햕@��,�ٿ܌���@��s4@�FMg��!?�B&K햕@�?���ٿ���P��@T�x�"4@�Q��!?,��&��@Q���ٿ5M����@���;�3@�5H�|�!?`Dh�@Q���ٿ5M����@���;�3@�5H�|�!?`Dh�@Q���ٿ5M����@���;�3@�5H�|�!?`Dh�@Q���ٿ5M����@���;�3@�5H�|�!?`Dh�@Q���ٿ5M����@���;�3@�5H�|�!?`Dh�@#�#�u�ٿ�K��Y�@��&G��3@�0�"�!?������@���DK�ٿ��}�n��@qN���3@7۪�]�!?r� �2�@f@C�ٿ�6��@0j�(�3@l��
p�!?\��:ٕ@f@C�ٿ�6��@0j�(�3@l��
p�!?\��:ٕ@f@C�ٿ�6��@0j�(�3@l��
p�!?\��:ٕ@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@(i]��ٿ{h3�r�@[F��@64@P�y�s�!?�#m�Z��@�:��ٿ�=&�h�@>�0]4@9|��!?�]PE��@�:��ٿ�=&�h�@>�0]4@9|��!?�]PE��@�:��ٿ�=&�h�@>�0]4@9|��!?�]PE��@�:��ٿ�=&�h�@>�0]4@9|��!?�]PE��@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@�j�墘ٿ�����-�@-���BH4@�}��z�!?u�����@b�p.�ٿ�y�"��@g���'4@hu�"��!?�9>z��@�m�I[�ٿ=���=�@���p4@���ĉ�!?��t�2�@���n��ٿ�b)��R�@x0��w4@�ɓ�y�!?�����@���n��ٿ�b)��R�@x0��w4@�ɓ�y�!?�����@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@���3��ٿ�!ú��@�Y/׀v4@��#^w�!?��x��@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@IBs��ٿ�fA����@kM=xr�4@K4� z�!?fQ��E�@�ݥK�ٿI5���@�#�H�b4@�:�
��!?m����@�ݥK�ٿI5���@�#�H�b4@�:�
��!?m����@�ݥK�ٿI5���@�#�H�b4@�:�
��!?m����@�ݥK�ٿI5���@�#�H�b4@�:�
��!?m����@�ݥK�ٿI5���@�#�H�b4@�:�
��!?m����@8άc��ٿ�"��	�@����{4@��v���!?�qN��@8άc��ٿ�"��	�@����{4@��v���!?�qN��@8άc��ٿ�"��	�@����{4@��v���!?�qN��@(v�zr�ٿ��vmɍ�@��+T�t4@l=7]t�!?�6�\��@�#�ٿG�2\a��@����DI4@TA�U�!?�l�Σr�@�:��
�ٿ����q*�@��
�xM4@THv��!?#�`N̕@�:��
�ٿ����q*�@��
�xM4@THv��!?#�`N̕@�:��
�ٿ����q*�@��
�xM4@THv��!?#�`N̕@P��`�ٿ<Q勰��@����k4@�?�:G�!?�[%���@�HZ{Y�ٿ*�A$��@tm�azq4@��:�U�!?Eb��!�@�HZ{Y�ٿ*�A$��@tm�azq4@��:�U�!?Eb��!�@�HZ{Y�ٿ*�A$��@tm�azq4@��:�U�!?Eb��!�@�HZ{Y�ٿ*�A$��@tm�azq4@��:�U�!?Eb��!�@�HZ{Y�ٿ*�A$��@tm�azq4@��:�U�!?Eb��!�@�G�)�ٿD��S��@��X[�g4@�P�D�!?���3F�@�G�)�ٿD��S��@��X[�g4@�P�D�!?���3F�@0Ŝ���ٿ�
��X�@S8�:44@�%�$m�!?Y	���@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@����d�ٿt�#4�@񂧂�3@5$����!?N�֔ѱ�@buI8
�ٿ�qv�ݯ�@ha٨�3@���y�!??��@��t�D�ٿ|�j���@?$��74@b?j�!?-�Nʢ�@��t�D�ٿ|�j���@?$��74@b?j�!?-�Nʢ�@��t�D�ٿ|�j���@?$��74@b?j�!?-�Nʢ�@��t�D�ٿ|�j���@?$��74@b?j�!?-�Nʢ�@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@S�җ�ٿ�2&�@%�AIP4@R��J��!?�?���@a�w�y�ٿ��Q�.�@l��3�C4@:��Kѐ!?W~.2H��@~����ٿm���N7�@v�]�0K4@s�昝�!?	��Ir�@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@~�2�ٿx������@_c��X>4@�|�W�!?G�W��@�W*�i�ٿwUW���@1Fq�+4@2xt�1�!?���%�k�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@ѭ9�ʜٿ��G�l'�@	$yR.4@FW7�;�!?W�梅�@df9#A�ٿ�@���@c�ֵ�84@'�#(*�!?P_!��x�@df9#A�ٿ�@���@c�ֵ�84@'�#(*�!?P_!��x�@��s".�ٿ$m��e��@���O
4@�I;e�!?�*�S�@��s".�ٿ$m��e��@���O
4@�I;e�!?�*�S�@��s".�ٿ$m��e��@���O
4@�I;e�!?�*�S�@��~B�ٿ8K��,��@�>��$64@�Cm*�!?�ͷMPk�@��~B�ٿ8K��,��@�>��$64@�Cm*�!?�ͷMPk�@��~B�ٿ8K��,��@�>��$64@�Cm*�!?�ͷMPk�@��~B�ٿ8K��,��@�>��$64@�Cm*�!?�ͷMPk�@n��֡ٿ$
ʉ���@�����4@�<mx��!?�~;�"�@n��֡ٿ$
ʉ���@�����4@�<mx��!?�~;�"�@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@IlGy�ٿ|aJZ�Y�@hJ%K�44@�� ���!?����7ݕ@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��ϙ�ٿ�6�0:~�@rK�B4@�[},��!?wuK�>�@��$��ٿ-}���[�@84J�4@B��炐!?|\j�*ؕ@��$��ٿ-}���[�@84J�4@B��炐!?|\j�*ؕ@��$��ٿ-}���[�@84J�4@B��炐!?|\j�*ؕ@��$��ٿ-}���[�@84J�4@B��炐!?|\j�*ؕ@��Q/"�ٿ*��<W��@$��V�3@<A��!?a�*���@��Q/"�ٿ*��<W��@$��V�3@<A��!?a�*���@��Q/"�ٿ*��<W��@$��V�3@<A��!?a�*���@��Q/"�ٿ*��<W��@$��V�3@<A��!?a�*���@��Q/"�ٿ*��<W��@$��V�3@<A��!?a�*���@�y�
�ٿ�%f��@�E?��3@�']I�!?��.ٕ@�y�
�ٿ�%f��@�E?��3@�']I�!?��.ٕ@�9t�I�ٿ��O�@�7f��T4@,;�!?KT��4�@�9t�I�ٿ��O�@�7f��T4@,;�!?KT��4�@�9t�I�ٿ��O�@�7f��T4@,;�!?KT��4�@��imj�ٿ��ݰ���@�ąD;4@��SV�!?_����͕@��imj�ٿ��ݰ���@�ąD;4@��SV�!?_����͕@ ?_�5�ٿf/�ie
�@3U,!�4@4���F�!?��BN��@ ?_�5�ٿf/�ie
�@3U,!�4@4���F�!?��BN��@�b���ٿ������@U�2�5!4@�j�� �!?��"��@�b���ٿ������@U�2�5!4@�j�� �!?��"��@���ٿc�=���@d�[�.4@���'�!?	�d-�5�@���ٿc�=���@d�[�.4@���'�!?	�d-�5�@K���ٿ��ٞ���@����?4@�䦰b�!?�(�֕@ jmC�ٿ��T�3��@��y+4@�p(k�!?Aŗ	�@ jmC�ٿ��T�3��@��y+4@�p(k�!?Aŗ	�@5>tO��ٿZ��74�@�i02	4@���;�!?���鿕@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@;Wd�ٿ���0�@yD4@0�e}�!?�
`ۜ��@U �7ʚٿQ{H����@���!|84@_s�".�!?��3�Ǖ@U �7ʚٿQ{H����@���!|84@_s�".�!?��3�Ǖ@U �7ʚٿQ{H����@���!|84@_s�".�!?��3�Ǖ@�o���ٿ��~@�@��1L�H4@�I��i�!?�l{����@t6�ٿ��i�S�@�*�GK4@A�!?��G��@t6�ٿ��i�S�@�*�GK4@A�!?��G��@t6�ٿ��i�S�@�*�GK4@A�!?��G��@t6�ٿ��i�S�@�*�GK4@A�!?��G��@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@L#�ٿv���"��@Ǖ��NQ4@uD6v�!?|� �
�@�jt���ٿ�h�C�@�/��m4@��p��!?���R�@�jt���ٿ�h�C�@�/��m4@��p��!?���R�@�jt���ٿ�h�C�@�/��m4@��p��!?���R�@�kvژٿ�ԭ-r:�@@h�i4@\=���!?���|���@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@��L �ٿ�h�c�	�@�CB4@��Bt��!?��Ld��@���.�ٿd�K@���@�c��4@(����!?#���&��@���.�ٿd�K@���@�c��4@(����!?#���&��@���.�ٿd�K@���@�c��4@(����!?#���&��@���.�ٿd�K@���@�c��4@(����!?#���&��@���.�ٿd�K@���@�c��4@(����!?#���&��@�Ls`d�ٿ�H��S��@�}Κ�@4@sb��z�!?���J�{�@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@��m���ٿ6�EZw��@��til4@41uA�!?r�{���@���ٿ(E՟�;�@�XQ��4@��_�9�!?g�X�t�@���ٿ(E՟�;�@�XQ��4@��_�9�!?g�X�t�@���ٿ(E՟�;�@�XQ��4@��_�9�!?g�X�t�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�B�ϲ�ٿg����
�@�7��Q4@��N0.�!? �L"�O�@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@�ޑ�R�ٿ��v����@����64@��#��!??����ƕ@r��ٿ�����@)e2�J4@)�A��!?���s�U�@Vi��A�ٿ�4����@�$.׽�3@�ڳ�!?�����@Vi��A�ٿ�4����@�$.׽�3@�ڳ�!?�����@Vi��A�ٿ�4����@�$.׽�3@�ڳ�!?�����@Vi��A�ٿ�4����@�$.׽�3@�ڳ�!?�����@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@��G�l�ٿH!��@�I"��<4@��=�!?_A��	�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@{gu���ٿ$V�����@;�fԑ*4@
��ǯ�!?wB���8�@��ث�ٿ4�(A���@���x�&4@N�.n�!?W�r�@��ث�ٿ4�(A���@���x�&4@N�.n�!?W�r�@��ث�ٿ4�(A���@���x�&4@N�.n�!?W�r�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@JD�0��ٿN���_�@��EA�H4@�w�T�!?)���~�@�ڌz �ٿY7+��@a�1ujc4@ãh���!?ON��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@Z�O#�ٿXf�I���@ȭ��Q4@p�a�!?�vO��@@r����ٿyGEqǠ�@X�����3@ oN�!?��n�/�@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@bJ;�ٿ�|��@�z�3@#�ʁ�!?�޾%��@��h�B�ٿŖ�!�;�@>�24@��Ա�!?�G� ��@��h�B�ٿŖ�!�;�@>�24@��Ա�!?�G� ��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@@w�f�ٿ�.�I��@W���;4@yX?8�!?m�Sh��@9��ٿ�?�����@s��8�4@�&�3�!?�S� �9�@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@mv�_�ٿl'5�3G�@t�x�-4@8a�9�!?9��1��@�`�D��ٿ��u�p�@ׇ�
�#4@�~ �A�!?�:^��@�`�D��ٿ��u�p�@ׇ�
�#4@�~ �A�!?�:^��@�`�D��ٿ��u�p�@ׇ�
�#4@�~ �A�!?�:^��@�;f�:�ٿ_o�]��@���54@�2g{F�!?��d��@�;f�:�ٿ_o�]��@���54@�2g{F�!?��d��@fN�� �ٿ�à��F�@���u�4@|Ǉ:�!?<�t��@fN�� �ٿ�à��F�@���u�4@|Ǉ:�!?<�t��@fN�� �ٿ�à��F�@���u�4@|Ǉ:�!?<�t��@fN�� �ٿ�à��F�@���u�4@|Ǉ:�!?<�t��@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@����ٿ��	�Q��@�u�24@��J.�!?+����@P'ú�ٿ��'�@z(�+4@����!?����@P'ú�ٿ��'�@z(�+4@����!?����@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@��@e�ٿyo�����@�~z��4@dנZQ�!?�O��]�@fO����ٿ���}���@���4@55rd�!?X%����@fO����ٿ���}���@���4@55rd�!?X%����@fO����ٿ���}���@���4@55rd�!?X%����@V�Ġٿ}ߋ�.�@�����4@U ���!?��
���@_�a���ٿ�e�Nb~�@���A�4@\�$=��!?xEm����@_�a���ٿ�e�Nb~�@���A�4@\�$=��!?xEm����@_�a���ٿ�e�Nb~�@���A�4@\�$=��!?xEm����@_�a���ٿ�e�Nb~�@���A�4@\�$=��!?xEm����@_�a���ٿ�e�Nb~�@���A�4@\�$=��!?xEm����@��Jw��ٿ!��WX�@�Si��3@�Q+p7�!?E��:땕@��Jw��ٿ!��WX�@�Si��3@�Q+p7�!?E��:땕@�*�N�ٿ��Q�#'�@�}�H4@B�R�@�!? rf�h�@�*�N�ٿ��Q�#'�@�}�H4@B�R�@�!? rf�h�@�*�N�ٿ��Q�#'�@�}�H4@B�R�@�!? rf�h�@�*�N�ٿ��Q�#'�@�}�H4@B�R�@�!? rf�h�@fv�zŞٿ|��b��@w��R��3@�7hX�!?��2]y{�@fv�zŞٿ|��b��@w��R��3@�7hX�!?��2]y{�@fv�zŞٿ|��b��@w��R��3@�7hX�!?��2]y{�@����Q�ٿ��]x��@P\�[�3@$56ٛ�!?ҳ��ൕ@����Q�ٿ��]x��@P\�[�3@$56ٛ�!?ҳ��ൕ@ۈ`�ٿ��k���@+�����3@���)Z�!?����@ۈ`�ٿ��k���@+�����3@���)Z�!?����@ۈ`�ٿ��k���@+�����3@���)Z�!?����@ۈ`�ٿ��k���@+�����3@���)Z�!?����@ۈ`�ٿ��k���@+�����3@���)Z�!?����@c/\k��ٿv�A�}�@3��>��3@�bSj��!?a:��W֕@�|AB�ٿ��ԓPy�@q�b��3@E��ݟ�!?�T;#���@�|AB�ٿ��ԓPy�@q�b��3@E��ݟ�!?�T;#���@�|AB�ٿ��ԓPy�@q�b��3@E��ݟ�!?�T;#���@�|AB�ٿ��ԓPy�@q�b��3@E��ݟ�!?�T;#���@�|AB�ٿ��ԓPy�@q�b��3@E��ݟ�!?�T;#���@���K�ٿ.3߉���@z
��3@��{�!?L��YL�@���K�ٿ.3߉���@z
��3@��{�!?L��YL�@�E���ٿI�f?�T�@#�e��4@3~O��!?m
<ؕ@�E���ٿI�f?�T�@#�e��4@3~O��!?m
<ؕ@�E���ٿI�f?�T�@#�e��4@3~O��!?m
<ؕ@�E���ٿI�f?�T�@#�e��4@3~O��!?m
<ؕ@�E���ٿI�f?�T�@#�e��4@3~O��!?m
<ؕ@5�a��ٿ�`�>V��@w�X4@f�+W^�!?���!;�@5�a��ٿ�`�>V��@w�X4@f�+W^�!?���!;�@5�a��ٿ�`�>V��@w�X4@f�+W^�!?���!;�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��Pk�ٿ�Ii��@%�J��3@N��^�!?rp�1�@��r�W�ٿګM���@��{�&�3@A�!�!?��`�PI�@��r�W�ٿګM���@��{�&�3@A�!�!?��`�PI�@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@�\����ٿs8��AL�@:m*p4@�4,ޏ!?�*��@q��ܠٿ�S+��
�@��2DR4@[��W��!?,��mv��@q��ܠٿ�S+��
�@��2DR4@[��W��!?,��mv��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@�Z�;>�ٿ��-�1��@��24@�|��!?H��!s��@��t�ٿ/������@S)0��N4@�H���!?�(����@��^��ٿ+���@�s��D)4@E6~狐!?�;����@Z$G$ךٿ>��X��@��p�R�3@k�lB{�!?>t7#� �@Z$G$ךٿ>��X��@��p�R�3@k�lB{�!?>t7#� �@Z$G$ךٿ>��X��@��p�R�3@k�lB{�!?>t7#� �@�`^�ٿ��e&y�@��5ZN 4@1;����!?���5C̕@�`^�ٿ��e&y�@��5ZN 4@1;����!?���5C̕@�`^�ٿ��e&y�@��5ZN 4@1;����!?���5C̕@�`^�ٿ��e&y�@��5ZN 4@1;����!?���5C̕@�`^�ٿ��e&y�@��5ZN 4@1;����!?���5C̕@u�-°�ٿ����*�@��
/4@��rƐ!?�i�!#ܕ@u�-°�ٿ����*�@��
/4@��rƐ!?�i�!#ܕ@u�-°�ٿ����*�@��
/4@��rƐ!?�i�!#ܕ@u�-°�ٿ����*�@��
/4@��rƐ!?�i�!#ܕ@�ke���ٿ^��F�i�@�l.�174@6;Y���!?^�g���@�ke���ٿ^��F�i�@�l.�174@6;Y���!?^�g���@�ke���ٿ^��F�i�@�l.�174@6;Y���!?^�g���@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@+�l)�ٿL�l�K�@-�F�24@ؽ�⏐!?�� +�@��NL��ٿ��>��@�-C4@T�"��!?�Y1Qk�@��NL��ٿ��>��@�-C4@T�"��!?�Y1Qk�@��NL��ٿ��>��@�-C4@T�"��!?�Y1Qk�@��NL��ٿ��>��@�-C4@T�"��!?�Y1Qk�@��NL��ٿ��>��@�-C4@T�"��!?�Y1Qk�@�5h�u�ٿw����,�@�7�H?4@Z�nH�!?���풖@�5h�u�ٿw����,�@�7�H?4@Z�nH�!?���풖@�5h�u�ٿw����,�@�7�H?4@Z�nH�!?���풖@��)��ٿ%fWҨO�@�d�h 4@
*��V�!?�¶-�@��)��ٿ%fWҨO�@�d�h 4@
*��V�!?�¶-�@��)��ٿ%fWҨO�@�d�h 4@
*��V�!?�¶-�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@���w*�ٿ�?�:��@7y4@�+�I1�!?*pr(�@��Df�ٿej�B�@�@k޹_4@^�ͣP�!?O[+�ݕ@��Df�ٿej�B�@�@k޹_4@^�ͣP�!?O[+�ݕ@���̝�ٿ�i=��@fF�	&4@�(B��!?����s�@���̝�ٿ�i=��@fF�	&4@�(B��!?����s�@���̝�ٿ�i=��@fF�	&4@�(B��!?����s�@���̝�ٿ�i=��@fF�	&4@�(B��!?����s�@���̝�ٿ�i=��@fF�	&4@�(B��!?����s�@)��>��ٿ��+��@l��wS�3@c�J�!?�c�4)?�@*
�q�ٿz]A���@��4�<4@������!?)�6 G�@*
�q�ٿz]A���@��4�<4@������!?)�6 G�@*
�q�ٿz]A���@��4�<4@������!?)�6 G�@b@�V�ٿ>�G�Y�@���^4@M�NW��!?y�Q���@TJNÚٿ���4���@wb��4@^@��!?�u�%�N�@TJNÚٿ���4���@wb��4@^@��!?�u�%�N�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@R�%4�ٿ�U�Q��@�:�]4@�?:E�!?�56!n�@�Q���ٿ-�zw�5�@tP��3@�0��@�!?���6�<�@�Q���ٿ-�zw�5�@tP��3@�0��@�!?���6�<�@�Q���ٿ-�zw�5�@tP��3@�0��@�!?���6�<�@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��1�ؠٿ����i�@�>I�4@�P�@s�!?�u7Z���@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@��~4D�ٿ���ʩZ�@}'���4@ПKH�!?^I�M�@	[�ҚٿE?�|Jm�@#�]P^4@?|T+�!?(|���S�@	[�ҚٿE?�|Jm�@#�]P^4@?|T+�!?(|���S�@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@��P@��ٿ�R�g�b�@��J�f�3@�ExZ��!?K;Y�ו@ЃMK�ٿЬ��T�@�y�_Q4@�+:�N�!? x����@��z'�ٿ��� �p�@�*Q84@�ƙ�_�!?�Kg@WB�@FODĤٿSn]�_�@�-�<�3@f���D�!?�.��� �@�v���ٿi)�_2�@�:�[`N4@����;�!?��W'0Õ@���lA�ٿ�m���@��E��*4@�sr�P�!?�[�9:l�@���lA�ٿ�m���@��E��*4@�sr�P�!?�[�9:l�@���lA�ٿ�m���@��E��*4@�sr�P�!?�[�9:l�@���lA�ٿ�m���@��E��*4@�sr�P�!?�[�9:l�@��#9�ٿ����}�@d���<4@n:&W��!?�.oR�@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@��A��ٿ��� ��@̘ b 4@L���(�!??�����@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@.���ٿ�& ��@�|�� 4@��Ba�!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@rwn��ٿ!s�- ��@ڪ� 4@`"����!?������@ �,���ٿ2� 0 ��@Cy�m 4@f����!?����@ �,���ٿ2� 0 ��@Cy�m 4@f����!?����@e�2<��ٿ<�D ��@���P 4@�@M=�!?<5���@�|�L��ٿ���N ��@}X� 4@� ��,�!?1�����@�|�L��ٿ���N ��@}X� 4@� ��,�!?1�����@k����ٿ��\ ��@Cw}� 4@�<f��!?]5���@k����ٿ��\ ��@Cw}� 4@�<f��!?]5���@L� ��ٿ�1J\ ��@��� 4@[�r9��!?ID����@L� ��ٿ�1J\ ��@��� 4@[�r9��!?ID����@L� ��ٿ�1J\ ��@��� 4@[�r9��!?ID����@L� ��ٿ�1J\ ��@��� 4@[�r9��!?ID����@�qT��ٿ���W ��@uZe� 4@dLwrq�!?]�I���@����ٿ�xLb ��@�o�D 4@�`k�3�!?�+{���@����ٿ�xLb ��@�o�D 4@�`k�3�!?�+{���@����ٿ�xLb ��@�o�D 4@�`k�3�!?�+{���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@�!=+��ٿ�a�U ��@02A 4@��H�c�!?3M���@F{N���ٿ۝*I ��@�I� 4@���V�!?������@F{N���ٿ۝*I ��@�I� 4@���V�!?������@F{N���ٿ۝*I ��@�I� 4@���V�!?������@F{N���ٿ۝*I ��@�I� 4@���V�!?������@�x�"��ٿS�3H ��@���� 4@�G��!?#8q���@��$ц�ٿ���5 ��@�� h 4@g���!?�����@/rbW��ٿNg�3 ��@�!U� 4@q�S��!?wRr���@/rbW��ٿNg�3 ��@�!U� 4@q�S��!?wRr���@P�%6��ٿI��3 ��@���� 4@,�"��!?Y.����@P�%6��ٿI��3 ��@���� 4@,�"��!?Y.����@P�%6��ٿI��3 ��@���� 4@,�"��!?Y.����@P�%6��ٿI��3 ��@���� 4@,�"��!?Y.����@=��R��ٿ�$�- ��@�k�W 4@��mF�!?V�����@=��R��ٿ�$�- ��@�k�W 4@��mF�!?V�����@=��R��ٿ�$�- ��@�k�W 4@��mF�!?V�����@=��R��ٿ�$�- ��@�k�W 4@��mF�!?V�����@��ي�ٿyJ�2 ��@�x$ 4@�m�i��!?�����@�]y��ٿ�L�4 ��@f+�* 4@Ʈ���!?Y����@�]y��ٿ�L�4 ��@f+�* 4@Ʈ���!?Y����@L��Z��ٿv?�5 ��@iSv 4@�0PP��!?�;���@�T�ދ�ٿ/��> ��@�� 4@r:p�!?3*���@%{ػ��ٿ��@ ��@*G�9 4@�WCV��!?�i���@��ʐ��ٿ�)�I ��@�M%� 4@�0��!?.Nٿ��@��ʐ��ٿ�)�I ��@�M%� 4@�0��!?.Nٿ��@��ʐ��ٿ�)�I ��@�M%� 4@�0��!?.Nٿ��@�y���ٿd��J ��@��U� 4@-� >j�!?_y����@��ٿ���E ��@נ� 4@���Zc�!?��;���@��ٿ���E ��@נ� 4@���Zc�!?��;���@��:�ٿ�� C ��@��c� 4@~��\ۏ!?��m���@��z���ٿB�C ��@��B 4@m���L�!?������@��z���ٿB�C ��@��B 4@m���L�!?������@��z���ٿB�C ��@��B 4@m���L�!?������@��z���ٿB�C ��@��B 4@m���L�!?������@��z���ٿB�C ��@��B 4@m���L�!?������@ǲ���ٿ0�D ��@��?� 4@�� 5�!?Z�r��@�9+���ٿK�kF ��@Z��5 4@/=�⤐!?X	�z��@�9+���ٿK�kF ��@Z��5 4@/=�⤐!?X	�z��@�9+���ٿK�kF ��@Z��5 4@/=�⤐!?X	�z��@��dC��ٿ_��H ��@�f 4@ &�ҭ�!?/����@��dC��ٿ_��H ��@�f 4@ &�ҭ�!?/����@�{%��ٿ��F ��@�� 4@��[^�!?;�'���@��l$��ٿ���K ��@�9 4@M�(ؐ!?�T���@� p��ٿ$��F ��@�L�D 4@�����!?�����@�h"�ٿ­�E ��@���� 4@dT^�B�!?�sؖ��@�h"�ٿ­�E ��@���� 4@dT^�B�!?�sؖ��@�h"�ٿ­�E ��@���� 4@dT^�B�!?�sؖ��@ N�w��ٿ"r�H ��@)_�s 4@/Љ^n�!?������@�V���ٿ� H ��@5�ӕ 4@T��|�!?�����@�/�꒙ٿ�$@ ��@Sg� 4@�S*+A�!?!^���@������ٿ�? ��@�<J� 4@�ɢ�]�!?ם��@������ٿM< ��@�` 4@S;QM�!?'�����@������ٿ^��? ��@T�~ 4@5��!?�����@������ٿ^��? ��@T�~ 4@5��!?�����@�m�b��ٿt�A ��@
�� 4@��q�!?!���@�m�b��ٿt�A ��@
�� 4@��q�!?!���@�m�b��ٿt�A ��@
�� 4@��q�!?!���@`�k��ٿ�D ��@:��� 4@-&Q�T�!?i�����@��j��ٿ��wF ��@��n� 4@.��Z�!?l�D���@��j��ٿ��wF ��@��n� 4@.��Z�!?l�D���@��j��ٿ��wF ��@��n� 4@.��Z�!?l�D���@<�.H��ٿ�VI ��@Ƭ�� 4@�S􇇐!?J�]���@�yRl��ٿ�XvG ��@l�`| 4@��S7�!?�H���@!>D3��ٿ�08G ��@o�|� 4@JJ�+�!?������@���W��ٿ��H ��@2,� 4@�]:�!?�]s���@Xߚ�ٿ�*K ��@�,N� 4@?SƳ�!?(o����@Xߚ�ٿ�*K ��@�,N� 4@?SƳ�!?(o����@������ٿ��H ��@:�� 4@nw%��!?#"t���@������ٿ��H ��@:�� 4@nw%��!?#"t���@������ٿ��H ��@:�� 4@nw%��!?#"t���@������ٿ��H ��@:�� 4@nw%��!?#"t���@i�ٔ�ٿ�IN ��@�y
� 4@��%��!?X����@\bߐ�ٿ6~�Q ��@ r�� 4@�KRX�!?I����@�銙ٿ�YP ��@��Em 4@64����!?#pA���@bV�E��ٿ�K]S ��@��B� 4@e!����!?�t����@���ℙٿ��O ��@�d 4@��h��!?�b����@���ℙٿ��O ��@�d 4@��h��!?�b����@�"d��ٿ���K ��@ϲ�� 4@��!.z�!?{�����@�"d��ٿ���K ��@ϲ�� 4@��!.z�!?{�����@�"d��ٿ���K ��@ϲ�� 4@��!.z�!?{�����@/��匙ٿݵ�O ��@�G|� 4@��C9�!?y%���@�Ϭ���ٿE��U ��@gs� 4@����9�!?�ΐ��@��P��ٿE�3Q ��@U� 4@(�q��!?Lm���@:a����ٿ�']Q ��@��^  4@ֺñ?�!?��6���@�
9K��ٿ�U ��@>�� 4@j���Y�!?�S���@��ٿ��VX ��@	(9� 4@윃�W�!?�%����@͉ʆ��ٿ.��W ��@���P 4@�adQ�!?�;���@�q*���ٿg�W ��@�>a 4@f/dA�!?�����@��Q〙ٿKKb ��@y�ȳ 4@h2A��!?�����@��Q〙ٿKKb ��@y�ȳ 4@h2A��!?�����@~�
���ٿ�o_ ��@q9�� 4@�ށg�!?ّ���@I�����ٿ��c ��@�q�� 4@P�Jn�!?p?.���@I�����ٿ��c ��@�q�� 4@P�Jn�!?p?.���@I�����ٿ��c ��@�q�� 4@P�Jn�!?p?.���@I�����ٿ��c ��@�q�� 4@P�Jn�!?p?.���@ �4*��ٿ�Y_ ��@lM� 4@�[z\�!?7ڷ��@ �4*��ٿ�Y_ ��@lM� 4@�[z\�!?7ڷ��@�(��ٿ�7^ ��@�Uj� 4@��5�!?�3���@�(��ٿ�7^ ��@�Uj� 4@��5�!?�3���@�(��ٿ�7^ ��@�Uj� 4@��5�!?�3���@Ȗ`���ٿY�<\ ��@��� 4@�h�W�!?@i����@=�Y푙ٿ��X ��@��� 4@*���S�!?�����@�ː�ٿ��Z ��@Y�_� 4@ 7�/�!?-� ���@F����ٿ��ba ��@�
z  4@�p�G�!?�O����@n�S|��ٿhg ��@"��P 4@�����!?`W;���@�pSٿwU�_ ��@���� 4@vN��=�!?�N���@H�~�ٿ��\ ��@�%�� 4@t�CV�!?y�e��@�"�M��ٿ�}F\ ��@��a� 4@}]B�?�!?o7����@I�
��ٿN[ ��@g�� 4@�� me�!?������@I�
��ٿN[ ��@g�� 4@�� me�!?������@�d����ٿ��7Y ��@��> 4@1q�!?̒k���@`�<՜�ٿ�� [ ��@��I� 4@���\�!?RB����@����ٿ�,` ��@"[�� 4@�s৕�!?�����@`�Ȓ�ٿ�#}Z ��@��� 4@N��Yː!?~8����@'�䔙ٿ�{�Z ��@e�= 4@���!?c�3���@'�䔙ٿ�{�Z ��@e�= 4@���!?c�3���@�ƙ�ٿ���U ��@G� 4@�DN"̐!?�����@�ƙ�ٿ���U ��@G� 4@�DN"̐!?�����@��!��ٿ̈kR ��@�h�� 4@��ɧ�!?M�m���@��!��ٿ̈kR ��@�h�� 4@��ɧ�!?M�m���@��!��ٿ̈kR ��@�h�� 4@��ɧ�!?M�m���@��!��ٿ̈kR ��@�h�� 4@��ɧ�!?M�m���@��!��ٿ̈kR ��@�h�� 4@��ɧ�!?M�m���@�n㙙ٿ�|L ��@̵s� 4@�P��t�!?�����@7o�ț�ٿ��J ��@�'� 4@(�p_�!?{	���@�"�Q��ٿE}�J ��@�� 4@���E�!?��]���@	$��ٿ�vNH ��@�2� 4@�>|�!?Tk�z��@=b�e��ٿ ,A ��@bm�p 4@�"�n�!?�V���@u�ꠙٿ���< ��@� 4@6f��G�!?6bFs��@U�A���ٿ�	D ��@�`� 4@:��R�!?&Ι���@>��u��ٿ�(C ��@=|�� 4@߅2�!?z����@���F��ٿ��/? ��@ǲ�� 4@dL��!?S���@���F��ٿ��/? ��@ǲ�� 4@dL��!?S���@���F��ٿ��/? ��@ǲ�� 4@dL��!?S���@�3���ٿ�i�? ��@�rd� 4@܌��!?�3���@�;Ӣ�ٿ:��K ��@މ0� 4@�K �!?�Z����@ X�p��ٿ��L ��@�'�{ 4@
A�n
�!?pͪ���@�E��ٿI�	\ ��@�Y� 4@�x/\8�!?�7����@�)K���ٿ�1V ��@�Ѕ� 4@��0.�!?�/���@���\��ٿ�r�W ��@u�� 4@����+�!?�V����@�����ٿR
S ��@O>Q 4@zһ��!?�����@�g����ٿ{��J ��@ҙ*� 4@�(��!?�����@��7���ٿJ4I ��@��� 4@[���p�!?Ժ���@%o̹��ٿ���I ��@�2]� 4@��)X��!?�����@�?���ٿ�o|I ��@��4l 4@Y�����!?t�X���@
�
 ��ٿ�I�N ��@�Rlj 4@�p�;�!?�ʧ���@ nSb��ٿ1aV ��@���Y 4@!
�>�!?�d\���@���و�ٿ�9Y ��@�0R� 4@�K�	�!?)���@�fIΊ�ٿP��U ��@;�d� 4@��	�2�!?`����@�fIΊ�ٿP��U ��@;�d� 4@��	�2�!?`����@��1Y��ٿ�D] ��@�U 4@�}��K�!?�e����@[����ٿ[�
e ��@LW� 4@3�g�8�!?!�����@�9��ٿR(Jb ��@tҰ� 4@x#N�!?Jr_���@�ޗ���ٿ
�O ��@֛-m 4@�K9;�!?C!+���@H�(���ٿp��\ ��@:�6/ 4@�|�K�!?M>m���@c�乄�ٿ�<[ ��@�ƣ 4@��U#4�!?�����@��:~�ٿ�D\ ��@6mf 4@�m�T�!?����@��g�o�ٿ�e ��@�/� 4@��^~�!?G����@F�E�d�ٿ`�h ��@0�� 4@�۲�!?�1l��@N)p�c�ٿ �*c ��@��o 4@@��fT�!?��HZ��@&�T1r�ٿ�b�a ��@�.(� 4@�'3�@�!? �����@&�T1r�ٿ�b�a ��@�.(� 4@�'3�@�!? �����@b�v�ٿ���[ ��@��c. 4@�xRo�!?��n��@x\bs�ٿPwR ��@�.� 4@� k}��!?���T��@T{�j{�ٿ�P O ��@H��� 4@_��m�!?��gz��@�t s�ٿ��%S ��@|�i� 4@%ގ�b�!?�27���@��z7��ٿ���G ��@��y 4@-�� v�!?�9����@�:Ԅ�ٿ��3I ��@��?� 4@�f�lG�!?��u���@��#�ٿ���B ��@ft�� 4@0N���!?��Uk��@��r{�ٿ, �= ��@��� 4@���m�!?�lW_��@U��#l�ٿC#E ��@��[  4@w٭�W�!?;h�b��@�.�@l�ٿV��D ��@,X�� 4@��[Ш�!?ă6o��@�>�k�ٿ_t
= ��@���J 4@Y���u�!?mF�d��@�>�k�ٿ_t
= ��@���J 4@Y���u�!?mF�d��@�>�k�ٿ_t
= ��@���J 4@Y���u�!?mF�d��@?�7hn�ٿ�>0 ��@r�d� 4@�=�A~�!?SP7c��@Ƿ%eq�ٿ�6�' ��@HX� 4@(���-�!?�E_��@�S;RN�ٿ6 ��@��o� 4@�Q�T��!?&���@���5Y�ٿ�ݙ$ ��@ׅ'x 4@�i�x�!?s����@�Z�[�ٿ=�J< ��@��� 4@�_�?�!?�qW��@��c�ٿ��E ��@��D. 4@z�'$�!?E��z��@z(��W�ٿKSP: ��@��
� 4@�fDl{�!?�Q�h��@1���B�ٿ�I�) ��@*dL� 4@	���p�!?HQ�1��@1���B�ٿ�I�) ��@*dL� 4@	���p�!?HQ�1��@J�!�+�ٿC3 ��@8&os 4@jn­X�!?��S���@J�!�+�ٿC3 ��@8&os 4@jn­X�!?��S���@V�}�!�ٿ��!1 ��@�bnq 4@�6��A�!?�ȩ���@X���2�ٿKT�B ��@���Q 4@{2u�!?������@�G�z��ٿk7 ��@?�y� 4@�^����!?H�͎��@��{:�ٿ��{9 ��@gtGe 4@m��kU�!?��C��@��{:�ٿ��{9 ��@gtGe 4@m��kU�!?��C��@�'j@�ٿ���K ��@:5� 4@h�*K�!?������@|�w%�ٿ-ϷC ��@���; 4@�Ѯ���!?[Қ���@���ٿk��M ��@>	�� 4@�]�[�!?!�q���@Uݺ��ٿ���U ��@A&rG 4@0��q�!?A����@�N��6�ٿd��v ��@z1� 4@6��OR�!?Hz��@�N���ٿ��[ ��@2�� 4@
Rey��!?�֘��@���I�ٿ�7` ��@��'� 4@bP��y�!?�%q���@�{���ٿs�4n ��@!�s 4@���Rx�!?['����@|�S�ٿ�h ��@�OM 4@?X���!?L�0��@ϛ�`*�ٿ��A| ��@-�\� 4@��H̀�!?`�A���@Zw�꺘ٿ}	�� ��@��	 4@�����!?�I�/��@�[mw{�ٿ��z� ��@�b��	 4@�bT؊�!?����@�[mw{�ٿ��z� ��@�b��	 4@�bT؊�!?����@�A�2F�ٿ{�g� ��@Ώ�
 4@Ud攐!?���a��@�a�v�ٿ|>� ��@p"�S	 4@S�8�a�!?������@�mo�ٿEL� ��@���) 4@���ʎ�!?A�&��@dic� �ٿ���,��@s��� 4@��Oe�!?|�3���@MD�G��ٿ:͝� ��@��]o
 4@=�Ϗ�!?�n�6��@|$?$�ٿhf� ��@
��
 4@��)�F�!?n����@|$?$�ٿhf� ��@
��
 4@��)�F�!?n����@|$?$�ٿhf� ��@
��
 4@��)�F�!?n����@��p�ٿ�	�� ��@���, 4@����@�!?~�U��@���o��ٿ∻� ��@�Z�~
 4@m&J�!?~a&K��@g��E�ٿ|i��@)� 4@ڻ;�7�!?��.���@g��E�ٿ|i��@)� 4@ڻ;�7�!?��.���@�$�<�ٿ�1s� ��@O�� 4@��!�)�!?�s��@�$�<�ٿ�1s� ��@O�� 4@��!�)�!?�s��@���Y7�ٿ�,�� ��@l��g 4@�� ��!?�jbb��@���Y7�ٿ�,�� ��@l��g 4@�� ��!?�jbb��@UV���ٿ�T6� ��@}��� 4@�F�Y�!?bPɭ��@UV���ٿ�T6� ��@}��� 4@�F�Y�!?bPɭ��@e��(=�ٿ��޳ ��@(��
 4@�	iQ �!?P��V��@e��(=�ٿ��޳ ��@(��
 4@�	iQ �!?P��V��@0�z�ٿB�=� ��@J��@ 4@��	E�!?�
���@������ٿ��V ��@�f� 4@�9�{�!?�|܋��@��!�W�ٿ:i�� ��@���w
 4@��_sI�!?�Mgw��@�.�]��ٿN� ��@kZ�� 4@BU�TP�!?��i���@��j�'�ٿ{������@1�X� 4@���B�!?�E8���@�G�vޘٿ,	����@�T\ 4@[�@<�!?`���@�G�vޘٿ,	����@�T\ 4@[�@<�!?`���@g�H=�ٿ�F����@y� 4@4���4�!?
����@���>/�ٿ�M�����@ϼ�� 4@cIzfd�!?�1X���@3u٘ٿ��+ ��@��e=	 4@vJuM�!?m�?���@�|k��ٿ1ʹ: ��@(�~d	 4@5b�H�!??^�t��@lXۍ�ٿf�4� ��@��$� 4@$Aҋe�!?q��m��@lXۍ�ٿf�4� ��@��$� 4@$Aҋe�!?q��m��@��+G�ٿ���� ��@��� 4@1OXqr�!?�����@��+G�ٿ���� ��@��� 4@1OXqr�!?�����@,$jp��ٿV;�� ��@�벙 4@�#��q�!?ڠK���@��͟J�ٿ\
3� ��@I悭 4@��zj��!?]�����@N���ʕٿAD_� ��@l��] 4@zsz�\�!?8���@����2�ٿ�]� ��@�x4 4@c; ��!?���K��@db���ٿ:�KD��@$~"n 4@�k���!?�����@��s<��ٿCZz���@&�L� 4@H���!?4z�a��@��s<��ٿCZz���@&�L� 4@H���!?4z�a��@��s<��ٿCZz���@&�L� 4@H���!?4z�a��@����B�ٿ��%� ��@6�� 4@U�\ �!?�H9��@����B�ٿ��%� ��@6�� 4@U�\ �!?�H9��@���ٿqN:R ��@�g`
 4@$�t�,�!?�����@���ٿqN:R ��@�g`
 4@$�t�,�!?�����@���ٿqN:R ��@�g`
 4@$�t�,�!?�����@����ٿt�� ��@���Z
 4@tE�d�!?�� ���@�/2�y�ٿ�r� ��@a�v" 4@,x��!?��"���@�/2�y�ٿ�r� ��@a�v" 4@,x��!?��"���@�/2�y�ٿ�r� ��@a�v" 4@,x��!?��"���@@� ���ٿ�s>[��@���
 4@�9A�*�!?��:���@@� ���ٿ�s>[��@���
 4@�9A�*�!?��:���@��K҂�ٿ�m ��@���� 4@���݇�!?������@��K҂�ٿ�m ��@���� 4@���݇�!?������@�)��ޗٿ�?~��@�Ę 4@��j'�!?Rx����@�)��ޗٿ�?~��@�Ę 4@��j'�!?Rx����@/����ٿ�����@�+�� 4@�K.�!?�g����@/����ٿ�����@�+�� 4@�K.�!?�g����@O��X�ٿ\#:���@]�6 4@T@"(#�!?�Ф���@�庰�ٿ�
S� ��@ۍz� 4@��q�e�!?K����@�`��ٿ�V$V ��@�� 4@⃋i�!?wPx���@�&��y�ٿ������@�,� 4@�X9�!?J٢e��@�&��y�ٿ������@�,� 4@�X9�!?J٢e��@.l�h>�ٿU��1��@��� 4@@�`3�!?�ޛ���@|Z���ٿ���� ��@ E 4@�,��;�!?��.}��@��32c�ٿ�n�t��@�&0� 4@v�.Gy�!?R�O>��@��32c�ٿ�n�t��@�&0� 4@v�.Gy�!?R�O>��@��32c�ٿ�n�t��@�&0� 4@v�.Gy�!?R�O>��@��32c�ٿ�n�t��@�&0� 4@v�.Gy�!?R�O>��@���ٿ��K'��@��� 4@WP�څ�!?H���@4�';ٿ�C3��@�i/ 4@ew�Ő!?">���@{?Qu[�ٿ3�_���@̷�N 4@��ng�!?���B��@{?Qu[�ٿ3�_���@̷�N 4@��ng�!?���B��@�P���ٿmw���@�y�9 4@��SL��!?�Łs��@�P���ٿmw���@�y�9 4@��SL��!?�Łs��@�P���ٿmw���@�y�9 4@��SL��!?�Łs��@:��'�ٿ΍N���@�B�}��3@*�V�!?�yh.��@,kx,��ٿ��+%���@ƶ���3@�HNN`�!?3&�F��@,kx,��ٿ��+%���@ƶ���3@�HNN`�!?3&�F��@,kx,��ٿ��+%���@ƶ���3@�HNN`�!?3&�F��@��8�M�ٿ��+9 ��@h܋���3@ٔpM��!?�ؐ��@��8�M�ٿ��+9 ��@h܋���3@ٔpM��!?�ؐ��@y��m��ٿ������@��-��3@2�}d�!?5�m ��@y��m��ٿ������@��-��3@2�}d�!?5�m ��@y��m��ٿ������@��-��3@2�}d�!?5�m ��@:�k
ߚٿ��q���@�6����3@�!�+�!?yt#s��@:�k
ߚٿ��q���@�6����3@�!�+�!?yt#s��@:�k
ߚٿ��q���@�6����3@�!�+�!?yt#s��@4�T���ٿ)�G����@�����3@k}��!?��K���@!�;V��ٿev ���@��|���3@�Gأ`�!?������@!�;V��ٿev ���@��|���3@�Gأ`�!?������@��˜�ٿ�N>����@�)�g��3@�N+@��!?ho,�@��6�j�ٿ������@t�mY��3@ǔ]�!?A�����@ݍ֟ٿ?�%"���@��-���3@��_���!?�\�H��@ݍ֟ٿ?�%"���@��-���3@��_���!?�\�H��@�$F?�ٿ�B_���@в���3@�VFC�!?8Cjg��@�$F?�ٿ�B_���@в���3@�VFC�!?8Cjg��@;�D^�ٿ{ʐx���@�����3@����!?��c1��@-S�$��ٿ�P�y��@�b	 4@��E7�!?�_���@-S�$��ٿ�P�y��@�b	 4@��E7�!?�_���@-S�$��ٿ�P�y��@�b	 4@��E7�!?�_���@���>ȡٿ��d���@�T_;��3@[�Yv�!?�
���@�:�T�ٿz��r ��@��~��3@�5S���!?useK��@�:�T�ٿz��r ��@��~��3@�5S���!?useK��@�:�T�ٿz��r ��@��~��3@�5S���!?useK��@���_w�ٿX�� ��@���  4@�6�2��!?۠���@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@����5�ٿ+� ��@N_� 4@2�!x8�!?0����@�y�&B�ٿ<v����@W�  4@b@pk�!?=r����@s~���ٿ��'���@���" 4@��;9�!?��K���@s~���ٿ��'���@���" 4@��;9�!?��K���@��iI�ٿ������@@N����3@��ُ!?�(��@��iI�ٿ������@@N����3@��ُ!?�(��@��iI�ٿ������@@N����3@��ُ!?�(��@��iI�ٿ������@@N����3@��ُ!?�(��@���ٿ��1���@
e���3@ɏ�U�!?�����@���ٿ��1���@
e���3@ɏ�U�!?�����@���ٿ��1���@
e���3@ɏ�U�!?�����@���ٿ��1���@
e���3@ɏ�U�!?�����@���ٿ��1���@
e���3@ɏ�U�!?�����@�_���ٿ)/}����@R�U���3@(u	r�!?����@�_���ٿ)/}����@R�U���3@(u	r�!?����@�_���ٿ)/}����@R�U���3@(u	r�!?����@�_���ٿ)/}����@R�U���3@(u	r�!?����@�_���ٿ)/}����@R�U���3@(u	r�!?����@�狒�ٿ�$�0���@Q����3@+}��!?(����@t�؍z�ٿف����@����3@q���!?2�N0��@kM2�ٟٿ��ie���@VB"��3@�+�5��!?%�Z+��@kM2�ٟٿ��ie���@VB"��3@�+�5��!?%�Z+��@kM2�ٟٿ��ie���@VB"��3@�+�5��!?%�Z+��@kM2�ٟٿ��ie���@VB"��3@�+�5��!?%�Z+��@�b����ٿB}{����@�ѩ��3@�cX5X�!?;z���@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@gL�'V�ٿ�Cy����@�Q���3@�x25�!?���^��@4��ٿ�0"���@�	<��3@eX#)�!?ِR���@4��ٿ�0"���@�	<��3@eX#)�!?ِR���@��f���ٿU�Zf���@�0I��3@��5�!?""����@���O8�ٿ������@	��3@��]�O�!?�9/���@���O8�ٿ������@	��3@��]�O�!?�9/���@���O8�ٿ������@	��3@��]�O�!?�9/���@���O8�ٿ������@	��3@��]�O�!?�9/���@���O8�ٿ������@	��3@��]�O�!?�9/���@���O8�ٿ������@	��3@��]�O�!?�9/���@~�}��ٿC8:���@�Vh0��3@[��[�!?b�IB��@jZ��˟ٿsn����@
�$VR�3@FO�o��!?(�u/��@jZ��˟ٿsn����@
�$VR�3@FO�o��!?(�u/��@jZ��˟ٿsn����@
�$VR�3@FO�o��!?(�u/��@�_��ٿĜ.x��@D �3@���U�!?c8����@��R}�ٿV������@�)e��3@jDQ��!?{%����@��R}�ٿV������@�)e��3@jDQ��!?{%����@N5/_��ٿҿ6܇�@�H���3@o���!?�wY��@N5/_��ٿҿ6܇�@�H���3@o���!?�wY��@N5/_��ٿҿ6܇�@�H���3@o���!?�wY��@N5/_��ٿҿ6܇�@�H���3@o���!?�wY��@24{��ٿ�:"0���@�퓈��3@2�0'�!?������@24{��ٿ�:"0���@�퓈��3@2�0'�!?������@24{��ٿ�:"0���@�퓈��3@2�0'�!?������@����ϟٿ`0����@6�	���3@#s �u�!?�~A	��@�˕��ٿt�Z����@I�No��3@P}s
8�!?�TT��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@X� ��ٿ2����@���4�3@f��i�!?]��g��@�߫ٿl�3��@V����3@V���!?��l��@�߫ٿl�3��@V����3@V���!?��l��@�߫ٿl�3��@V����3@V���!?��l��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@���8��ٿ-�N��@ ��(�3@�c��l�!?�M��@+�3B�ٿ��B?��@3���3@�o7�ސ!?0����@�D0<�ٿ��S���@�$�h��3@o��TÐ!?v�) �@���ٿT�����@�����3@M-�!?�< �@���ٿT�����@�����3@M-�!?�< �@m�ͽ��ٿ���◄�@��X��3@�NNĐ!?���0# �@%�Q|ӟٿ����@�KVܦ�3@C���!?�$����@%�Q|ӟٿ����@�KVܦ�3@C���!?�$����@{1%S�ٿZ�*XP��@m.�t
4@�Vw:�!?Ÿ�}i�@{1%S�ٿZ�*XP��@m.�t
4@�Vw:�!?Ÿ�}i�@կ�(�ٿA�\`��@wk�4@rߩ��!?�kҪ�@կ�(�ٿA�\`��@wk�4@rߩ��!?�kҪ�@<��*�ٿi~�dӉ�@�t'kt4@�t� ~�!?�V0��@M��+�ٿ�Ldm��@C��Qb�3@�(U[�!?s����@M��+�ٿ�Ldm��@C��Qb�3@�(U[�!?s����@M��+�ٿ�Ldm��@C��Qb�3@�(U[�!?s����@M��+�ٿ�Ldm��@C��Qb�3@�(U[�!?s����@M��+�ٿ�Ldm��@C��Qb�3@�(U[�!?s����@A�[���ٿ�dHK��@(G��@�3@�E�;�!?���Z-�@A�[���ٿ�dHK��@(G��@�3@�E�;�!?���Z-�@A�[���ٿ�dHK��@(G��@�3@�E�;�!?���Z-�@A�[���ٿ�dHK��@(G��@�3@�E�;�!?���Z-�@��h�ٿb�X��@$��Ώ�3@�����!?�?G���@��h�ٿb�X��@$��Ώ�3@�����!?�?G���@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@T���ߠٿ-!<�.��@v�.�4@�?�G�!?��u�u�@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@�4~�	�ٿW��lԈ�@�8�4@�jW�n�!?`�vZ��@oD��z�ٿ�ua���@/^Q,�4@d�^h_�!?�4��@oD��z�ٿ�ua���@/^Q,�4@d�^h_�!?�4��@oD��z�ٿ�ua���@/^Q,�4@d�^h_�!?�4��@oD��z�ٿ�ua���@/^Q,�4@d�^h_�!?�4��@ZqoK��ٿ#�0�#��@��v)4@m�mr�!??+�*�@ZqoK��ٿ#�0�#��@��v)4@m�mr�!??+�*�@C��Y.�ٿ�DN�(��@�G�H�3@+!EΆ�!?$�-�@:����ٿ -m�g��@��a��
4@b�;���!?�0���@#�]r�ٿ+��Z@��@Z.p��3@:'͙(�!?�����@#�]r�ٿ+��Z@��@Z.p��3@:'͙(�!?�����@#�]r�ٿ+��Z@��@Z.p��3@:'͙(�!?�����@#�]r�ٿ+��Z@��@Z.p��3@:'͙(�!?�����@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@~��<�ٿ9�^����@�sY'��3@�B"Ȳ�!?���" �@�Op��ٿ�*̹i��@R�Hw�3@8�>��!?�꠬��@�Op��ٿ�*̹i��@R�Hw�3@8�>��!?�꠬��@D��2\�ٿ���sI��@F	�5�3@�<z�!?��J�@��*��ٿS�^ޣ��@iyk�\<4@��EH�!?�dRK��@w֖� �ٿ� �5���@�j�&4@JѹtK�!?=�W"�@ Y�C��ٿ�a����@�vU G4@���]�!?���Rt�@ Y�C��ٿ�a����@�vU G4@���]�!?���Rt�@#�lq�ٿ���W���@�!��4@Hd���!?ɦ��@��b�ٿ��t���@/�(�'4@zNd�!?C��9�	�@��b�ٿ��t���@/�(�'4@zNd�!?C��9�	�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@��u�ٿ)�� ��@8�C84@��2�"�!?sgc[�@f3��+�ٿe��׏�@�߱>4@�����!?�俠��@f3��+�ٿe��׏�@�߱>4@�����!?�俠��@\]��ٿ�ы��@Ep4�/4@� ��:�!?ښ����@\]��ٿ�ы��@Ep4�/4@� ��:�!?ښ����@��ro˜ٿ���N���@h☠�-4@~d]��!?.���u
�@��ro˜ٿ���N���@h☠�-4@~d]��!?.���u
�@?[��єٿ��*��@`خ�4@���>�!?�+��&�@?[��єٿ��*��@`خ�4@���>�!?�+��&�@?[��єٿ��*��@`خ�4@���>�!?�+��&�@?ىٿ����$��@b��h�04@56��!?I8���
�@+�q��ٿk������@�Qwg�4@J�ZI�!?�	%���@+�q��ٿk������@�Qwg�4@J�ZI�!?�	%���@+�q��ٿk������@�Qwg�4@J�ZI�!?�	%���@^P��9�ٿq�뗃�@A50���3@x��Rp�!?�ta%��@^P��9�ٿq�뗃�@A50���3@x��Rp�!?�ta%��@^P��9�ٿq�뗃�@A50���3@x��Rp�!?�ta%��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@\(H�Ҟٿ>�i����@������3@$�h�0�!?g�mn��@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@Z��-l�ٿ�|0<���@>%���3@�<.��!?T�3���@>M]�ٿ��^t��@4ooZ��3@��!?�hav=�@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�O�ʠٿ��et��@�2����3@t<��d�!?EvP����@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@�,_�s�ٿ�h5L���@2�.��3@$�o?�!?�W�x�@����ٿ�:,L{��@���4@� �>�!?��O��@����ٿ�:,L{��@���4@� �>�!?��O��@����ٿ�:,L{��@���4@� �>�!?��O��@����ٿ�:,L{��@���4@� �>�!?��O��@����ٿ�:,L{��@���4@� �>�!?��O��@����ٿ�:,L{��@���4@� �>�!?��O��@�6 �*�ٿ��%̲��@���+4@��v@Z�!?L��)��@�6 �*�ٿ��%̲��@���+4@��v@Z�!?L��)��@�6 �*�ٿ��%̲��@���+4@��v@Z�!?L��)��@�d���ٿ[�����@б� 4@!�t�6�!?#O��@�d���ٿ[�����@б� 4@!�t�6�!?#O��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@g�'�1�ٿT>�
>��@!=.�;�3@��Q�!??�?��@���?��ٿ��<~Ї�@͍ܴ��3@D�G`T�!?9�����@p.IEm�ٿ��TN��@^�5~��3@R�zS�!?�(G��@^��l�ٿ=�@wK��@P%�v�3@ (��i�!?R�����@^��l�ٿ=�@wK��@P%�v�3@ (��i�!?R�����@�]��؟ٿ��f\��@�e��]�3@\�S�H�!?/���}��@�]��؟ٿ��f\��@�e��]�3@\�S�H�!?/���}��@�]��؟ٿ��f\��@�e��]�3@\�S�H�!?/���}��@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@K��|�ٿj4 ��@��p�4@ ]lL:�!?���t%�@�谛΢ٿ�g��&��@�H���
4@��e�!?O9h��@}=�5�ٿ�d����@���Xq	4@!@��ؐ!?J����@}=�5�ٿ�d����@���Xq	4@!@��ؐ!?J����@}=�5�ٿ�d����@���Xq	4@!@��ؐ!?J����@}=�5�ٿ�d����@���Xq	4@!@��ؐ!?J����@\D�Z@�ٿ����#��@'�24@}կ`��!?�i��
�@\D�Z@�ٿ����#��@'�24@}կ`��!?�i��
�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@�|!�]�ٿ/���g��@���<+4@$�RB�!?�s���	�@yv\�\�ٿ>_�K��@	�t��3@�W��6�!?����@yv\�\�ٿ>_�K��@	�t��3@�W��6�!?����@yv\�\�ٿ>_�K��@	�t��3@�W��6�!?����@yv\�\�ٿ>_�K��@	�t��3@�W��6�!?����@�P���ٿ�����@w1�4@w�=�z�!?d���Z�@�A�~�ٿ�'yC��@��7;�4@?��A5�!?���M��@�A�~�ٿ�'yC��@��7;�4@?��A5�!?���M��@�A�~�ٿ�'yC��@��7;�4@?��A5�!?���M��@�A�~�ٿ�'yC��@��7;�4@?��A5�!?���M��@�3Q忠ٿ3�N�#��@&�~��4@�d-�R�!?�KP	�@�3Q忠ٿ3�N�#��@&�~��4@�d-�R�!?�KP	�@�3Q忠ٿ3�N�#��@&�~��4@�d-�R�!?�KP	�@����+�ٿ�u+���@	�.2Y4@8����!?�7@�@u�Ѣ:�ٿ�������@s����94@�F^�!?F�ځ�@�9����ٿt�cgx��@��D4@Ӡ'���!?>7D�@[�(՚ٿu=b���@*v�14@�vL��!? 6_�_
�@[�(՚ٿu=b���@*v�14@�vL��!? 6_�_
�@[�(՚ٿu=b���@*v�14@�vL��!? 6_�_
�@./��:�ٿY)�7��@!����p4@xVM�>�!?�Հ;7�@9�c��ٿc �ms��@��
qgT4@��IpϏ!?�1�{�@9�c��ٿc �ms��@��
qgT4@��IpϏ!?�1�{�@�l21�ٿ�������@�?b^4@'|�j��!?�@v���@:4��ڗٿb�p�T{�@b�G���3@@�5��!?�Tpˎ��@ˎG��ٿm`�e��@�k���3@�W�N��!?���� �@ˎG��ٿm`�e��@�k���3@�W�N��!?���� �@ˎG��ٿm`�e��@�k���3@�W�N��!?���� �@�k4
~�ٿ��kx���@�n����3@O)yؐ!?�{i���@�k4
~�ٿ��kx���@�n����3@O)yؐ!?�{i���@�k4
~�ٿ��kx���@�n����3@O)yؐ!?�{i���@���ud�ٿ��^b��@*G3�34@�S��!??�p��@���ud�ٿ��^b��@*G3�34@�S��!??�p��@���ud�ٿ��^b��@*G3�34@�S��!??�p��@���ud�ٿ��^b��@*G3�34@�S��!??�p��@���ud�ٿ��^b��@*G3�34@�S��!??�p��@���ud�ٿ��^b��@*G3�34@�S��!??�p��@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@�V��B�ٿb�Bu
��@ �P�/\4@�%�C�!?1ad���@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@9V��ٿ`��Ѝ�@��t�24@4����!?@��	�@��Z^��ٿ�}u���@Ph�*4@�_�\�!?LwY�	�@��Z^��ٿ�}u���@Ph�*4@�_�\�!?LwY�	�@��Z^��ٿ�}u���@Ph�*4@�_�\�!?LwY�	�@J��i�ٿ^�\N���@6q��c4@��Be!�!?�"�Q�@J��i�ٿ^�\N���@6q��c4@��Be!�!?�"�Q�@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@�� ?�ٿ�z��|�@�뭧3@�6)Ӽ�!?�t�F���@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@���lݨٿ��4�_��@���w�3@���g�!?c�ut, �@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@�u�.��ٿ�QK��@�N�E�Y4@i���؏!?g����@Iץ���ٿ(�[���@�)��Q4@J^ɗ��!?'����@�����ٿO�����@�!M��44@)�����!?�dMQ�@�����ٿO�����@�!M��44@)�����!?�dMQ�@�����ٿO�����@�!M��44@)�����!?�dMQ�@z�X&��ٿ@Ǯ|т�@��6��3@�c��ؐ!?1�;���@z�X&��ٿ@Ǯ|т�@��6��3@�c��ؐ!?1�;���@z�X&��ٿ@Ǯ|т�@��6��3@�c��ؐ!?1�;���@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@i	@�ٿ��_����@9��J��3@�r:p!�!?��ӭ�@��l�k�ٿ��,()��@��h���3@���x�!?�"m �@��l�k�ٿ��,()��@��h���3@���x�!?�"m �@��l�k�ٿ��,()��@��h���3@���x�!?�"m �@��l�k�ٿ��,()��@��h���3@���x�!?�"m �@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@x�T���ٿ7((�d��@*�Q2��3@��ÄI�!?�?����@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@�WCE�ٿq�?��@p�Ҥ-4@>Z�;H�!?'Fg
�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@��� ^�ٿr_pC���@����Z:4@爴���!?��7k:�@�q%R˚ٿZ��a���@Y�x�0�3@� ~��!?ßˊ�@e��Ϙٿ�7~=ό�@0���&4@�B���!?a�5	�@�Wܹ�ٿ�`W^e��@���4@]]��h�!?����@�Wܹ�ٿ�`W^e��@���4@]]��h�!?����@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@�}�V��ٿ|����@瑬7�4@Z�{�~�!?VP��@ι󡌜ٿ)"	Eۍ�@iT0��)4@��D:�!?��+Y7�@ι󡌜ٿ)"	Eۍ�@iT0��)4@��D:�!?��+Y7�@ι󡌜ٿ)"	Eۍ�@iT0��)4@��D:�!?��+Y7�@���ga�ٿ�S;���@jQ�3�3@����!?������@���ga�ٿ�S;���@jQ�3�3@����!?������@����l�ٿFq}<�|�@��[�3@����̏!?�!W���@����l�ٿFq}<�|�@��[�3@����̏!?�!W���@����l�ٿFq}<�|�@��[�3@����̏!?�!W���@����l�ٿFq}<�|�@��[�3@����̏!?�!W���@yg�ٿa�_����@n@|�3@�H�PΏ!?��S�;��@yg�ٿa�_����@n@|�3@�H�PΏ!?��S�;��@yg�ٿa�_����@n@|�3@�H�PΏ!?��S�;��@��#U>�ٿ�����@�ˬ�5�3@�Ͼ��!?��1���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@+!��8�ٿ�^���@떊���3@�,H��!?'�"���@��go�ٿ��"�3��@kѶ�P�3@d��ka�!?WH�S�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@#��ãٿgq���@"�<��,4@��j��!?��N3
�@�.�p	�ٿ�YHB��@���4@"=�!?��/��@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@o`>���ٿ��Z����@�!؟%4@��X-�!?��[	�@��>^m�ٿ���	 ��@
����3@QC�,�!?�I.[%�@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@l@�j�ٿ�w���@]5����3@����!?n��_��@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@2����ٿ.�����@As`���3@Xx*U�!?{�T�f�@ZSan�ٿ�D�YC��@�L�ip�3@>��Q�!?�;��@���v�ٿ&Na3щ�@���?�3@۝�
�!?����@���v�ٿ&Na3щ�@���?�3@۝�
�!?����@���v�ٿ&Na3щ�@���?�3@۝�
�!?����@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@������ٿ
�;�ʋ�@�GV"t4@|֌\�!?�6 �_�@)����ٿn�F��@}*"s4@�vk�b�!?�/R�@)����ٿn�F��@}*"s4@�vk�b�!?�/R�@)����ٿn�F��@}*"s4@�vk�b�!?�/R�@���O.�ٿX]�.��@��){04@8%��B�!?T��� �@���O.�ٿX]�.��@��){04@8%��B�!?T��� �@���O.�ٿX]�.��@��){04@8%��B�!?T��� �@��� �ٿ���{��@	1(�)4@�����!?ˇ�����@��� �ٿ���{��@	1(�)4@�����!?ˇ�����@��� �ٿ���{��@	1(�)4@�����!?ˇ�����@��� �ٿ���{��@	1(�)4@�����!?ˇ�����@��� �ٿ���{��@	1(�)4@�����!?ˇ�����@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@3b�矠ٿo������@Fw��3@���Om�!?�$�� �@�ќ \�ٿ�\$�4��@��_a
4@��~�h�!?�a7 ��@�ќ \�ٿ�\$�4��@��_a
4@��~�h�!?�a7 ��@�x$<�ٿo�9u��@����+�3@'��N�!?Q߭<m�@�x$<�ٿo�9u��@����+�3@'��N�!?Q߭<m�@�x$<�ٿo�9u��@����+�3@'��N�!?Q߭<m�@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�;�H��ٿ�����@����3@����[�!?5d.��@�{�p��ٿ}Լ���@{�L���3@����:�!?�0q�@�{�p��ٿ}Լ���@{�L���3@����:�!?�0q�@�{�p��ٿ}Լ���@{�L���3@����:�!?�0q�@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@�U��Y�ٿ�9��Z��@��hm%4@j#_�g�!?�����@kb5J�ٿ���e��@z<k��4@����e�!?S��@kb5J�ٿ���e��@z<k��4@����e�!?S��@kb5J�ٿ���e��@z<k��4@����e�!?S��@�l��Q�ٿ�c�c��@V���24@��{�b�!?��F����@�l��Q�ٿ�c�c��@V���24@��{�b�!?��F����@�l��Q�ٿ�c�c��@V���24@��{�b�!?��F����@5vR�ٿ�.u��@��	�w�3@�WY�%�!?���Z���@5vR�ٿ�.u��@��	�w�3@�WY�%�!?���Z���@$��d�ٿ1t�Ҁ�@�U{2�3@p�?P�!?c�x��@$��d�ٿ1t�Ҁ�@�U{2�3@p�?P�!?c�x��@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@�_�3	�ٿ�B�?��@J����3@V���P�!?
����@A\�ۘٿ�qz��@pғ��3@��d�!?���9�@A\�ۘٿ�qz��@pғ��3@��d�!?���9�@���Q��ٿ0���|�@:c%��3@D	�8�!?�@{S�@���Q��ٿ0���|�@:c%��3@D	�8�!?�@{S�@N���ٿ���:�x�@o��N� 4@�X¸��!?�74�B��@N���ٿ���:�x�@o��N� 4@�X¸��!?�74�B��@N���ٿ���:�x�@o��N� 4@�X¸��!?�74�B��@N���ٿ���:�x�@o��N� 4@�X¸��!?�74�B��@J+���ٿr�S�hw�@��R��4@����!?��^�|ږ@J+���ٿr�S�hw�@��R��4@����!?��^�|ږ@J+���ٿr�S�hw�@��R��4@����!?��^�|ږ@J+���ٿr�S�hw�@��R��4@����!?��^�|ږ@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@���z�ٿ�A=����@��Һ04@�����!?�}{���@׆o���ٿkF�]��@�G�s��3@YҼ��!?���	�@0�٪��ٿ��4���@��X��3@�鬦G�!?[��)#�@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@㓎�7�ٿ��d���@�����4@�6�؏!?�:����@p�U{��ٿ�P��pv�@}�_�=C4@�}�\R�!?���`Ζ@p�U{��ٿ�P��pv�@}�_�=C4@�}�\R�!?���`Ζ@p�U{��ٿ�P��pv�@}�_�=C4@�}�\R�!?���`Ζ@p�U{��ٿ�P��pv�@}�_�=C4@�}�\R�!?���`Ζ@�U�![�ٿ���CH��@!��w@>4@@�-MR�!?��Ck��@�U�![�ٿ���CH��@!��w@>4@@�-MR�!?��Ck��@�U�![�ٿ���CH��@!��w@>4@@�-MR�!?��Ck��@��&D;�ٿ�@e��@u9�0�3@N-���!?M'*�=�@��&D;�ٿ�@e��@u9�0�3@N-���!?M'*�=�@Du��W�ٿ���u�@�����3@��  �!?Y����@Du��W�ٿ���u�@�����3@��  �!?Y����@���3O�ٿY<�Oe�@K�����3@��?��!?�x̸��@�3��ٿ���s[�@�ŵ��3@N?�-̏!?�h���@c�����ٿ�&��_b�@kAE�3@�a��!?G��o[��@NI�#��ٿ���rj}�@޸�L�3@����Q�!?g#��F�@̝����ٿ�X,�j��@����3@P�����!?�B�4���@̝����ٿ�X,�j��@����3@P�����!?�B�4���@̝����ٿ�X,�j��@����3@P�����!?�B�4���@�U$5�ٿ��Cn�@gEh�3@fҙ;y�!?-�*�ʖ@�U$5�ٿ��Cn�@gEh�3@fҙ;y�!?-�*�ʖ@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�fS�[�ٿ�&�,Bf�@���C�;4@Q��!?�Ir��@�����ٿ��=��K�@K�צ�K4@�E�Z�!?����r�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@�I߹ޖٿd��9�@�O�@(64@'[J�:�!?&T���I�@?�hs�ٿ�O�@&�h~4@[>u.�!?��"��@?�hs�ٿ�O�@&�h~4@[>u.�!?��"��@?�hs�ٿ�O�@&�h~4@[>u.�!?��"��@�$��6�ٿX��T��@{z����3@����!?����w�@��6�ܦٿ�[����@;�E�E4@�E5�!?�o��˕@�a6�ٿҞ8*���@�}�J�U4@�]�!?��N�g��@�a6�ٿҞ8*���@�}�J�U4@�]�!?��N�g��@�a6�ٿҞ8*���@�}�J�U4@�]�!?��N�g��@�a6�ٿҞ8*���@�}�J�U4@�]�!?��N�g��@|�u��ٿ��n����@��4�Vb4@<�)��!?Bi��R�@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�����ٿk鬒���@ۏ��+4@�%5�!?��A���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@�1�ٿ��8���@�
�/�M4@���!?0�W���@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@>�/��ٿ7��cbq�@���|�3@G�ifI�!?y����ɖ@���JL�ٿ��j�1�@�0�4��3@�8��%�!?p{�*S?�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@爩�m�ٿ3���H�@��mj��3@� 8�!?�n[hDk�@l�O�g�ٿ�O:C��@�cI�3@��٤��!?�˄�ȕ@l�O�g�ٿ�O:C��@�cI�3@��٤��!?�˄�ȕ@l�O�g�ٿ�O:C��@�cI�3@��٤��!?�˄�ȕ@l�O�g�ٿ�O:C��@�cI�3@��٤��!?�˄�ȕ@l�O�g�ٿ�O:C��@�cI�3@��٤��!?�˄�ȕ@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�n�0�ٿI%��<�@��o4@!��i�!?�)nf�Y�@�AP�ٿ��	�2�@�M4�Z4@�-����!?�'Ӹp;�@p���L�ٿ �ƞ,4�@rԜ��14@M+�qj�!?��f�yN�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�(÷Дٿ�)�C�+�@I辉�54@[#��(�!?dW��^;�@�zHw��ٿ��W��7�@P,�N�3@���Ώ!?����M�@�zHw��ٿ��W��7�@P,�N�3@���Ώ!?����M�@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@��c4�ٿ�%*���@i},Z4@�C�C֏!?i<���@�F�GY�ٿ(i�� ��@Z-��&4@[�1��!?n�*Â�@�F�GY�ٿ(i�� ��@Z-��&4@[�1��!?n�*Â�@�F�GY�ٿ(i�� ��@Z-��&4@[�1��!?n�*Â�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@i����ٿ]]�H�f�@J����3@���:B�!?K��Ǯ�@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@�ZK��ٿ�x�����@�'���4@��Ht;�!?�t��Ǖ@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@:�;ޛٿ����@0�)4@�j����!?���an�@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@2%��џٿ@[�!�@?��4@^[)+�!?HF��@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@8sZRЛٿ�>Vw �@"���4@Һ J��!?�0�z� �@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@a�p��ٿR�E��@�ĵ�4@Dt��!?J�Yޡ��@���"֖ٿ������@�n)A4@#LV��!?��c���@���"֖ٿ������@�n)A4@#LV��!?��c���@���"֖ٿ������@�n)A4@#LV��!?��c���@���"֖ٿ������@�n)A4@#LV��!?��c���@���"֖ٿ������@�n)A4@#LV��!?��c���@� {�W�ٿ�Ψ�v��@�ْ#��3@�N��ޏ!?�ݛ0��@� {�W�ٿ�Ψ�v��@�ْ#��3@�N��ޏ!?�ݛ0��@� {�W�ٿ�Ψ�v��@�ْ#��3@�N��ޏ!?�ݛ0��@� {�W�ٿ�Ψ�v��@�ْ#��3@�N��ޏ!?�ݛ0��@��v�v�ٿ:�D�a�@��	<�3@G5}�!?g������@��v�v�ٿ:�D�a�@��	<�3@G5}�!?g������@ �)�F�ٿ��r
	%�@��kb��3@�I��R�!?O��@ �)�F�ٿ��r
	%�@��kb��3@�I��R�!?O��@G"{�:�ٿ��"��@=˼4@�I>㩐!?��z��@G"{�:�ٿ��"��@=˼4@�I>㩐!?��z��@G"{�:�ٿ��"��@=˼4@�I>㩐!?��z��@G"{�:�ٿ��"��@=˼4@�I>㩐!?��z��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@]��Q�ٿ���\���@��)(�4@�4�I�!?�;K�'��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@@�:�ؘٿ�D�2���@/��w<4@X!��-�!?.V�1��@�2����ٿ�#y.��@sՕ\K4@����!?:�u�Ε@�2����ٿ�#y.��@sՕ\K4@����!?:�u�Ε@�2����ٿ�#y.��@sՕ\K4@����!?:�u�Ε@hQtM��ٿlX�n��@����4@�J�&�!?��z�@hQtM��ٿlX�n��@����4@�J�&�!?��z�@hQtM��ٿlX�n��@����4@�J�&�!?��z�@hQtM��ٿlX�n��@����4@�J�&�!?��z�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@�lpi=�ٿ�k�-�@GӢ1&4@�Yڒ6�!?��FsD�@B��ٿ����"�@��z���3@ԝ� ��!?��c$�@B��ٿ����"�@��z���3@ԝ� ��!?��c$�@n~k�ٿ�nJ<��@�-�5�3@��Mp�!?y�E�c�@3���X�ٿkQ=���@��2��3@��r���!?B�Dw(��@3���X�ٿkQ=���@��2��3@��r���!?B�Dw(��@I�}��ٿ��E��!�@�Y�
�3@��\�!?��-���@��>��ٿ���1�?�@W��0�4@��Ȁ��!?+�xn�@��>��ٿ���1�?�@W��0�4@��Ȁ��!?+�xn�@�����ٿO�t��@G���-�3@����!?wZ߽��@�����ٿO�t��@G���-�3@����!?wZ߽��@�����ٿO�t��@G���-�3@����!?wZ߽��@�����ٿO�t��@G���-�3@����!?wZ߽��@��k��ٿMk�L��@p��5�3@��3��!?��5<���@��k��ٿMk�L��@p��5�3@��3��!?��5<���@��k��ٿMk�L��@p��5�3@��3��!?��5<���@��k��ٿMk�L��@p��5�3@��3��!?��5<���@��k��ٿMk�L��@p��5�3@��3��!?��5<���@��k��ٿMk�L��@p��5�3@��3��!?��5<���@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@*��)�ٿl����@1;�ؘ4@��_�.�!?ǫj��@o?'��ٿ�7�@��Eze�3@�򨴑�!?B���
�@o?'��ٿ�7�@��Eze�3@�򨴑�!?B���
�@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@���ٿ�*"U��@t�{��+4@.�x+S�!?��cRV��@��W#��ٿ�nSy�@g4�'4@��2/�!?̺���@��W#��ٿ�nSy�@g4�'4@��2/�!?̺���@�jX��ٿ�8X��@�`�?
4@:k�9Ő!?�Q!�@�jX��ٿ�8X��@�`�?
4@:k�9Ő!?�Q!�@�jX��ٿ�8X��@�`�?
4@:k�9Ő!?�Q!�@�jX��ٿ�8X��@�`�?
4@:k�9Ő!?�Q!�@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@p�φӘٿ�,� S��@*o����3@~H���!?�U�yu��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@yF�B�ٿDp"�#�@�,2�4@f
{e�!?%�n��@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@i`Bg��ٿ#f��s �@��6^.'4@*��d�!?ĮK�Е@�_}�s�ٿ*(8¤�@�����3@���
��!?z�ri��@�n����ٿ��c 	�@��*�i/4@4`.�!?���u|ܕ@�n����ٿ��c 	�@��*�i/4@4`.�!?���u|ܕ@�n����ٿ��c 	�@��*�i/4@4`.�!?���u|ܕ@�n����ٿ��c 	�@��*�i/4@4`.�!?���u|ܕ@�n����ٿ��c 	�@��*�i/4@4`.�!?���u|ܕ@�Bԉ��ٿ��ּ���@S$n�!4@p*�~�!?� �4��@�Bԉ��ٿ��ּ���@S$n�!4@p*�~�!?� �4��@�Bԉ��ٿ��ּ���@S$n�!4@p*�~�!?� �4��@�Bԉ��ٿ��ּ���@S$n�!4@p*�~�!?� �4��@�Bԉ��ٿ��ּ���@S$n�!4@p*�~�!?� �4��@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@�+��S�ٿ܃�ҫ�@q� ��Z4@�:�,o�!?
�EwK�@rX��ٿ��|W
�@aM���I4@d���!?��spՕ@�N`ߡ�ٿ�s��1��@ZY^�J4@�C�Xe�!?�0�*�@�N`ߡ�ٿ�s��1��@ZY^�J4@�C�Xe�!?�0�*�@��0Тٿ#����@�ڭ�Th4@|�£:�!?b��}O�@��0Тٿ#����@�ڭ�Th4@|�£:�!?b��}O�@��0Тٿ#����@�ڭ�Th4@|�£:�!?b��}O�@��0Тٿ#����@�ڭ�Th4@|�£:�!?b��}O�@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@�| ��ٿ��y���@]�n�[4@]�'�!?�t9���@<��W)�ٿX�[��@e}�4�3@�C�(�!?�_�jBR�@
D/-X�ٿ�Z��� �@(�I0�3@ڿ�>V�!?xl`6���@
D/-X�ٿ�Z��� �@(�I0�3@ڿ�>V�!?xl`6���@
D/-X�ٿ�Z��� �@(�I0�3@ڿ�>V�!?xl`6���@
D/-X�ٿ�Z��� �@(�I0�3@ڿ�>V�!?xl`6���@מ���ٿZ4���M�@�s���3@�v+���!?���kFZ�@מ���ٿZ4���M�@�s���3@�v+���!?���kFZ�@����E�ٿƁ7�c[�@/�fy�%4@�W_���!?�� �p�@����E�ٿƁ7�c[�@/�fy�%4@�W_���!?�� �p�@����E�ٿƁ7�c[�@/�fy�%4@�W_���!?�� �p�@H v�ٿ�'��{�@ŷ�|4@E�8i�!?C�;S���@H v�ٿ�'��{�@ŷ�|4@E�8i�!?C�;S���@H v�ٿ�'��{�@ŷ�|4@E�8i�!?C�;S���@i1y�E�ٿS�U�5�@��,�3@Ը�琐!?ӿZ���@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@M����ٿE-����@8�[���3@a��!?��&Y�@�P���ٿ쨌F���@џ��=4@���U#�!?K`8=���@�P���ٿ쨌F���@џ��=4@���U#�!?K`8=���@�4>�ٿ�B���@�����#4@���cU�!?9��R;�@�4>�ٿ�B���@�����#4@���cU�!?9��R;�@�4>�ٿ�B���@�����#4@���cU�!?9��R;�@�68W�ٿN�K��@Y�L��4@��biH�!?϶�Q_�@�68W�ٿN�K��@Y�L��4@��biH�!?϶�Q_�@�68W�ٿN�K��@Y�L��4@��biH�!?϶�Q_�@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�y�ٿ�Jˣ
�@�x�:��3@�U�dQ�!?f�_��ԕ@�ohK�ٿ��&��4�@$�]Y�4@�"�9�!?�}���@�ohK�ٿ��&��4�@$�]Y�4@�"�9�!?�}���@[0����ٿTl2�$�@��U	*4@d4a�K�!?;\^P��@{�f!��ٿ��1�)�@�y��J-4@�
k�!?��'�05�@{�f!��ٿ��1�)�@�y��J-4@�
k�!?��'�05�@{�f!��ٿ��1�)�@�y��J-4@�
k�!?��'�05�@{�f!��ٿ��1�)�@�y��J-4@�
k�!?��'�05�@4�M��ٿ�,�@;?|�K4@꧅���!?k�A��@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@;>�k9�ٿ�������@ %�w�3@�.�rx�!? kz쭕@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@��U��ٿU�o|�@S(��,4@��9Y�!?Bf�����@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@���ٿ"� H���@�\�!4@�e(P�!?t�N�7s�@����f�ٿ&��{ �@#Ꮺ4@��G�6�!?h	�r-��@I�n�ٿ+��YY�@FB2j
4@F�c��!?p-�����@I�n�ٿ+��YY�@FB2j
4@F�c��!?p-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�`7ĝٿQrNOv'�@"�R�{4@h[9|�!?-�����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@�s.��ٿۢu�R�@'עe�	4@��Ɖ��!?��<����@ո��ٿ��sX�@"��ً.4@�0q�!?�ǋd�Е@S�;놛ٿ�%6섾�@������3@},7(��!?���ĕ@S�;놛ٿ�%6섾�@������3@},7(��!?���ĕ@MY�ԧ�ٿ`]M�!��@o����4@8?[@�!?j6�v'�@MY�ԧ�ٿ`]M�!��@o����4@8?[@�!?j6�v'�@MY�ԧ�ٿ`]M�!��@o����4@8?[@�!?j6�v'�@MY�ԧ�ٿ`]M�!��@o����4@8?[@�!?j6�v'�@��:y�ٿ7��C~�@��y�E�3@m�n�!?<�~EK�@��:y�ٿ7��C~�@��y�E�3@m�n�!?<�~EK�@�ئ��ٿ��]~���@�5�3@$� ŏ�!?���=[ŕ@�ئ��ٿ��]~���@�5�3@$� ŏ�!?���=[ŕ@�[�w�ٿ1��&���@Y+Q��3@��\�F�!?��i�@�[�w�ٿ1��&���@Y+Q��3@��\�F�!?��i�@/SИٿ{���!��@i2i?T�3@g��O�!?tJ�Z%��@/SИٿ{���!��@i2i?T�3@g��O�!?tJ�Z%��@qrɔ�ٿ�.� ���@��t�Q4@���[�!?mU�u��@qrɔ�ٿ�.� ���@��t�Q4@���[�!?mU�u��@qrɔ�ٿ�.� ���@��t�Q4@���[�!?mU�u��@qrɔ�ٿ�.� ���@��t�Q4@���[�!?mU�u��@qrɔ�ٿ�.� ���@��t�Q4@���[�!?mU�u��@2����ٿ���,��@�l�c��3@�VLm�!?��u��@�S��9�ٿ
N�����@V¾\�!4@���4<�!?��~�@a�u���ٿy?�s���@j�G��4@�ļ�ː!?q�.�@b�@a�u���ٿy?�s���@j�G��4@�ļ�ː!?q�.�@b�@a�u���ٿy?�s���@j�G��4@�ļ�ː!?q�.�@b�@a�u���ٿy?�s���@j�G��4@�ļ�ː!?q�.�@b�@�� c��ٿ���@):X�3@����ڐ!?�v['0�@�� c��ٿ���@):X�3@����ڐ!?�v['0�@�� c��ٿ���@):X�3@����ڐ!?�v['0�@���@.�ٿ\�O"���@
�Ś4@T��lm�!?��E��@���@.�ٿ\�O"���@
�Ś4@T��lm�!?��E��@߼Oٯ�ٿ��C��@o��2=4@�lu�F�!?��`!x�@�u�0ҕٿH��G)��@O2���k4@�Y�!?qA -w�@� ɪ�ٿe�P���@}ܐZ�D4@ܥՌ��!?��,����@�'�J�ٿ�� ��f�@D�5��#4@�vg���!?��p��7�@�'�J�ٿ�� ��f�@D�5��#4@�vg���!?��p��7�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@���Šٿ"�,�}��@I��vET4@���!?7p�i\�@2M��ޣٿ�هT7��@r���44@�'���!?�g�ϔ�@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�Jѩ�ٿ��5���@�[���3@I,
F��!?�W���@�g,~�ٿ��ԟ(��@?l�/�4@�����!?a��r�a�@�g,~�ٿ��ԟ(��@?l�/�4@�����!?a��r�a�@1E�;�ٿ�x�Y��@����3@����=�!?T�M!0�@1,�$�ٿ~o����@���3@F˃�ܐ!?�K����@1,�$�ٿ~o����@���3@F˃�ܐ!?�K����@1,�$�ٿ~o����@���3@F˃�ܐ!?�K����@1,�$�ٿ~o����@���3@F˃�ܐ!?�K����@9���ٿ+S���W�@��Hb�	4@��)7{�!?)�lXHv�@9���ٿ+S���W�@��Hb�	4@��)7{�!?)�lXHv�@g��C��ٿa���6e�@4��`4@ݹ�!b�!?N���W�@g��C��ٿa���6e�@4��`4@ݹ�!b�!?N���W�@�֍I�ٿV�*��0�@�U'�p�3@�_�!?���];�@�0���ٿ;�1T���@ij���4@���X�!?�	zC�6�@�0���ٿ;�1T���@ij���4@���X�!?�	zC�6�@�0���ٿ;�1T���@ij���4@���X�!?�	zC�6�@XQ�ٿݧ�Z�@� ~,4@��!�!?1��eA�@��}H�ٿ� ���@�8��!�3@��X�v�!?�����@��}H�ٿ� ���@�8��!�3@��X�v�!?�����@��}H�ٿ� ���@�8��!�3@��X�v�!?�����@��}H�ٿ� ���@�8��!�3@��X�v�!?�����@on_W�ٿ��#�if�@�<ȟ(�3@m�r�P�!?k����D�@on_W�ٿ��#�if�@�<ȟ(�3@m�r�P�!?k����D�@on_W�ٿ��#�if�@�<ȟ(�3@m�r�P�!?k����D�@on_W�ٿ��#�if�@�<ȟ(�3@m�r�P�!?k����D�@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@'L���ٿG9+=��@3�~��4@*�D�!?k��>��@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@u��-רٿ�2c�2�@�k��3@=Ig=K�!?��1�-ʕ@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@��pt8�ٿ����e8�@$	ڠ��3@��p���!?�FV���@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@d9�>#�ٿ#4T���@���˼4@�+�NL�!?N!��k�@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@!����ٿV��⿽�@T��E�4@��^t��!?�A�7>��@���;8�ٿ�A?	�~�@Y�!���3@$t�g�!?�=��9�@����a�ٿ�<yZ�~�@�2�Im�3@���t�!?�KZ��@����a�ٿ�<yZ�~�@�2�Im�3@���t�!?�KZ��@����a�ٿ�<yZ�~�@�2�Im�3@���t�!?�KZ��@4�x~�ٿce����@Z=x��3@h7�vg�!?���e�@4�x~�ٿce����@Z=x��3@h7�vg�!?���e�@4�x~�ٿce����@Z=x��3@h7�vg�!?���e�@4�x~�ٿce����@Z=x��3@h7�vg�!?���e�@56�ٿ
��"��@�ʊ4@8�KRF�!?3o�Jg�@56�ٿ
��"��@�ʊ4@8�KRF�!?3o�Jg�@56�ٿ
��"��@�ʊ4@8�KRF�!?3o�Jg�@56�ٿ
��"��@�ʊ4@8�KRF�!?3o�Jg�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@D�w���ٿ���P���@�Z[E�(4@�ur�!?FL��s�@���a��ٿ&�Z1-$�@��yҏ4@��z�!?�����@���a��ٿ&�Z1-$�@��yҏ4@��z�!?�����@���a��ٿ&�Z1-$�@��yҏ4@��z�!?�����@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@��:�ٿ�CybW@�@�xc
�)4@{��$g�!?�F�cxX�@e���ٿ|��D�x�@aIԚP4@��dx�!?�~�6��@e���ٿ|��D�x�@aIԚP4@��dx�!?�~�6��@e���ٿ|��D�x�@aIԚP4@��dx�!?�~�6��@e���ٿ|��D�x�@aIԚP4@��dx�!?�~�6��@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@	 G;��ٿ�B�U�@H�m�4@�����!? ��͖@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@�c;,5�ٿƨ�����@)��wC 4@]�Z�!?.K1\ɕ@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@T���ٿ�Ԭg�@AL=f4@J���l�!?ݎ� �@q��oٝٿt��=�@~��ޭJ4@���Gs�!?�)�2�u�@q��oٝٿt��=�@~��ޭJ4@���Gs�!?�)�2�u�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@���Lݟٿ;�!���@�`JlH4@$�{Oa�!?Q{L��3�@56��ٿ����?�@W2	=4@6�1�^�!?!%2�ZՖ@56��ٿ����?�@W2	=4@6�1�^�!?!%2�ZՖ@$Y�v�ٿ'���zj�@�bi�4@��B�a�!?ϫ�^�@$Y�v�ٿ'���zj�@�bi�4@��B�a�!?ϫ�^�@$Y�v�ٿ'���zj�@�bi�4@��B�a�!?ϫ�^�@$Y�v�ٿ'���zj�@�bi�4@��B�a�!?ϫ�^�@$Y�v�ٿ'���zj�@�bi�4@��B�a�!?ϫ�^�@�f���ٿ����W��@�S&V84@Ӷ�T�!?��=fŕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@���袗ٿ�)����@���4@R�]]`�!?
T0ӨǕ@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@�z6�ٿ�i�;�@�k>��4@��w�a�!?#{s_�
�@��	�ٿ��E��@.�s{�4@�h �b�!?��R莖@��	�ٿ��E��@.�s{�4@�h �b�!?��R莖@��	�ٿ��E��@.�s{�4@�h �b�!?��R莖@7�����ٿ�����@Epq�(4@�����!?��\�&�@7�����ٿ�����@Epq�(4@�����!?��\�&�@7�����ٿ�����@Epq�(4@�����!?��\�&�@�dҢ�ٿ2�t3R��@h�mM�3@�$�Z:�!?�X��ˢ�@�dҢ�ٿ2�t3R��@h�mM�3@�$�Z:�!?�X��ˢ�@�dҢ�ٿ2�t3R��@h�mM�3@�$�Z:�!?�X��ˢ�@�dҢ�ٿ2�t3R��@h�mM�3@�$�Z:�!?�X��ˢ�@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@�(�=�ٿ��@�]��@>,w�4@۳U�8�!?���F��@%���ٿ�%�AvT�@u� 4@�cĶ��!?��9�]�@��ƈ�ٿ#G�Ij�@/���4@\37Ð!?K�A��@��ƈ�ٿ#G�Ij�@/���4@\37Ð!?K�A��@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@�dj���ٿ��F���@�ފ�4@�b_l�!?Ͱa7�@��͛�ٿ*p`90��@����i�3@[��N�!?;!�7��@��͛�ٿ*p`90��@����i�3@[��N�!?;!�7��@��͛�ٿ*p`90��@����i�3@[��N�!?;!�7��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@k���k�ٿ��A��@�O�� �3@3+\A��!?y��e$��@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@{Um���ٿ�HֶvT�@����94@��!m�!?���[6�@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@�	�u�ٿ�����@�'�#.�3@9�k�o�!?6S��ޕ@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���'ϡٿ�v�U���@����4@��5��!?��:��@���yx�ٿǭ��@�o#�a4@��;H�!?.G��U4�@���yx�ٿǭ��@�o#�a4@��;H�!?.G��U4�@���yx�ٿǭ��@�o#�a4@��;H�!?.G��U4�@���yx�ٿǭ��@�o#�a4@��;H�!?.G��U4�@��A�բٿn�t�G�@l�G�24@�{���!?
CO	��@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@���H�ٿ�@xl�l�@	�N!�*4@�#���!?7���@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@�a�H_�ٿ���&+��@���]g84@g\au�!?�Y���o�@9�!�ѠٿVW���@�S W&4@ P�]��!?����b�@9�!�ѠٿVW���@�S W&4@ P�]��!?����b�@9�!�ѠٿVW���@�S W&4@ P�]��!?����b�@�#\|��ٿ��o��@�!�
4@OM�?��!?�Iuʕ@�#\|��ٿ��o��@�!�
4@OM�?��!?�Iuʕ@�#\|��ٿ��o��@�!�
4@OM�?��!?�Iuʕ@�tSPe�ٿBu���@�j[���3@KSD���!?�:lM��@�tSPe�ٿBu���@�j[���3@KSD���!?�:lM��@�tSPe�ٿBu���@�j[���3@KSD���!?�:lM��@�tSPe�ٿBu���@�j[���3@KSD���!?�:lM��@� ��Śٿ�����/�@;��/�3@�@���!?םĪ(ӕ@� ��Śٿ�����/�@;��/�3@�@���!?םĪ(ӕ@� ��Śٿ�����/�@;��/�3@�@���!?םĪ(ӕ@i WWn�ٿ0��� ��@[��U�3@mqQ�g�!?cρ��ԕ@i WWn�ٿ0��� ��@[��U�3@mqQ�g�!?cρ��ԕ@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@� ����ٿk��"~��@� H��3@~ܡ��!?�}G�B2�@�p�Up�ٿr��:e��@6�]`�4@��¬��!?�>L��"�@�p�Up�ٿr��:e��@6�]`�4@��¬��!?�>L��"�@�p�Up�ٿr��:e��@6�]`�4@��¬��!?�>L��"�@�p�Up�ٿr��:e��@6�]`�4@��¬��!?�>L��"�@�p�Up�ٿr��:e��@6�]`�4@��¬��!?�>L��"�@��ߣٿ��6*�%�@
����3@��%��!?o9�]^�@��ߣٿ��6*�%�@
����3@��%��!?o9�]^�@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@o�
��ٿ�t,!��@�R���3@h6e�>�!?�N7��@�� �ߣٿ�.35��@�0��"4@Snt3��!?�����@�� �ߣٿ�.35��@�0��"4@Snt3��!?�����@�$k��ٿ�׊!
��@~���3@���g�!?~�8.ѕ@0�/�ٿ'r�$W�@�̹�4@�{����!?<�y�@0�/�ٿ'r�$W�@�̹�4@�{����!?<�y�@0�/�ٿ'r�$W�@�̹�4@�{����!?<�y�@0�/�ٿ'r�$W�@�̹�4@�{����!?<�y�@>�,-�ٿI�QH��@@�"�3@��e�!?�Bvy�@>�,-�ٿI�QH��@@�"�3@��e�!?�Bvy�@>�,-�ٿI�QH��@@�"�3@��e�!?�Bvy�@>�,-�ٿI�QH��@@�"�3@��e�!?�Bvy�@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��q*�ٿ\��Hm�@�ȍ#D�3@���&�!?�C�e�Ε@��|M�ٿ�D�/O�@QF�Pf/4@�7�
�!?�ʾ�|��@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@=Kݪ�ٿ�E��&�@��F�W4@��֓��!?ۇ�O���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�<��ٿ�*��U��@ ��?,4@?�����!?���`���@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@�!}�Ϙٿ3f�W���@��P��?4@�B3�n�!?Q=ꩽx�@c0�f̠ٿ���j�@�Q�gL$4@BR;n�!?6��¹�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@���=�ٿ�h�����@/�s��3@��{H�!?u��j�@��A��ٿ��[�< �@�=���3@I9τ&�!?��2��@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@�j�JǛٿ6����@�8z�4@��:�!?�{�s8�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@?�cΚٿ9�|K�W�@�^���?4@l8`��!?�W��G�@r׬�ٿϒ�k%
�@ ��`4@�>B�!?��R���@r׬�ٿϒ�k%
�@ ��`4@�>B�!?��R���@��tY@�ٿ_��r�@��2[�V4@F2�!?��{��@��tY@�ٿ_��r�@��2[�V4@F2�!?��{��@��tY@�ٿ_��r�@��2[�V4@F2�!?��{��@���"�ٿ."9=L>�@E?�WnQ4@D�P-��!?��[���@���"�ٿ."9=L>�@E?�WnQ4@D�P-��!?��[���@���Y��ٿ��Q���@�"��4@u�%�z�!?�3U5�6�@���Y��ٿ��Q���@�"��4@u�%�z�!?�3U5�6�@���Y��ٿ��Q���@�"��4@u�%�z�!?�3U5�6�@d�%_j�ٿ���9X��@���I4@Y"�䶐!?0{Z�k�@d�%_j�ٿ���9X��@���I4@Y"�䶐!?0{Z�k�@o�P�ٿ?����R�@�{~nX4@������!?��{~��@�iُV�ٿ��Za��@M~�QY4@G�}Gb�!?i_����@�iُV�ٿ��Za��@M~�QY4@G�}Gb�!?i_����@�iُV�ٿ��Za��@M~�QY4@G�}Gb�!?i_����@�iُV�ٿ��Za��@M~�QY4@G�}Gb�!?i_����@�iُV�ٿ��Za��@M~�QY4@G�}Gb�!?i_����@�5��N�ٿ�F-Et��@���4@���5��!?�q�pw��@G;�)B�ٿ�b��@V��$4@e4)w�!?���|)P�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@P��o�ٿ�R�����@���4@Bھ3��!?wB �_!�@ip�B�ٿp�k�Q�@ �3T�3@!�����!?��O�	�@��S���ٿ@�} k��@���=��3@�gC�!?��u�~Օ@��S���ٿ@�} k��@���=��3@�gC�!?��u�~Օ@���*��ٿ�6�j��@@G-X��3@���Z��!?�@hzՕ@������ٿ�	�B0��@LL$�'4@��9��!?�;�9�@������ٿ�	�B0��@LL$�'4@��9��!?�;�9�@������ٿ�	�B0��@LL$�'4@��9��!?�;�9�@������ٿ�	�B0��@LL$�'4@��9��!?�;�9�@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@y����ٿ����@�����4@�����!?�����@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@�Se�ٿ���%Q��@�r�p�4@0#q��!?�L���@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@c�򚈘ٿ%fpܴ�@in�ʎ�3@�AeJ�!?�n�z��@���<b�ٿND�c��@[q��b 4@!�<�!?i�d��@���<b�ٿND�c��@[q��b 4@!�<�!?i�d��@���<b�ٿND�c��@[q��b 4@!�<�!?i�d��@���<b�ٿND�c��@[q��b 4@!�<�!?i�d��@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@Jt`�ٿ���-��@�W�2�4@�>��!?�x��~�@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�;���ٿnnҲ��@	���3@eΩk$�!?�Eh����@�)(Nr�ٿPkA���@�
�;4@�;(�|�!?���I �@�)(Nr�ٿPkA���@�
�;4@�;(�|�!?���I �@����P�ٿ��Dg*�@�ġ��?4@����C�!?w0n��@����P�ٿ��Dg*�@�ġ��?4@����C�!?w0n��@����P�ٿ��Dg*�@�ġ��?4@����C�!?w0n��@լD*�ٿ�o �u�@e	�O�4@�XTa,�!?B{��&&�@��~���ٿ�]����@ӌ����3@cx_�e�!?9�m��@��~���ٿ�]����@ӌ����3@cx_�e�!?9�m��@��~���ٿ�]����@ӌ����3@cx_�e�!?9�m��@^1$ؖٿF;�aB�@r����4@�!�!?�G�6��@^1$ؖٿF;�aB�@r����4@�!�!?�G�6��@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@��&Y�ٿ������@�dۈ��3@�<j�!?W�1�E�@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@���ٿ��j�@�t�լ4@���@�!?75�;��@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@n�h�f�ٿ!�x�b��@�O�&�
4@~��t�!?�rEB�ە@y�HC�ٿ>�,	5��@��Md;4@�>R�!?J���Օ@y�HC�ٿ>�,	5��@��Md;4@�>R�!?J���Օ@y�HC�ٿ>�,	5��@��Md;4@�>R�!?J���Օ@�4~羽ٿ��4���@`؋x�/4@���� �!?�)�#�
�@&�n�7�ٿ�T���|�@Gß|�%4@�B#��!?dؖtG��@&�n�7�ٿ�T���|�@Gß|�%4@�B#��!?dؖtG��@�;6��ٿ�`��0�@a*{}�4@I�qBo�!?\�"ѕ@�K�ۣٿ0�d����@�$��4@�#F[�!?� a��Օ@oo�hݠٿ�ק ��@Z!�W4@Nzm���!?b�$����@oo�hݠٿ�ק ��@Z!�W4@Nzm���!?b�$����@����R�ٿv~^ϭ�@91se0�3@#�C��!?`�����@����R�ٿv~^ϭ�@91se0�3@#�C��!?`�����@����R�ٿv~^ϭ�@91se0�3@#�C��!?`�����@����R�ٿv~^ϭ�@91se0�3@#�C��!?`�����@wd��ǝٿ�<�Z��@g��3<4@�Ln踐!?�}.3z֕@wd��ǝٿ�<�Z��@g��3<4@�Ln踐!?�}.3z֕@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@b(�`�ٿ�ι��@�p���3@�չX̐!?M!��2/�@��Rk��ٿ���d�@���4@�`N�!?���R��@��Rk��ٿ���d�@���4@�`N�!?���R��@��Rk��ٿ���d�@���4@�`N�!?���R��@��Rk��ٿ���d�@���4@�`N�!?���R��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@="�x	�ٿ�t���@�2�R'4@O����!?��s��@�7�R��ٿԖz�4O�@���ҍM4@��B��!?7�J<���@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��~�ٿ��` �@�����54@&g`��!?m�KV �@��7�ٿ|L���@����e4@�g>�Đ!?Z)��ޕ@��7�ٿ|L���@����e4@�g>�Đ!?Z)��ޕ@��7�ٿ|L���@����e4@�g>�Đ!?Z)��ޕ@x�:��ٿ���2�@�c� `4@������!?l(�9�@x�:��ٿ���2�@�c� `4@������!?l(�9�@�>G�ٿ\�yK�@>�ٿ4@R���!?��R��@�>G�ٿ\�yK�@>�ٿ4@R���!?��R��@��S!�ٿvW"?�@�\�4@FL���!?6m��ƕ@��S!�ٿvW"?�@�\�4@FL���!?6m��ƕ@��S!�ٿvW"?�@�\�4@FL���!?6m��ƕ@��S!�ٿvW"?�@�\�4@FL���!?6m��ƕ@��S!�ٿvW"?�@�\�4@FL���!?6m��ƕ@�6H�ٿ���ۑM�@[竢�4@v���!?����aQ�@�P}�ٿg�ν���@�?�m�4@(��,��!?��?�VO�@�P}�ٿg�ν���@�?�m�4@(��,��!?��?�VO�@\�r�	�ٿ/e�=��@���G?4@�?���!?t�}���@\�r�	�ٿ/e�=��@���G?4@�?���!?t�}���@ՠ�u��ٿ~�M�a�@3;7��O4@��\,�!?A�����@ՠ�u��ٿ~�M�a�@3;7��O4@��\,�!?A�����@ՠ�u��ٿ~�M�a�@3;7��O4@��\,�!?A�����@ՠ�u��ٿ~�M�a�@3;7��O4@��\,�!?A�����@ՠ�u��ٿ~�M�a�@3;7��O4@��\,�!?A�����@S-�	}�ٿ`���
�@�V�V4@SSUIz�!? `����@��]Iɛٿ��)B��@;-]x/4@sj=	?�!?XYY�Ǖ@��]Iɛٿ��)B��@;-]x/4@sj=	?�!?XYY�Ǖ@��]Iɛٿ��)B��@;-]x/4@sj=	?�!?XYY�Ǖ@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@
�Z{��ٿ�ٟ�J�@c�w?�4@��]}�!?�`�H��@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�u�ٿԄ���@��r�3@��0�=�!?��=)�?�@�f��ٿ����@�#~.4@��84�!?�!s��@�f��ٿ����@�#~.4@��84�!?�!s��@�f��ٿ����@�#~.4@��84�!?�!s��@L��-�ٿ�[�!���@��4@�4*�!?�*PLĕ@t�5=&�ٿ������@�@��K4@ ��M�!?D5cI���@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@��� �ٿB���
 �@@5�+34@��'���!?�_�xb �@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@Am��T�ٿ��>�k��@�8[�4@ҒyC�!?�TY�Ż�@�Mhꮙٿ_ �!�>�@�1B�/4@�0,ߤ�!?m���1�@�Mhꮙٿ_ �!�>�@�1B�/4@�0,ߤ�!?m���1�@�>�
�ٿ�E}x���@�N�54@�{�ܥ�!?���@��^XٚٿV��&���@=�N�14@�!�j�!?��p���@)�샠ٿN�P���@�tM��;4@��r��!?rgP$���@)�샠ٿN�P���@�tM��;4@��r��!?rgP$���@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@�L�ٿ��%b(�@��t�F)4@��|@�!?%�բ�@a/����ٿ�A��A��@d(��#4@��c�!?4-�N�e�@a/����ٿ�A��A��@d(��#4@��c�!?4-�N�e�@a/����ٿ�A��A��@d(��#4@��c�!?4-�N�e�@��2�ٿ�r�T=�@�k��3@���\�!?XX�eЁ�@��2�ٿ�r�T=�@�k��3@���\�!?XX�eЁ�@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@&����ٿr&5��.�@꠬5d4@��'�!?��ԔA��@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@�=ߙٿ�4��@��@G34@�p�L�!?���S=̕@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@a�C��ٿG����@�~ĮE;4@>�*M��!?�����@�2��ٿ9�~��R�@�+��X94@/�S���!?❷aX�@�2��ٿ9�~��R�@�+��X94@/�S���!?❷aX�@�2��ٿ9�~��R�@�+��X94@/�S���!?❷aX�@�2��ٿ9�~��R�@�+��X94@/�S���!?❷aX�@��F0�ٿk9B���@/��%t84@� 	���!?ڰ�Nq��@��F0�ٿk9B���@/��%t84@� 	���!?ڰ�Nq��@��F0�ٿk9B���@/��%t84@� 	���!?ڰ�Nq��@��F0�ٿk9B���@/��%t84@� 	���!?ڰ�Nq��@��F0�ٿk9B���@/��%t84@� 	���!?ڰ�Nq��@hO��B�ٿa���ͭ�@f)�R04@�7��!?��f�j��@hO��B�ٿa���ͭ�@f)�R04@�7��!?��f�j��@hO��B�ٿa���ͭ�@f)�R04@�7��!?��f�j��@hO��B�ٿa���ͭ�@f)�R04@�7��!?��f�j��@�-Mϝٿ �<�f�@r�*��3@s��y�!?T���w�@�-Mϝٿ �<�f�@r�*��3@s��y�!?T���w�@�-Mϝٿ �<�f�@r�*��3@s��y�!?T���w�@9\���ٿ� ��~�@�1YM�>4@�K�v�!?�j���@9\���ٿ� ��~�@�1YM�>4@�K�v�!?�j���@9\���ٿ� ��~�@�1YM�>4@�K�v�!?�j���@9\���ٿ� ��~�@�1YM�>4@�K�v�!?�j���@9\���ٿ� ��~�@�1YM�>4@�K�v�!?�j���@�>0qY�ٿc�ԩ�M�@a�OKf�3@��6�l�!?)�

��@�>0qY�ٿc�ԩ�M�@a�OKf�3@��6�l�!?)�

��@�>0qY�ٿc�ԩ�M�@a�OKf�3@��6�l�!?)�

��@�>0qY�ٿc�ԩ�M�@a�OKf�3@��6�l�!?)�

��@�>0qY�ٿc�ԩ�M�@a�OKf�3@��6�l�!?)�

��@�^S���ٿz`W{z�@��e�3@Zj}:>�!?�.���
�@�^S���ٿz`W{z�@��e�3@Zj}:>�!?�.���
�@�^S���ٿz`W{z�@��e�3@Zj}:>�!?�.���
�@�^S���ٿz`W{z�@��e�3@Zj}:>�!?�.���
�@�E+��ٿ�+�|�@.�g'^4@�{cN�!?� �'�@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@���-�ٿ�D����@r|n�
4@.��;��!?'��ޕ@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@��&Üٿ��R��@��C'4@�Y�(s�!?C�
�j��@�}㽚ٿ�fU���@�'�z�4@0]"��!?�i��Jɕ@�}㽚ٿ�fU���@�'�z�4@0]"��!?�i��Jɕ@�}㽚ٿ�fU���@�'�z�4@0]"��!?�i��Jɕ@�}㽚ٿ�fU���@�'�z�4@0]"��!?�i��Jɕ@�}㽚ٿ�fU���@�'�z�4@0]"��!?�i��Jɕ@��x�ٿ�����@մ��+4@���:��!?��:��@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@_��K_�ٿ���T�@��?x4@S6O�!?��[h�@w�H��ٿ�UE+G��@PVDa4@�P���!?cz|/��@w�H��ٿ�UE+G��@PVDa4@�P���!?cz|/��@w�H��ٿ�UE+G��@PVDa4@�P���!?cz|/��@w�H��ٿ�UE+G��@PVDa4@�P���!?cz|/��@w�H��ٿ�UE+G��@PVDa4@�P���!?cz|/��@�`�3�ٿ�	�/��@�!��84@����'�!?�7�oȝ�@�`�3�ٿ�	�/��@�!��84@����'�!?�7�oȝ�@�`�3�ٿ�	�/��@�!��84@����'�!?�7�oȝ�@N)���ٿSD��e�@u[��4@�Ÿ.=�!?����@�7P}��ٿT,v�|��@�V`��4@nb�!?�]���@*��IL�ٿ��feN��@���f]4@�Dv���!?ޕ�4<��@*��IL�ٿ��feN��@���f]4@�Dv���!?ޕ�4<��@C*���ٿ�b:���@�-���34@���C�!?;�*�,�@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�:U�ٿ�����@�<�@K4@D��;͐!?�~�Y|��@�����ٿ"u�|��@��xxD4@��!r�!?�@�vO�@�����ٿ"u�|��@��xxD4@��!r�!?�@�vO�@t=k(�ٿ�=�h̃�@�5^N94@%n{�O�!?Ў(b�@t=k(�ٿ�=�h̃�@�5^N94@%n{�O�!?Ў(b�@t=k(�ٿ�=�h̃�@�5^N94@%n{�O�!?Ў(b�@t=k(�ٿ�=�h̃�@�5^N94@%n{�O�!?Ў(b�@t=k(�ٿ�=�h̃�@�5^N94@%n{�O�!?Ў(b�@?�&QJ�ٿ�P����@�F��p%4@��D�!?��n麣�@?�&QJ�ٿ�P����@�F��p%4@��D�!?��n麣�@?�&QJ�ٿ�P����@�F��p%4@��D�!?��n麣�@�@��آٿ���~��@��K��4@
�o�!?c?eە@&�,H��ٿ89�a��@�^,]�4@�ѿf��!?۔h�o��@��lO�ٿ��ĥ��@ �V�4@�[�.�!?>۶�p��@��lO�ٿ��ĥ��@ �V�4@�[�.�!?>۶�p��@��lO�ٿ��ĥ��@ �V�4@�[�.�!?>۶�p��@��lO�ٿ��ĥ��@ �V�4@�[�.�!?>۶�p��@#Li� �ٿ�v��g��@�yB��	4@��P;D�!?��rz��@�VD�X�ٿP����#�@T�GP�3@�J�@�!?����_ޕ@�VD�X�ٿP����#�@T�GP�3@�J�@�!?����_ޕ@�VD�X�ٿP����#�@T�GP�3@�J�@�!?����_ޕ@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@�Ĝ�i�ٿا�2;�@��4@��ƿq�!?���߯֕@5]�!�ٿl.�&��@�n� 4@S�s��!?+Kf�^�@5]�!�ٿl.�&��@�n� 4@S�s��!?+Kf�^�@5]�!�ٿl.�&��@�n� 4@S�s��!?+Kf�^�@Z���ٿ.�r?ha�@��l4@�h/5R�!?��}%��@�)�ٿ��;���@0s34@�\�2�!?��8\�ѕ@�)�ٿ��;���@0s34@�\�2�!?��8\�ѕ@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@ONV��ٿ�(�QV��@�W�D4@J����!?�7�w��@�o�ݞٿ��j�8��@4h��%"4@u��p�!?�ֈv/֕@�o�ݞٿ��j�8��@4h��%"4@u��p�!?�ֈv/֕@�o�ݞٿ��j�8��@4h��%"4@u��p�!?�ֈv/֕@�o�ݞٿ��j�8��@4h��%"4@u��p�!?�ֈv/֕@G%j*�ٿۿ��o]�@�D�Nj.4@%V�j{�!?�0]o��@��P���ٿ�Q����@�x}G4@�R�y�!?R>~��@�+�X�ٿ�_�> �@�"�04@�:,��!?�/���@5X�<k�ٿ�S���*�@j�]�4@neϐ!?�h���_�@5X�<k�ٿ�S���*�@j�]�4@neϐ!?�h���_�@�_ꗡٿ���rl��@��|�4@�n�]��!?/��~�@�����ٿ2��@��@9���;4@D��l�!?Z$�+ڕ@~%�d�ٿ9��J��@*n�XE4@1���[�!?$���@ѕ@U�&��ٿ{��X��@�^6�4@�CB"O�!?�3���2�@���q�ٿ�	>V-�@�%-`4@E}���!?h��`
�@���q�ٿ�	>V-�@�%-`4@E}���!?h��`
�@���q�ٿ�	>V-�@�%-`4@E}���!?h��`
�@
�ҚٿK,����@)���f84@\7]�!?�^�Z�@�kMt֛ٿߔn���@�Z���F4@X(W���!?g^�u�@�kMt֛ٿߔn���@�Z���F4@X(W���!?g^�u�@��a$|�ٿf�jG��@���<4@�CF���!?�7 %�@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@!�T�a�ٿK�8M�R�@Tg�4@�@�8�!?E��a��@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@g}�͝ٿ�X
��@N���z4@���!?�
�i
@�@BD�BA�ٿ� �8���@�����4@�}V��!?�BőWE�@BD�BA�ٿ� �8���@�����4@�}V��!?�BőWE�@BD�BA�ٿ� �8���@�����4@�}V��!?�BőWE�@BD�BA�ٿ� �8���@�����4@�}V��!?�BőWE�@u_O{��ٿ�f����@����3@�WU�!?��.��@u_O{��ٿ�f����@����3@�WU�!?��.��@�}볘�ٿ��苉�@��[Q 4@S� �~�!?PU1�Ew�@R��R�ٿ�����@t`)�3@i�2e�!?�I����@R��R�ٿ�����@t`)�3@i�2e�!?�I����@R��R�ٿ�����@t`)�3@i�2e�!?�I����@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@s�'��ٿ���9�@㚽�@4@F��}�!?� *�@�Б7��ٿ}�La�@!i$~��3@�-q��!?�mjy�@�Б7��ٿ}�La�@!i$~��3@�-q��!?�mjy�@�Б7��ٿ}�La�@!i$~��3@�-q��!?�mjy�@�Б7��ٿ}�La�@!i$~��3@�-q��!?�mjy�@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@��Ў�ٿ��.�(�@)���+4@�:W�!?E�tC甕@�f�f+�ٿy<�Tr��@�
���4@��w��!?������@�K|��ٿ�Ͽ߼�@�J!���3@��R�!?��e��ƕ@�K|��ٿ�Ͽ߼�@�J!���3@��R�!?��e��ƕ@�K|��ٿ�Ͽ߼�@�J!���3@��R�!?��e��ƕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@���?�ٿ~D��i��@C�{#�4@��2��!?sg�xٕ@ް����ٿƱ�����@S���[4@ܨ�nI�!?��4-(~�@ް����ٿƱ�����@S���[4@ܨ�nI�!?��4-(~�@�=z���ٿ��O���@5Í^�4@��)h�!?	6�k��@����ٿ`�s�L�@f3}�Z�3@j&β�!?W�Q��@����ٿ`�s�L�@f3}�Z�3@j&β�!?W�Q��@����ٿ`�s�L�@f3}�Z�3@j&β�!?W�Q��@`�|���ٿ�����@�?V)4@b}����!?����@`�|���ٿ�����@�?V)4@b}����!?����@`�|���ٿ�����@�?V)4@b}����!?����@��˝ٿSFQ�I��@~x�;4@c�ñ��!?l(�H��@��˝ٿSFQ�I��@~x�;4@c�ñ��!?l(�H��@��˝ٿSFQ�I��@~x�;4@c�ñ��!?l(�H��@�R[Fd�ٿ���Sn�@h�394@���!?j�P�3��@�R[Fd�ٿ���Sn�@h�394@���!?j�P�3��@��K�ٿ�!�:ק�@n!��4@?t����!?��x����@��K�ٿ�!�:ק�@n!��4@?t����!?��x����@��K�ٿ�!�:ק�@n!��4@?t����!?��x����@���[�ٿ���Z3��@��F 4@ғ����!?RM��7y�@���[�ٿ���Z3��@��F 4@ғ����!?RM��7y�@���[�ٿ���Z3��@��F 4@ғ����!?RM��7y�@�.�_��ٿ6�V�Sr�@Bx��3@������!?�a���@�.�_��ٿ6�V�Sr�@Bx��3@������!?�a���@�.�_��ٿ6�V�Sr�@Bx��3@������!?�a���@�.�_��ٿ6�V�Sr�@Bx��3@������!?�a���@:��ah�ٿ�����t�@�g�Z�4@4����!?�ә���@z簨d�ٿת +P�@���Ǌ�3@M�R�!?Wt�0ќ�@z簨d�ٿת +P�@���Ǌ�3@M�R�!?Wt�0ќ�@�	O�Ǜٿ��&k'&�@�a���3@�0Sϐ!?��k~�x�@�	O�Ǜٿ��&k'&�@�a���3@�0Sϐ!?��k~�x�@�	O�Ǜٿ��&k'&�@�a���3@�0Sϐ!?��k~�x�@ܓ���ٿ�B��D�@m$fW�3@�o��b�!?dn�M��@ܓ���ٿ�B��D�@m$fW�3@�o��b�!?dn�M��@ܓ���ٿ�B��D�@m$fW�3@�o��b�!?dn�M��@\��4��ٿYv����@ΉlY��3@���ː!?�GB�O*�@\��4��ٿYv����@ΉlY��3@���ː!?�GB�O*�@�_�(�ٿ�\ce��@�pE��3@���pԐ!?x�aW\�@�_�(�ٿ�\ce��@�pE��3@���pԐ!?x�aW\�@�_�(�ٿ�\ce��@�pE��3@���pԐ!?x�aW\�@�_�(�ٿ�\ce��@�pE��3@���pԐ!?x�aW\�@�	�� �ٿ��͖�@�׈��3@�8 ؐ!?��#�4d�@��ը��ٿp�!����@&��%�3@���)��!?�~B�U�@��F"��ٿi�?+�@�ڙ���3@ ^�t��!??��Bh�@��F"��ٿi�?+�@�ڙ���3@ ^�t��!??��Bh�@��F"��ٿi�?+�@�ڙ���3@ ^�t��!??��Bh�@��F"��ٿi�?+�@�ڙ���3@ ^�t��!??��Bh�@Zh�hC�ٿa�Y|��@*H����3@��F!�!?���?�;�@>�s��ٿ��K;��@x^���3@��r���!?FBK�@�� t�ٿH�Y��H�@��}���3@��n�j�!?P�EW�@�� t�ٿH�Y��H�@��}���3@��n�j�!?P�EW�@\�����ٿ�m�ʣ�@
��]	4@�f=��!?�����!�@\�����ٿ�m�ʣ�@
��]	4@�f=��!?�����!�@\�����ٿ�m�ʣ�@
��]	4@�f=��!?�����!�@\�����ٿ�m�ʣ�@
��]	4@�f=��!?�����!�@\�����ٿ�m�ʣ�@
��]	4@�f=��!?�����!�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@x�^�ٿ�8z���@�:���3@�J�!?�y:�6�@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@)�"��ٿ\\�3�U�@{C@L�3@>D�o��!?��D��@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@��R��ٿ�Q�v%�@��h�4@|X�^�!?������@l!�]�ٿ�I)23�@��3�4@L����!?��v�X�@l!�]�ٿ�I)23�@��3�4@L����!?��v�X�@l!�]�ٿ�I)23�@��3�4@L����!?��v�X�@l!�]�ٿ�I)23�@��3�4@L����!?��v�X�@���#��ٿ��<,w*�@�K�w@�3@ߩ=9�!?���ޭ�@���#��ٿ��<,w*�@�K�w@�3@ߩ=9�!?���ޭ�@���#��ٿ��<,w*�@�K�w@�3@ߩ=9�!?���ޭ�@R��ٿP�%V]��@(�.4@K� Y�!?�{�7>
�@R��ٿP�%V]��@(�.4@K� Y�!?�{�7>
�@R��ٿP�%V]��@(�.4@K� Y�!?�{�7>
�@�!I?!�ٿ�x� !�@���%�3@K"N�:�!?���ƕ@�!I?!�ٿ�x� !�@���%�3@K"N�:�!?���ƕ@�!I?!�ٿ�x� !�@���%�3@K"N�:�!?���ƕ@�1vD͝ٿ�*/��q�@2����4@�%�B�!?iM�8eƕ@�1vD͝ٿ�*/��q�@2����4@�%�B�!?iM�8eƕ@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@X�0�,�ٿ �E�&�@��y��/4@=�Q�J�!?��N���@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@�l����ٿ��u���@2w�KJ4@��/x��!?�OXFȕ@z(:/�ٿ�4rn�+�@�M�4@VY���!?��$u֕@z(:/�ٿ�4rn�+�@�M�4@VY���!?��$u֕@z(:/�ٿ�4rn�+�@�M�4@VY���!?��$u֕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@J�3�<�ٿDa�����@��@a��3@!��o�!?w�-r姕@�)q�U�ٿz.�,���@ת$W0�3@	�jL�!?���3�@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@��,�.�ٿW���K�@�Y��1 4@p�LSO�!?��@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@|	|���ٿ��bǦ�@b3
�4@��k�}�!?>��9�@$H�n�ٿ�Mќ��@�[8�r"4@�oK��!?^���R&�@$H�n�ٿ�Mќ��@�[8�r"4@�oK��!?^���R&�@h�Gb�ٿ�C����@�Q�1wJ4@G����!?L��%�@h�Gb�ٿ�C����@�Q�1wJ4@G����!?L��%�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@̥MJ�ٿ*]�o�@Ig���14@���!?�����8�@��i���ٿ�r.�@����4@�۞�!?iM����@��i���ٿ�r.�@����4@�۞�!?iM����@��i���ٿ�r.�@����4@�۞�!?iM����@��i���ٿ�r.�@����4@�۞�!?iM����@��i���ٿ�r.�@����4@�۞�!?iM����@:���ٿ*�cf{��@�#7�\4@'�̌�!?L�(�7�@ǧ[�V�ٿp){����@��aQ{4@�=|N��!?��L�Oޕ@ǧ[�V�ٿp){����@��aQ{4@�=|N��!?��L�Oޕ@\�^ir�ٿ�u²�\�@K���;4@���{�!?>��0��@����.�ٿ�O�U��@�mj�,4@_�x���!?R3�Î��@�c�
�ٿ�~�ڈ��@��,v�3@U�}�l�!?�Q;�1�@�c�
�ٿ�~�ڈ��@��,v�3@U�}�l�!?�Q;�1�@�c�
�ٿ�~�ڈ��@��,v�3@U�}�l�!?�Q;�1�@�c�
�ٿ�~�ڈ��@��,v�3@U�}�l�!?�Q;�1�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@�3�zџٿ/{�h�@��	3�3@.���3�!?7��p+�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@��j��ٿ���O��@px2}��3@DH�!?�*�g-�@J���ٿ�B���`�@_�F��4@��}t�!?3��K�ƕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@���V��ٿ���Q�@a����/4@��s�!?�ϧR�ȕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�[+l�ٿB�Y��@��*�T4@�V�<��!?�@UyЕ@�ԏFѠٿnc��@lP�W4@m%����!?�b�Kk�@�y�T�ٿ؜F�@�9}
`4@�����!?s�sҕ@�y�T�ٿ؜F�@�9}
`4@�����!?s�sҕ@�y�T�ٿ؜F�@�9}
`4@�����!?s�sҕ@�y�T�ٿ؜F�@�9}
`4@�����!?s�sҕ@��-�ٿSx����@�Q�j.4@��_H��!?PV�vM�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@,���ٿ�y����@����4@�E6��!?Z�Ps3�@��$�ٿ�V� C��@��
��4@�m5{l�!?H2�>�@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@���AԖٿO����D�@!�@��4@�޽���!?s[��@�ȹ��ٿ��w��9�@>��A	4@�<��!?��{&w�@�ȹ��ٿ��w��9�@>��A	4@�<��!?��{&w�@�ȹ��ٿ��w��9�@>��A	4@�<��!?��{&w�@����ٿ�p�;���@�`$�3@��L��!?�<+MV�@����ٿ�p�;���@�`$�3@��L��!?�<+MV�@����ٿ�p�;���@�`$�3@��L��!?�<+MV�@놦⠘ٿVշ܀��@u�HA4@?�Fؐ!?�5�ǀ�@놦⠘ٿVշ܀��@u�HA4@?�Fؐ!?�5�ǀ�@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@>�<�ٿ[M�����@�QC04@q�6���!?S����@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@Q��k�ٿ6�+8���@�ﳧq4@b����!?��𓋕@�F�A�ٿ��Ugs�@��y��P4@����.�!?�N��ە@�F�A�ٿ��Ugs�@��y��P4@����.�!?�N��ە@�F�A�ٿ��Ugs�@��y��P4@����.�!?�N��ە@�F�A�ٿ��Ugs�@��y��P4@����.�!?�N��ە@�F�A�ٿ��Ugs�@��y��P4@����.�!?�N��ە@w�\��ٿ*�����@],[�
4@��p0��!?,bP|>�@w�\��ٿ*�����@],[�
4@��p0��!?,bP|>�@w�\��ٿ*�����@],[�
4@��p0��!?,bP|>�@w�\��ٿ*�����@],[�
4@��p0��!?,bP|>�@�O*�ȡٿ��&G�@�:�0�3@^!煟�!?��o�
/�@�O*�ȡٿ��&G�@�:�0�3@^!煟�!?��o�
/�@��`��ٿƞdV�@�*��)4@�����!?�4~J?�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@ؤ�/�ٿ���g?�@���l<4@'�|�!?1)��:�@S�O �ٿ�u۽1m�@��,u�B4@�kA���!?�
���@S�O �ٿ�u۽1m�@��,u�B4@�kA���!?�
���@S�O �ٿ�u۽1m�@��,u�B4@�kA���!?�
���@>�����ٿ�e)��k�@=�}xH4@�Z9�̐!?�= �h�@>�����ٿ�e)��k�@=�}xH4@�Z9�̐!?�= �h�@>�����ٿ�e)��k�@=�}xH4@�Z9�̐!?�= �h�@��R,�ٿ����r�@e�e%'4@��ِ!?7l(�%�@��R,�ٿ����r�@e�e%'4@��ِ!?7l(�%�@��R,�ٿ����r�@e�e%'4@��ِ!?7l(�%�@��R,�ٿ����r�@e�e%'4@��ِ!?7l(�%�@��R,�ٿ����r�@e�e%'4@��ِ!?7l(�%�@R�ژٿ�㊀ݗ�@��-�k4@Ï�v�!? ����@R�ژٿ�㊀ݗ�@��-�k4@Ï�v�!? ����@R�ژٿ�㊀ݗ�@��-�k4@Ï�v�!? ����@R�ژٿ�㊀ݗ�@��-�k4@Ï�v�!? ����@nM�ٿ֠�#ѭ�@ ���4@�����!?����@nM�ٿ֠�#ѭ�@ ���4@�����!?����@nM�ٿ֠�#ѭ�@ ���4@�����!?����@�]r6�ٿ�i�^`��@�E* �3@v�ai�!?J_�?"�@1,KJ)�ٿ�L�1�@=�!��3@`'g�!?W�CP�@1,KJ)�ٿ�L�1�@=�!��3@`'g�!?W�CP�@/"o�١ٿ:<����@�S	4@g�"�*�!? Ì����@/"o�١ٿ:<����@�S	4@g�"�*�!? Ì����@/"o�١ٿ:<����@�S	4@g�"�*�!? Ì����@/"o�١ٿ:<����@�S	4@g�"�*�!? Ì����@/"o�١ٿ:<����@�S	4@g�"�*�!? Ì����@ Otͣٿ:����@
]�|4@)%�;o�!?�
/�A�@HԼ蹣ٿ&��)";�@�nQ9�4@{o�N��!?��/�.�@�u��'�ٿ��_v?�@xM�g��3@x�ӂ�!?��Xǅ��@�=B�ٿ���t�H�@N���.4@/*@S�!?�k�䕖@�=B�ٿ���t�H�@N���.4@/*@S�!?�k�䕖@�=B�ٿ���t�H�@N���.4@/*@S�!?�k�䕖@�=B�ٿ���t�H�@N���.4@/*@S�!?�k�䕖@�=B�ٿ���t�H�@N���.4@/*@S�!?�k�䕖@Ȯh��ٿ��s'ݸ�@9�:4@v{e��!?t����@�^`�ٝٿ�4Y P��@���@J4@��C�!?�U��1��@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@����ٿ�}�p�f�@��v��U4@=��m��!?�6rimE�@���ٿ��B��@zƑ�\4@c3��W�!?(M�ǩ��@9�R�ٿ�I�$ո�@�s!�3@ɲ�Rˏ!?�y4��@9�R�ٿ�I�$ո�@�s!�3@ɲ�Rˏ!?�y4��@,"�o�ٿ�#"��e�@9�$zŭ3@M���^�!?�ë��@^s [�ٿn���*�@So u�3@�p� &�!?K$�V�@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@Q��I`�ٿL�)h��@�w[�d�3@�4cv)�!?oz�"Zѕ@��Ո4�ٿȆڤ��@�P|�f�3@,��b�!?&鬑Ӥ�@��Ո4�ٿȆڤ��@�P|�f�3@,��b�!?&鬑Ӥ�@��Ո4�ٿȆڤ��@�P|�f�3@,��b�!?&鬑Ӥ�@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@>��S��ٿ>q9U��@�!4@������!?�=]���@��+�M�ٿ3r�D�@�F���3@ސ�R��!?{ȆE���@��+�M�ٿ3r�D�@�F���3@ސ�R��!?{ȆE���@M��8D�ٿGn�:���@�e;4@`ߗ9.�!?~%M%v�@M��8D�ٿGn�:���@�e;4@`ߗ9.�!?~%M%v�@M��8D�ٿGn�:���@�e;4@`ߗ9.�!?~%M%v�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@�ૠ�ٿ�c��NY�@��n�� 4@����!?=l��1�@X���ٿ��m�:)�@_�V�Y�3@kPUr�!?Ч���@X���ٿ��m�:)�@_�V�Y�3@kPUr�!?Ч���@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��]c��ٿd�*��@��]��3@���p;�!?g��Kו@��B�m�ٿ�g<vԶ�@A��̓�3@W�f곐!?0�aP�@�_S#k�ٿwE�G_��@�a)��3@;�� Ґ!?04�D�?�@�_S#k�ٿwE�G_��@�a)��3@;�� Ґ!?04�D�?�@�_S#k�ٿwE�G_��@�a)��3@;�� Ґ!?04�D�?�@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@���|�ٿ`���%h�@?^�D�3@�"0(��!?�>�D��@�����ٿ}�0\���@�*b�:�3@%iđ�!?VtH�2�@�����ٿ}�0\���@�*b�:�3@%iđ�!?VtH�2�@�����ٿ}�0\���@�*b�:�3@%iđ�!?VtH�2�@�����ٿ}�0\���@�*b�:�3@%iđ�!?VtH�2�@�A��ٿ0��v7B�@�V��3@����!?�e��Y�@�A��ٿ0��v7B�@�V��3@����!?�e��Y�@�A��ٿ0��v7B�@�V��3@����!?�e��Y�@�A��ٿ0��v7B�@�V��3@����!?�e��Y�@�A��ٿ0��v7B�@�V��3@����!?�e��Y�@������ٿ�f�i��@Jә��3@����!?XEX�@ѕ@������ٿ�f�i��@Jә��3@����!?XEX�@ѕ@������ٿ�f�i��@Jә��3@����!?XEX�@ѕ@ɔ��ٿ1{�l��@;T��3@����i�!?u6da,&�@ɔ��ٿ1{�l��@;T��3@����i�!?u6da,&�@ɔ��ٿ1{�l��@;T��3@����i�!?u6da,&�@ɔ��ٿ1{�l��@;T��3@����i�!?u6da,&�@ɔ��ٿ1{�l��@;T��3@����i�!?u6da,&�@;{�:�ٿ�2bp��@��[��3@�[�!?FC��X�@�8ĸ�ٿ�f���@���)� 4@(3꣐!?sA��@F*�h�ٿ����3��@���5 4@q��D��!?�-`]�T�@F*�h�ٿ����3��@���5 4@q��D��!?�-`]�T�@F*�h�ٿ����3��@���5 4@q��D��!?�-`]�T�@?H1 k�ٿ���>�@B\R4@,J����!?��wp�@?H1 k�ٿ���>�@B\R4@,J����!?��wp�@?H1 k�ٿ���>�@B\R4@,J����!?��wp�@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@I��Mݡٿ*�v�Й�@Xe! �3@����!?��P&��@�r�乤ٿ��ө�f�@�u��4@��(�0�!?4���� �@�r�乤ٿ��ө�f�@�u��4@��(�0�!?4���� �@���c��ٿ�� ��@�OJ�*4@5�Я�!?Ym����@���c��ٿ�� ��@�OJ�*4@5�Я�!?Ym����@���c��ٿ�� ��@�OJ�*4@5�Я�!?Ym����@���c��ٿ�� ��@�OJ�*4@5�Я�!?Ym����@���c��ٿ�� ��@�OJ�*4@5�Я�!?Ym����@��y0V�ٿ<:�5I�@U)��?4@z�d���!?>_�N��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@5� P>�ٿ���G�@sʦ\54@�^ʏ!?kqӴ��@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@��e��ٿy�A��@�12�T4@�Ii�C�!?U���@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@�*��y�ٿ�\ ����@]����64@hw�h1�!?>�v{��@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@��(�(�ٿ��A^k�@����hP4@!�G�s�!?�ܸ/g=�@׷���ٿ���J�@}��=��3@@[m��!?5����@ݗ���ٿi86�w�@��)��4@#�^,b�!?K`G
�@ݗ���ٿi86�w�@��)��4@#�^,b�!?K`G
�@�n)�ߟٿ���"p��@�'��T�3@Lo�Mv�!?�~����@�n)�ߟٿ���"p��@�'��T�3@Lo�Mv�!?�~����@�n)�ߟٿ���"p��@�'��T�3@Lo�Mv�!?�~����@�n)�ߟٿ���"p��@�'��T�3@Lo�Mv�!?�~����@�n)�ߟٿ���"p��@�'��T�3@Lo�Mv�!?�~����@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@K̿;�ٿ�Q��6��@�)>_034@��jr�!?N�p�@���~��ٿ���%�0�@�+N�4@å+��!?�=2�&�@���~��ٿ���%�0�@�+N�4@å+��!?�=2�&�@���~��ٿ���%�0�@�+N�4@å+��!?�=2�&�@���~��ٿ���%�0�@�+N�4@å+��!?�=2�&�@v�cK�ٿ�[�4��@p۰���3@�Ų���!?�nO�u�@v�cK�ٿ�[�4��@p۰���3@�Ų���!?�nO�u�@v�cK�ٿ�[�4��@p۰���3@�Ų���!?�nO�u�@"�ٲg�ٿ�Uـxx�@��:z4@0���!?�����@"�ٲg�ٿ�Uـxx�@��:z4@0���!?�����@"�ٲg�ٿ�Uـxx�@��:z4@0���!?�����@"�ٲg�ٿ�Uـxx�@��:z4@0���!?�����@"�ٲg�ٿ�Uـxx�@��:z4@0���!?�����@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@+���ٿ��D���@g o��4@D 뤘�!?H�@�ߕ@�F��Y�ٿD�^���@�'�C��3@Uu��x�!?[I�XC1�@�F��Y�ٿD�^���@�'�C��3@Uu��x�!?[I�XC1�@�F��Y�ٿD�^���@�'�C��3@Uu��x�!?[I�XC1�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@�Y|`��ٿ�]����@�d�o��3@�"Ft�!?��{/f�@
�m�k�ٿ0A�?q��@�T.!�3@�Q���!?v�u�<�@
�m�k�ٿ0A�?q��@�T.!�3@�Q���!?v�u�<�@
�m�k�ٿ0A�?q��@�T.!�3@�Q���!?v�u�<�@
�m�k�ٿ0A�?q��@�T.!�3@�Q���!?v�u�<�@
�m�k�ٿ0A�?q��@�T.!�3@�Q���!?v�u�<�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@#3P�i�ٿ��7TH�@~T�g>4@�^���!?o�d.(�@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�s:�v�ٿ-���@�q>��A4@a�(�0�!?u6�>��@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@�G��W�ٿL/i���@�wY4@�#�q��!?>a�ȕ@~�2�@�ٿ2~���@�F���54@��6��!?�#(���@~�2�@�ٿ2~���@�F���54@��6��!?�#(���@~�2�@�ٿ2~���@�F���54@��6��!?�#(���@~�2�@�ٿ2~���@�F���54@��6��!?�#(���@���<��ٿC_���@��2��#4@�SV�=�!?$'}����@���<��ٿC_���@��2��#4@�SV�=�!?$'}����@���<��ٿC_���@��2��#4@�SV�=�!?$'}����@���<��ٿC_���@��2��#4@�SV�=�!?$'}����@���<��ٿC_���@��2��#4@�SV�=�!?$'}����@S��W�ٿ��k� ��@�eg��4@�B:���!?��V2-�@S��W�ٿ��k� ��@�eg��4@�B:���!?��V2-�@S��W�ٿ��k� ��@�eg��4@�B:���!?��V2-�@S��W�ٿ��k� ��@�eg��4@�B:���!?��V2-�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@�]�ɡٿxV��Y�@�=QE4@�P���!?���IOF�@����ٿ��G=��@�P��-4@��0D=�!?��D���@����ٿ��G=��@�P��-4@��0D=�!?��D���@����ٿ��G=��@�P��-4@��0D=�!?��D���@sg/f�ٿH���b�@�b+Q�4@�=��!?���m�@sg/f�ٿH���b�@�b+Q�4@�=��!?���m�@sg/f�ٿH���b�@�b+Q�4@�=��!?���m�@wI��k�ٿ�g,~ �@)߭��4@A�+�!?ۚ꫁I�@wI��k�ٿ�g,~ �@)߭��4@A�+�!?ۚ꫁I�@wI��k�ٿ�g,~ �@)߭��4@A�+�!?ۚ꫁I�@wI��k�ٿ�g,~ �@)߭��4@A�+�!?ۚ꫁I�@wI��k�ٿ�g,~ �@)߭��4@A�+�!?ۚ꫁I�@8Di�x�ٿ�f8�Y��@OB��9�3@��ӿ;�!?��G8�@QJB<ޤٿn��{
��@P��H��3@�T`Y�!?Xw��ѕ@�Y:��ٿ��7li�@Υc���3@��K�c�!?Ԓ�u�6�@�Y:��ٿ��7li�@Υc���3@��K�c�!?Ԓ�u�6�@�Y:��ٿ��7li�@Υc���3@��K�c�!?Ԓ�u�6�@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@s�i�ٿy�0�	=�@�ז:��3@��L��!?*pB�ە@�=֠ٿ�i�ס��@���S�3@�q���!?) 4���@�=֠ٿ�i�ס��@���S�3@�q���!?) 4���@�=֠ٿ�i�ס��@���S�3@�q���!?) 4���@o����ٿ�Yq(��@<}�4@/+����!?cbI����@o����ٿ�Yq(��@<}�4@/+����!?cbI����@o����ٿ�Yq(��@<}�4@/+����!?cbI����@o����ٿ�Yq(��@<}�4@/+����!?cbI����@o����ٿ�Yq(��@<}�4@/+����!?cbI����@o����ٿ�Yq(��@<}�4@/+����!?cbI����@,X�ٿ��иW�@E���4@$;gƐ!?R��d�@kqu�\�ٿ�*}p`4�@�4@4@>���!?"�k���@kqu�\�ٿ�*}p`4�@�4@4@>���!?"�k���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�E�q��ٿy��o���@�Tj�)4@o��Y�!?���$���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@�G%s?�ٿI���$5�@c W��4@�2Y(.�!?rB���@���o��ٿcN�%�R�@��'�54@%ρ��!?yz����@��~��ٿG���	-�@�����F4@��+�׏!?��zߕ@��~��ٿG���	-�@�����F4@��+�׏!?��zߕ@��7c�ٿ���^b�@���	94@*
�[�!?.��O�V�@��7c�ٿ���^b�@���	94@*
�[�!?.��O�V�@�N@�c�ٿ��نһ�@��3�'54@x���A�!?b��PDk�@�N@�c�ٿ��نһ�@��3�'54@x���A�!?b��PDk�@.�kY�ٿ���mlE�@�D�E44@��>5�!?����<�@.�kY�ٿ���mlE�@�D�E44@��>5�!?����<�@��6�U�ٿ�Rq#N��@%�Z�4@�*���!?�)`�fi�@��6�U�ٿ�Rq#N��@%�Z�4@�*���!?�)`�fi�@��6�U�ٿ�Rq#N��@%�Z�4@�*���!?�)`�fi�@��6�U�ٿ�Rq#N��@%�Z�4@�*���!?�)`�fi�@��6�U�ٿ�Rq#N��@%�Z�4@�*���!?�)`�fi�@�Tk�Οٿ��H�@���(3*4@QW�.��!?�<J��ƕ@�Tk�Οٿ��H�@���(3*4@QW�.��!?�<J��ƕ@�Tk�Οٿ��H�@���(3*4@QW�.��!?�<J��ƕ@�Tk�Οٿ��H�@���(3*4@QW�.��!?�<J��ƕ@�Tk�Οٿ��H�@���(3*4@QW�.��!?�<J��ƕ@���ٿĹ�|��@]0��!�3@Oթ�.�!?+uiϕ@���ٿĹ�|��@]0��!�3@Oթ�.�!?+uiϕ@�����ٿ�8�����@��-F4@�00L�!?g��/x�@�����ٿ�8�����@��-F4@�00L�!?g��/x�@�����ٿ�8�����@��-F4@�00L�!?g��/x�@�*Lv�ٿsc���@:߄g�3@�lK�'�!?:����K�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@N&�uߠٿ�y��T&�@=�&c�	4@�Zz+/�!?��F�3Z�@�s�z�ٿ7��'��@�>��<4@��m�s�!?6(p�Ny�@�s�z�ٿ7��'��@�>��<4@��m�s�!?6(p�Ny�@�.��ߠٿ�k���@B�,34@9�R�e�!?�	�Ңѕ@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@���i�ٿ��g�R�@�4�o?4@&p��q�!?/EG࢕@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�<.ҠٿM���h��@��
�l,4@F �N��!?~ ���@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@�G#�;�ٿ���`��@js���4@��Y��!?Q��F�@Y�iԛٿ�As�E�@r��4@/��!?r����N�@@j��|�ٿ���eS�@����3@��F-�!?RF;/��@@j��|�ٿ���eS�@����3@��F-�!?RF;/��@�<���ٿ��d��@iŽ�W4@Q�H8�!?��Ƣ�`�@�<���ٿ��d��@iŽ�W4@Q�H8�!?��Ƣ�`�@�<���ٿ��d��@iŽ�W4@Q�H8�!?��Ƣ�`�@��O4ҚٿH��5��@7�M^�"4@&W��D�!?��ꗝ�@��O4ҚٿH��5��@7�M^�"4@&W��D�!?��ꗝ�@��O4ҚٿH��5��@7�M^�"4@&W��D�!?��ꗝ�@�@�/�ٿ�h���J�@�>2)4@/�Z�!?a;�疶�@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@�.	ʟٿ�9"���@ ,�hX4@�zċ�!?HX���@W���ٿ������@�I�h4@���N(�!?�@����@W���ٿ������@�I�h4@���N(�!?�@����@W���ٿ������@�I�h4@���N(�!?�@����@xeo���ٿ<ue�<�@�+�!4@����q�!?�]�ż�@xeo���ٿ<ue�<�@�+�!4@����q�!?�]�ż�@xeo���ٿ<ue�<�@�+�!4@����q�!?�]�ż�@xeo���ٿ<ue�<�@�+�!4@����q�!?�]�ż�@xeo���ٿ<ue�<�@�+�!4@����q�!?�]�ż�@0KX�ٿ�x<����@�P�Y�3@�(B>i�!?O�(���@0KX�ٿ�x<����@�P�Y�3@�(B>i�!?O�(���@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@9�5�֝ٿ:'LI��@��5X(4@��?��!?����H@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�j�|��ٿ���y��@�.�V�*4@���U�!?i���̕@�«�ٿ
���@�@C��Z'4@���"��!?������@�«�ٿ
���@�@C��Z'4@���"��!?������@�����ٿԭu���@Vd	x,74@M�%��!?yV`�Cڕ@�����ٿԭu���@Vd	x,74@M�%��!?yV`�Cڕ@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@�����ٿri�)�@'4a4@	^��b�!?)�SgP,�@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@Z#���ٿRN�"��@x��F�4@�t�g��!?GxҔ?��@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@���[��ٿz{)~E��@�~7���3@2x��u�!?�Xf���@�R�ٿ4�X����@p^dy)4@��%P�!?��$9��@�R�ٿ4�X����@p^dy)4@��%P�!?��$9��@�R�ٿ4�X����@p^dy)4@��%P�!?��$9��@�hC�ٿ�C� g�@3��D�74@�iۉ�!?�ͨߕ@�hC�ٿ�C� g�@3��D�74@�iۉ�!?�ͨߕ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@/����ٿ�D[���@P��!�D4@ޒjM�!?)A�c&Õ@�K�O�ٿ���U��@��BĂ54@/H�j�!?wiLW��@�K�O�ٿ���U��@��BĂ54@/H�j�!?wiLW��@#����ٿ�a�$��@!���g#4@��溍�!?�^��L��@#����ٿ�a�$��@!���g#4@��溍�!?�^��L��@(Ѵ�0�ٿ|� �@��Ծ.4@׿�"q�!?��c���@0��ٿ��ں��@�82�%4@��G%M�!?��lSK�@0��ٿ��ں��@�82�%4@��G%M�!?��lSK�@0��ٿ��ں��@�82�%4@��G%M�!?��lSK�@��G�ٿ�k�i�n�@,l�O/4@�`C��!?7�����@��G�ٿ�k�i�n�@,l�O/4@�`C��!?7�����@��G�ٿ�k�i�n�@,l�O/4@�`C��!?7�����@��G�ٿ�k�i�n�@,l�O/4@�`C��!?7�����@��G�ٿ�k�i�n�@,l�O/4@�`C��!?7�����@l��):�ٿ3b����@BW����3@�<o)Đ!?�kz�왕@#9�y�ٿ������@����B4@�(�d�!?�1��ɕ@#9�y�ٿ������@����B4@�(�d�!?�1��ɕ@#9�y�ٿ������@����B4@�(�d�!?�1��ɕ@�u܁�ٿ��)��c�@%0��!4@�.�!?�V׺��@�u܁�ٿ��)��c�@%0��!4@�.�!?�V׺��@�u܁�ٿ��)��c�@%0��!4@�.�!?�V׺��@�>�uD�ٿoD�����@e��;4@Y�6�!?o�:����@�>�uD�ٿoD�����@e��;4@Y�6�!?o�:����@�<�3��ٿW�<+�f�@Y�R�[4@\�<ZB�!?J�VX�ؕ@�<�3��ٿW�<+�f�@Y�R�[4@\�<ZB�!?J�VX�ؕ@�<�3��ٿW�<+�f�@Y�R�[4@\�<ZB�!?J�VX�ؕ@Cm<�S�ٿP4WG�@��c��?4@3u��T�!?�<@c�@Cm<�S�ٿP4WG�@��c��?4@3u��T�!?�<@c�@�s��5�ٿc�N����@|�2��,4@X�� ��!?� ���@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@ 0����ٿZ,��I�@u�<TO=4@Ő�<��!?R�F��@�z)��ٿ��al��@����04@�����!?���W�ٕ@�z)��ٿ��al��@����04@�����!?���W�ٕ@�z)��ٿ��al��@����04@�����!?���W�ٕ@�z)��ٿ��al��@����04@�����!?���W�ٕ@:b���ٿ��4��A�@�S�8G"4@qQ���!?��O��@:b���ٿ��4��A�@�S�8G"4@qQ���!?��O��@���X��ٿ�X,��w�@h!�HD4@�C%�~�!?%�����@���X��ٿ�X,��w�@h!�HD4@�C%�~�!?%�����@�l*���ٿ��^ؕn�@G��[l4@��7�o�!?�A���@�l*���ٿ��^ؕn�@G��[l4@��7�o�!?�A���@�l*���ٿ��^ؕn�@G��[l4@��7�o�!?�A���@�l*���ٿ��^ؕn�@G��[l4@��7�o�!?�A���@�l*���ٿ��^ؕn�@G��[l4@��7�o�!?�A���@��ط�ٿt;�o��@pu��4@���k��!?}��F�ו@��ط�ٿt;�o��@pu��4@���k��!?}��F�ו@��ط�ٿt;�o��@pu��4@���k��!?}��F�ו@��ط�ٿt;�o��@pu��4@���k��!?}��F�ו@�z`�6�ٿ�1&$�@��#ٮ�3@di�Y�!?��)��@�z`�6�ٿ�1&$�@��#ٮ�3@di�Y�!?��)��@�8#�C�ٿ��
���@�q�!��3@'�&W��!?��63�Õ@�lH�Q�ٿ�k�ȍ�@&���3@�7���!?�4Iw��@�lH�Q�ٿ�k�ȍ�@&���3@�7���!?�4Iw��@G��؛ٿ�ٳ�a�@��c�H4@��/��!?� \0}ޕ@G��؛ٿ�ٳ�a�@��c�H4@��/��!?� \0}ޕ@�&V<��ٿ*jQ���@ܷ4@'���!?�{�ӹ�@�B%<�ٿ�$2r%C�@��Sg�
4@N��ߚ�!?n1 ��@�B%<�ٿ�$2r%C�@��Sg�
4@N��ߚ�!?n1 ��@�B%<�ٿ�$2r%C�@��Sg�
4@N��ߚ�!?n1 ��@�B%<�ٿ�$2r%C�@��Sg�
4@N��ߚ�!?n1 ��@�B%<�ٿ�$2r%C�@��Sg�
4@N��ߚ�!?n1 ��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����g�ٿw�j=��@}���3@*q��!?Nc��@����Оٿ�:�O��@Z"
���3@���^�!?,MBQ�@����Оٿ�:�O��@Z"
���3@���^�!?,MBQ�@����Оٿ�:�O��@Z"
���3@���^�!?,MBQ�@����Оٿ�:�O��@Z"
���3@���^�!?,MBQ�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@�I^��ٿ�O���@�`~5��3@A��.E�!?���l�V�@A<�Țٿ�~�/�r�@jݟy�4@���a4�!?�A�q�@A<�Țٿ�~�/�r�@jݟy�4@���a4�!?�A�q�@A<�Țٿ�~�/�r�@jݟy�4@���a4�!?�A�q�@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@��Y�ٿ0�P�"_�@�<�F�"4@��;�3�!?��]���@�X�K��ٿ0�Հ��@�7rC4@to�!?�b_���@�X�K��ٿ0�Հ��@�7rC4@to�!?�b_���@�X�K��ٿ0�Հ��@�7rC4@to�!?�b_���@=r�.R�ٿ���(N4�@�X�@�%4@�Y_\|�!?��&��ɕ@=r�.R�ٿ���(N4�@�X�@�%4@�Y_\|�!?��&��ɕ@��_��ٿ�0B���@��w�4@*͒�M�!?ViC�tו@��_��ٿ�0B���@��w�4@*͒�M�!?ViC�tו@���Úٿ��!ʴy�@�-��44@f;�O��!?sޤ�d�@���Úٿ��!ʴy�@�-��44@f;�O��!?sޤ�d�@�$Öٿ(	�g�@��L��*4@8y��!?��_S�Ε@�$Öٿ(	�g�@��L��*4@8y��!?��_S�Ε@9SEg_�ٿ�0�B�@�=r4@�V�!?dZ 
�@K�[�v�ٿ/q�b�@�#�ñ�3@��ܔ3�!?��B(��@K�[�v�ٿ/q�b�@�#�ñ�3@��ܔ3�!?��B(��@K�[�v�ٿ/q�b�@�#�ñ�3@��ܔ3�!?��B(��@K�[�v�ٿ/q�b�@�#�ñ�3@��ܔ3�!?��B(��@d�Ģ��ٿ�V*���@�0�n4@^�ν&�!?����e��@�x��*�ٿN�$���@���E�3@�8$���!?���5��@�x��*�ٿN�$���@���E�3@�8$���!?���5��@�x��*�ٿN�$���@���E�3@�8$���!?���5��@�x��*�ٿN�$���@���E�3@�8$���!?���5��@�x��*�ٿN�$���@���E�3@�8$���!?���5��@\P��ٿS��`�O�@<(~�24@XRu��!?	Gr�ѕ@�1��A�ٿ}��*�@s����24@����!?H0��@�1��A�ٿ}��*�@s����24@����!?H0��@�1��A�ٿ}��*�@s����24@����!?H0��@�1��A�ٿ}��*�@s����24@����!?H0��@�1��A�ٿ}��*�@s����24@����!?H0��@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�e�w}�ٿ� �(�@Y�hvF4@�䨪��!?��`��m�@�E��v�ٿe�t�*e�@��;4@}���5�!?����}3�@�E��v�ٿe�t�*e�@��;4@}���5�!?����}3�@�E��v�ٿe�t�*e�@��;4@}���5�!?����}3�@�E��v�ٿe�t�*e�@��;4@}���5�!?����}3�@�tB�M�ٿ�čL��@���z�3@��Zv^�!?)33<(\�@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@"�R�ٿ��6�0D�@�w9���3@��ȃp�!?�T�:���@X���b�ٿ��!��@�O����3@��G�ɐ!?;v����@v��[�ٿ�����@}IDgd	4@���ڐ!?},�[�v�@�����ٿ���C[[�@y4�	,�3@bQ�3v�!?E��ήÕ@��Y�ٿ6�p��@Χ��i4@�{�u�!?�j��ܕ@h��a�ٿ���\r �@�I}�4@���D�!?52�abQ�@h��a�ٿ���\r �@�I}�4@���D�!?52�abQ�@h��a�ٿ���\r �@�I}�4@���D�!?52�abQ�@h��a�ٿ���\r �@�I}�4@���D�!?52�abQ�@h��a�ٿ���\r �@�I}�4@���D�!?52�abQ�@��̚ٿ)C��x��@���U4@�KT�!?@p�2
#�@�.W�ٿ��P9-�@��EF�C4@Gs�!?�!�=�@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@��S�i�ٿ���u	��@Y�  �?4@I�eJ�!?�׽�֕@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@�+�3��ٿ��3��@X��14@�!4ɓ�!?o�MrЕ@H�r�?�ٿ�H�_�:�@�mI߂?4@����[�!?�?|)ҕ@|a5֜�ٿ �E���@wD��4@�M%q;�!?-���@|a5֜�ٿ �E���@wD��4@�M%q;�!?-���@m�K��ٿ� [b��@#GH�$+4@�}�z(�!?N�40��@�Yf�5�ٿ��v���@F��4@*H]GS�!?���Bj��@�Yf�5�ٿ��v���@F��4@*H]GS�!?���Bj��@������ٿ��r��@�0�v��3@>��=�!?5���@�VZ��ٿ����@J	^�u4@°-�f�!?� �n�@�VZ��ٿ����@J	^�u4@°-�f�!?� �n�@�VZ��ٿ����@J	^�u4@°-�f�!?� �n�@�VZ��ٿ����@J	^�u4@°-�f�!?� �n�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@�Y:�ٿ�P:hOl�@��y��4@z3-�K�!?'���Z
�@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@8��:�ٿ<ʗ~\�@�k!]�3@�q�g�!?p����@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@��L�X�ٿ��_���@0��H�3@{�>!r�!?E:L%��@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�QE��ٿ[ꃡ��@ˎ(m	4@�����!?�j¦� �@�(3���ٿe��E;�@DS	'��3@	2�oG�!?�;����@3b�z�ٿ8������@�\�O4@6t��]�!?�H@"�@3b�z�ٿ8������@�\�O4@6t��]�!?�H@"�@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��!�ٿ��^�H�@�嚪~4@IA���!?�I >��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@��W��ٿa�]�X�@SX�7��3@��`mH�!?�C��~��@K/�.�ٿK���U-�@��"ef�3@��ok�!?�*�ҕ@K/�.�ٿK���U-�@��"ef�3@��ok�!?�*�ҕ@K/�.�ٿK���U-�@��"ef�3@��ok�!?�*�ҕ@�y&9Z�ٿ?��Y��@�J����3@�aޜ4�!?��h�ĕ@���ׇ�ٿ���(��@�m��3@�B��6�!?z�>���@���ׇ�ٿ���(��@�m��3@�B��6�!?z�>���@���ׇ�ٿ���(��@�m��3@�B��6�!?z�>���@���ׇ�ٿ���(��@�m��3@�B��6�!?z�>���@��_TI�ٿp�����@vD0Ӿ�3@'`�?R�!?z4��@��_TI�ٿp�����@vD0Ӿ�3@'`�?R�!?z4��@�*	�Ǜٿ	Q���@M���3@�1$��!?-�\@
�@7n��ٿt��A�-�@��=�:�3@��F���!?#Y�}ҷ�@7n��ٿt��A�-�@��=�:�3@��F���!?#Y�}ҷ�@7n��ٿt��A�-�@��=�:�3@��F���!?#Y�}ҷ�@7n��ٿt��A�-�@��=�:�3@��F���!?#Y�}ҷ�@(��N#�ٿ�ѱ���@��$4@��u�n�!?���n��@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�^�*��ٿ�bv_D�@����3@��{�!?��-�|p�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@�wO+�ٿ��m�h��@�6	4@lM��`�!?���C�t�@��k��ٿ1��z��@wٔ VC4@��B��!?k���{h�@��k��ٿ1��z��@wٔ VC4@��B��!?k���{h�@�qk~@�ٿ@!�g�@kW���Y4@A�ߏ!?	?���Ǖ@)���|�ٿ�$ߎs�@�kŔ^C4@"~g��!?c��t���@�X�,�ٿ���~���@^c�I�4@QS�T�!?�����@�X�,�ٿ���~���@^c�I�4@QS�T�!?�����@j���^�ٿ|�Ӊo��@�Y`��3@�7�@�!?��18F��@j���^�ٿ|�Ӊo��@�Y`��3@�7�@�!?��18F��@j���^�ٿ|�Ӊo��@�Y`��3@�7�@�!?��18F��@j���^�ٿ|�Ӊo��@�Y`��3@�7�@�!?��18F��@��_Z�ٿH�I$�L�@$�Ga9�3@6;��!?R�a���@��_Z�ٿH�I$�L�@$�Ga9�3@6;��!?R�a���@��_Z�ٿH�I$�L�@$�Ga9�3@6;��!?R�a���@��_Z�ٿH�I$�L�@$�Ga9�3@6;��!?R�a���@��ڇ��ٿhQ,���@7�; �=4@��܏!?�I��x�@��ڇ��ٿhQ,���@7�; �=4@��܏!?�I��x�@�ӑ"N�ٿ[L����@�Ø��4@�nf�!?8��@�ӑ"N�ٿ[L����@�Ø��4@�nf�!?8��@�ӑ"N�ٿ[L����@�Ø��4@�nf�!?8��@�ӑ"N�ٿ[L����@�Ø��4@�nf�!?8��@�ӑ"N�ٿ[L����@�Ø��4@�nf�!?8��@.}��'�ٿ������@��P+04@6�K
��!?X�.W��@.}��'�ٿ������@��P+04@6�K
��!?X�.W��@�Ȥe�ٿ^sER�q�@@��04@��x�!?��e'�L�@¯1F�ٿ븉�~��@Y���N4@e�Cw�!?k��V�A�@¯1F�ٿ븉�~��@Y���N4@e�Cw�!?k��V�A�@E��y�ٿ�=�����@)�9Mes4@�����!?O[���@E��y�ٿ�=�����@)�9Mes4@�����!?O[���@E��y�ٿ�=�����@)�9Mes4@�����!?O[���@��]�֟ٿ���@e�>7R4@�0%���!?L{]��@��]�֟ٿ���@e�>7R4@�0%���!?L{]��@��]�֟ٿ���@e�>7R4@�0%���!?L{]��@��I�ٿ������@�=��l4@�;���!?�Dp⁖@��I�ٿ������@�=��l4@�;���!?�Dp⁖@��I�ٿ������@�=��l4@�;���!?�Dp⁖@�>���ٿ ~��i7�@z+K�DP4@��� >�!?8�gGg6�@�>���ٿ ~��i7�@z+K�DP4@��� >�!?8�gGg6�@c�o���ٿJm:�]��@/��I4@"���!?Z�3���@c�o���ٿJm:�]��@/��I4@"���!?Z�3���@c�o���ٿJm:�]��@/��I4@"���!?Z�3���@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@V��J�ٿQ�X ّ�@:�434@�%�!?}��0�@��b�ٿ%��pd�@�i����3@���[�!?_�W��k�@LP����ٿ�%�����@1���Y4@��6�e�!?8d=��%�@LP����ٿ�%�����@1���Y4@��6�e�!?8d=��%�@LP����ٿ�%�����@1���Y4@��6�e�!?8d=��%�@LP����ٿ�%�����@1���Y4@��6�e�!?8d=��%�@LP����ٿ�%�����@1���Y4@��6�e�!?8d=��%�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@�u���ٿ�Ѐp��@�S޵r4@YrQO�!?5�)=/3�@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@)���̠ٿNrſ�@�:�%�4@�#'b�!?(6�����@��>���ٿm���@�P4�[�3@��d�9�!?{ښ��@ޜ){D�ٿu1X��s�@��E��3@ ��,�!?�RvK��@ޜ){D�ٿu1X��s�@��E��3@ ��,�!?�RvK��@ޜ){D�ٿu1X��s�@��E��3@ ��,�!?�RvK��@��a��ٿ�?�^���@�X狕�3@�d�E�!?cYt�͕@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@��!C�ٿ�o�N���@Pngj�+4@�]�g�!?��_�ʕ@�<s䒜ٿ� 5�{�@B+���4@���-�!?U�+?H�@�<s䒜ٿ� 5�{�@B+���4@���-�!?U�+?H�@�<s䒜ٿ� 5�{�@B+���4@���-�!?U�+?H�@ې���ٿL�%���@y<f�*4@<�VzV�!?�\ת6.�@ې���ٿL�%���@y<f�*4@<�VzV�!?�\ת6.�@ې���ٿL�%���@y<f�*4@<�VzV�!?�\ת6.�@xTAԙٿD���^��@��} -4@3$��y�!?�4�@xTAԙٿD���^��@��} -4@3$��y�!?�4�@xTAԙٿD���^��@��} -4@3$��y�!?�4�@īR���ٿw$h���@�ml54@���L��!?*�>���@īR���ٿw$h���@�ml54@���L��!?*�>���@īR���ٿw$h���@�ml54@���L��!?*�>���@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@��0<�ٿ� ��n�@�b���3@����ʐ!?�k�}�֕@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@����ٿ�d�3�@�`ڍ�14@`�*��!?271:�@p���ٿC1B;��@�����54@i��j��!?Bh���ٕ@p���ٿC1B;��@�����54@i��j��!?Bh���ٕ@p���ٿC1B;��@�����54@i��j��!?Bh���ٕ@p���ٿC1B;��@�����54@i��j��!?Bh���ٕ@H��6�ٿ�i̙��@�Q���+4@�
���!?�7z�@H��6�ٿ�i̙��@�Q���+4@�
���!?�7z�@H��6�ٿ�i̙��@�Q���+4@�
���!?�7z�@H��6�ٿ�i̙��@�Q���+4@�
���!?�7z�@H��6�ٿ�i̙��@�Q���+4@�
���!?�7z�@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@�vֱ	�ٿ����$=�@B�@^94@��?1b�!?U�c��@��[�ٿ�^��@<���W)4@���f��!?C�P�K��@�����ٿ�nO>�@gT�:"4@S�D�b�!?��s�u�@�����ٿ�nO>�@gT�:"4@S�D�b�!?��s�u�@�����ٿ�nO>�@gT�:"4@S�D�b�!?��s�u�@�����ٿ�nO>�@gT�:"4@S�D�b�!?��s�u�@c��E��ٿb�|t��@`��Z4@�N勐!?�@�)�@0ny��ٿe����@�@
�gK4@/�F��!?y�	ƱD�@0ny��ٿe����@�@
�gK4@/�F��!?y�	ƱD�@0ny��ٿe����@�@
�gK4@/�F��!?y�	ƱD�@���ٿ�:����@��|�?44@|i:���!?C=� ܕ@���ٿ�:����@��|�?44@|i:���!?C=� ܕ@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@��g�ٿ5���s�@�6��BL4@,�F�!?���S��@'�8���ٿ@"(M���@c?{B�4@{��r�!?��� �@'�8���ٿ@"(M���@c?{B�4@{��r�!?��� �@'�8���ٿ@"(M���@c?{B�4@{��r�!?��� �@Fa��M�ٿ��5���@�WDM4@Ǳ�j|�!?�y�Pc��@Fa��M�ٿ��5���@�WDM4@Ǳ�j|�!?�y�Pc��@Fa��M�ٿ��5���@�WDM4@Ǳ�j|�!?�y�Pc��@�K$��ٿ�'y���@K�E��24@k�6mk�!?y��~��@�K$��ٿ�'y���@K�E��24@k�6mk�!?y��~��@�K$��ٿ�'y���@K�E��24@k�6mk�!?y��~��@� ����ٿ� ���@���m94@��/�!?�,Mlzߕ@� ����ٿ� ���@���m94@��/�!?�,Mlzߕ@yUj��ٿC�8m��@P�}�4@7:���!?+y_N�ŕ@yUj��ٿC�8m��@P�}�4@7:���!?+y_N�ŕ@EjϚ3�ٿk�����@0e{|+4@��A�I�!?v!(Ϳ=�@U����ٿ嬆@\��@���
4@���(y�!?>܂!9��@U����ٿ嬆@\��@���
4@���(y�!?>܂!9��@U����ٿ嬆@\��@���
4@���(y�!?>܂!9��@U����ٿ嬆@\��@���
4@���(y�!?>܂!9��@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@�}�신ٿ�ѯ7s��@����4@+D\�!?rEgFە@���t��ٿԖOJ��@�b.?��3@va�!?�,�m̕@���t��ٿԖOJ��@�b.?��3@va�!?�,�m̕@���t��ٿԖOJ��@�b.?��3@va�!?�,�m̕@���t��ٿԖOJ��@�b.?��3@va�!?�,�m̕@���t��ٿԖOJ��@�b.?��3@va�!?�,�m̕@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@��� �ٿ�����@~cXE4@A
[�\�!?7X�(��@�{]�ٿ&|��X�@h���3@bs_��!?G[r+��@�{]�ٿ&|��X�@h���3@bs_��!?G[r+��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@���Ϝ�ٿ\�/��@��(4@��3+�!?tϕN��@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@w��i�ٿV�>:��@�>v�#A4@m�]���!?���}Y)�@MIb��ٿ
�����@ֱ��!A4@���a�!??�w�`�@MIb��ٿ
�����@ֱ��!A4@���a�!??�w�`�@MIb��ٿ
�����@ֱ��!A4@���a�!??�w�`�@MIb��ٿ
�����@ֱ��!A4@���a�!??�w�`�@�km5�ٿ�3x���@Yߦ5��3@����!?n*P;%;�@NI�D�ٿQ����j�@Fv@c4@�����!?���X��@��.��ٿ�_RY��@b�YP	�3@���]�!?����
q�@��.��ٿ�_RY��@b�YP	�3@���]�!?����
q�@��.��ٿ�_RY��@b�YP	�3@���]�!?����
q�@��.��ٿ�_RY��@b�YP	�3@���]�!?����
q�@��.��ٿ�_RY��@b�YP	�3@���]�!?����
q�@̕��}�ٿ&�U���@H�x:4@,m� ��!?V��u�@̕��}�ٿ&�U���@H�x:4@,m� ��!?V��u�@̕��}�ٿ&�U���@H�x:4@,m� ��!?V��u�@̕��}�ٿ&�U���@H�x:4@,m� ��!?V��u�@���*>�ٿ��0��+�@�?�)4@@w%�j�!?�<0o�T�@~���ٿ�W�@�o��F4@�M�]�!?���^D7�@~���ٿ�W�@�o��F4@�M�]�!?���^D7�@�����ٿ)��U��@�n1i�W4@}d8G�!?�v�/�@@,���ٿG��Qkk�@X&���3@P W7C�!?F���@@,���ٿG��Qkk�@X&���3@P W7C�!?F���@-�kea�ٿܬ(v��@=�=<i4@d�<�!?a<ued��@-�kea�ٿܬ(v��@=�=<i4@d�<�!?a<ued��@-�kea�ٿܬ(v��@=�=<i4@d�<�!?a<ued��@OJD��ٿӇI���@����,4@v��(�!?�;��ߕ@OJD��ٿӇI���@����,4@v��(�!?�;��ߕ@OJD��ٿӇI���@����,4@v��(�!?�;��ߕ@OJD��ٿӇI���@����,4@v��(�!?�;��ߕ@OJD��ٿӇI���@����,4@v��(�!?�;��ߕ@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@�����ٿI������@܏U5q4@�ʬ�>�!?�y@z��@X�r���ٿ��1B^�@pZ!��'4@��ޙ�!?������@X�r���ٿ��1B^�@pZ!��'4@��ޙ�!?������@X�r���ٿ��1B^�@pZ!��'4@��ޙ�!?������@X�r���ٿ��1B^�@pZ!��'4@��ޙ�!?������@X�r���ٿ��1B^�@pZ!��'4@��ޙ�!?������@X�v�W�ٿ>{���@/6��54@�����!?���S��@X�v�W�ٿ>{���@/6��54@�����!?���S��@���y�ٿ��t���@�\{�H
4@Y�w���!?�ä�u�@���y�ٿ��t���@�\{�H
4@Y�w���!?�ä�u�@���y�ٿ��t���@�\{�H
4@Y�w���!?�ä�u�@���y�ٿ��t���@�\{�H
4@Y�w���!?�ä�u�@E����ٿ���Y��@�'y���3@O�\/�!?t �*�Е@��K��ٿ ���_��@�P� ��3@��No�!? ���H�@��K��ٿ ���_��@�P� ��3@��No�!? ���H�@�y<t�ٿO/0�c��@mt~L94@4��'k�!?R$O)_�@�y<t�ٿO/0�c��@mt~L94@4��'k�!?R$O)_�@�(�Y�ٿ��[���@Ԁ�@�D4@���?o�!?�_B��/�@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@��sA�ٿ�X;M]@�@yp��A94@U	�v�!?���Bٕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@s���ٿ:2+���@&��4@�A�Su�!?D|ݮ[ܕ@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@+^�:�ٿbmA��R�@�4
|��3@~§pr�!?k�(��
�@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@cM\[�ٿ�d��Q��@"�̉��3@Q��W�!?�{`k�ڕ@,�wqp�ٿ�s<�>�@����3@+��M�!?}Rs��@,�wqp�ٿ�s<�>�@����3@+��M�!?}Rs��@,�wqp�ٿ�s<�>�@����3@+��M�!?}Rs��@,�wqp�ٿ�s<�>�@����3@+��M�!?}Rs��@,�wqp�ٿ�s<�>�@����3@+��M�!?}Rs��@�����ٿ�B�i1�@wH(��#4@jl�R�!?M�1u�6�@�����ٿ�B�i1�@wH(��#4@jl�R�!?M�1u�6�@�����ٿ�B�i1�@wH(��#4@jl�R�!?M�1u�6�@�����ٿ�B�i1�@wH(��#4@jl�R�!?M�1u�6�@�����ٿ�B�i1�@wH(��#4@jl�R�!?M�1u�6�@PZ%�X�ٿ_��9��@cMM+F4@Y�7�:�!?�6R5�@�����ٿ9=��j�@3:@?WW4@���3�!?X(�N��@�����ٿ9=��j�@3:@?WW4@���3�!?X(�N��@ �ԎΟٿbY����@��ˀ�/4@�v�q�!?�MX����@ �ԎΟٿbY����@��ˀ�/4@�v�q�!?�MX����@���ٿ-���@8�V{�U4@j��S�!?>-�����@���ٿ-���@8�V{�U4@j��S�!?>-�����@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@V�.ly�ٿ���PP�@�4���[4@���B��!?����£�@�𬞜ٿ�+���+�@e蕒b4@���\�!?��h����@�𬞜ٿ�+���+�@e蕒b4@���\�!?��h����@�𬞜ٿ�+���+�@e蕒b4@���\�!?��h����@��m3�ٿ��K��@X���e4@�g �u�!?����O��@��m3�ٿ��K��@X���e4@�g �u�!?����O��@��m3�ٿ��K��@X���e4@�g �u�!?����O��@��m3�ٿ��K��@X���e4@�g �u�!?����O��@��m3�ٿ��K��@X���e4@�g �u�!?����O��@��m3�ٿ��K��@X���e4@�g �u�!?����O��@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@6��6��ٿ[�ڙGf�@$y��U4@������!?̇�a���@�W����ٿ/��_�n�@�x���,4@`Q�Ԑ!?l}�0쬕@�W����ٿ/��_�n�@�x���,4@`Q�Ԑ!?l}�0쬕@�W����ٿ/��_�n�@�x���,4@`Q�Ԑ!?l}�0쬕@����F�ٿ���@$4/��3@Jc��6�!?
y��*�@����F�ٿ���@$4/��3@Jc��6�!?
y��*�@����F�ٿ���@$4/��3@Jc��6�!?
y��*�@cDA}�ٿ% Cy�C�@~��s4@c{�N�!?S�:w%�@cDA}�ٿ% Cy�C�@~��s4@c{�N�!?S�:w%�@cDA}�ٿ% Cy�C�@~��s4@c{�N�!?S�:w%�@cDA}�ٿ% Cy�C�@~��s4@c{�N�!?S�:w%�@�dt~Q�ٿ����m��@#��Ӄ4@u`3b�!?����J�@�dt~Q�ٿ����m��@#��Ӄ4@u`3b�!?����J�@������ٿ�^���@�	�xw�3@x(W=�!?��No���@������ٿ�^���@�	�xw�3@x(W=�!?��No���@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@����ٿ��9@�@�X��%%4@�.��B�!?��n�.��@�P����ٿ2k8�^��@fJc��3@K�)�8�!?��nJ��@�P����ٿ2k8�^��@fJc��3@K�)�8�!?��nJ��@�P����ٿ2k8�^��@fJc��3@K�)�8�!?��nJ��@�P����ٿ2k8�^��@fJc��3@K�)�8�!?��nJ��@�P����ٿ2k8�^��@fJc��3@K�)�8�!?��nJ��@�`��(�ٿ�2�6_��@�|֛�3@l^��*�!?����/�@�`��(�ٿ�2�6_��@�|֛�3@l^��*�!?����/�@��`Lޜٿ쇾�K�@�g�f�3@�-&�O�!?�f���@��`Lޜٿ쇾�K�@�g�f�3@�-&�O�!?�f���@�Uۥ.�ٿ����@���VP�3@)*T猐!?���O�@�Uۥ.�ٿ����@���VP�3@)*T猐!?���O�@�Uۥ.�ٿ����@���VP�3@)*T猐!?���O�@�Uۥ.�ٿ����@���VP�3@)*T猐!?���O�@�e}dۚٿ%"Jy��@�H�[��3@�D�U�!?)�0h
�@�J�;�ٿ���?{�@Z�����3@�k(�}�!?���Fk�@�J�;�ٿ���?{�@Z�����3@�k(�}�!?���Fk�@����ٿ�lb��@��t��W4@�gė��!?Cꔒ��@����ٿ�lb��@��t��W4@�gė��!?Cꔒ��@����ٿ�lb��@��t��W4@�gė��!?Cꔒ��@E�Ƶx�ٿ�Uת�@H��N4@F�T��!?_n�;bϕ@E�Ƶx�ٿ�Uת�@H��N4@F�T��!?_n�;bϕ@E�Ƶx�ٿ�Uת�@H��N4@F�T��!?_n�;bϕ@�U�G�ٿQg^�[��@U�^�*4@����B�!?{�E�$�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@r"`�k�ٿaJ6%uR�@Wde�&4@�w�Z�!?}q�"�@-�����ٿ$������@�P�˴04@�c0J�!?G�~�:J�@-�����ٿ$������@�P�˴04@�c0J�!?G�~�:J�@-�����ٿ$������@�P�˴04@�c0J�!?G�~�:J�@-�����ٿ$������@�P�˴04@�c0J�!?G�~�:J�@�ᖟٿL��I��@_"h�S�3@2���"�!?˔�!R�@k!	_��ٿ���'�@�����L4@!a���!?��Z��@k!	_��ٿ���'�@�����L4@!a���!?��Z��@�$��ٿ����a��@���H4@XA��U�!?jo�����@�$��ٿ����a��@���H4@XA��U�!?jo�����@�$��ٿ����a��@���H4@XA��U�!?jo�����@��!�ٿ5'��@�Wjfy4@��l#>�!?`��C)�@��!�ٿ5'��@�Wjfy4@��l#>�!?`��C)�@��!�ٿ5'��@�Wjfy4@��l#>�!?`��C)�@���ٿr�	����@/\ �*I4@M�Y�@�!?=�$�f�@���ٿr�	����@/\ �*I4@M�Y�@�!?=�$�f�@���ٿr�	����@/\ �*I4@M�Y�@�!?=�$�f�@���ٿr�	����@/\ �*I4@M�Y�@�!?=�$�f�@��)��ٿ� 硥��@�	\\<4@�~�8�!?��u$C�@��)��ٿ� 硥��@�	\\<4@�~�8�!?��u$C�@��)��ٿ� 硥��@�	\\<4@�~�8�!?��u$C�@ps�Cژٿu�����@դF�3@�Fg5�!?)��0ߕ@ps�Cژٿu�����@դF�3@�Fg5�!?)��0ߕ@��W�ٿ��!+�@�\'4@gB�$;�!?����K��@��W�ٿ��!+�@�\'4@gB�$;�!?����K��@��W�ٿ��!+�@�\'4@gB�$;�!?����K��@�Ԋn��ٿ�{B�0��@�����4@kQ=ZW�!?v�B�?��@�;+�"�ٿ	�|No�@����94@�y<�!?
̃�aە@Ԝ���ٿ�~R�L�@�!J�k4@���2�!?d�'뵼�@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@��!I�ٿ��IL�@��u�3@����@�!?�� Е@rNr�ۗٿ\8�u�@GDBk��3@,�7�Y�!?h�rN$�@rNr�ۗٿ\8�u�@GDBk��3@,�7�Y�!?h�rN$�@rNr�ۗٿ\8�u�@GDBk��3@,�7�Y�!?h�rN$�@+�x^v�ٿ�ы���@]�G���3@l��0I�!?�~����@+�x^v�ٿ�ы���@]�G���3@l��0I�!?�~����@+�x^v�ٿ�ы���@]�G���3@l��0I�!?�~����@+�x^v�ٿ�ы���@]�G���3@l��0I�!?�~����@r0ݰ�ٿC�n�2�@O�e��44@���1��!?F�xz��@r0ݰ�ٿC�n�2�@O�e��44@���1��!?F�xz��@���F�ٿ���@�+�׽<4@�@<��!?o;�"t�@����ٿQ���m�@z����4@��
9�!?oe��{�@����ٿQ���m�@z����4@��
9�!?oe��{�@����ٿQ���m�@z����4@��
9�!?oe��{�@¶.���ٿ�Y�����@wUC�4@Y���!?�G�lҕ@¶.���ٿ�Y�����@wUC�4@Y���!?�G�lҕ@�����ٿDX����@uB���3@wg����!??WR���@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@�}f2�ٿ��,��@�����3@3|�"��!?��f	Q�@`M��Ԡٿ���N��@�b���4@��fLy�!?��[��h�@`M��Ԡٿ���N��@�b���4@��fLy�!?��[��h�@`M��Ԡٿ���N��@�b���4@��fLy�!?��[��h�@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�ʸ�F�ٿu���}��@�=�J!4@���BA�!?��^���@�%�ٿ�����@�`�,�4@=�>H�!?��A�3�@�%�ٿ�����@�`�,�4@=�>H�!?��A�3�@�%�ٿ�����@�`�,�4@=�>H�!?��A�3�@�%�ٿ�����@�`�,�4@=�>H�!?��A�3�@�%�ٿ�����@�`�,�4@=�>H�!?��A�3�@�����ٿ�4�6��@�?iD��3@D6� l�!?-��Ss�@	~�|�ٿQs/��@�s���"4@���'j�!?�|����@	~�|�ٿQs/��@�s���"4@���'j�!?�|����@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@C2f�ٿq*'Et�@Q.9L�"4@A^��u�!?���<"�@t�z�ٿW��g�@��y�6f4@�aGUv�!?���<�@���"-�ٿC �2�@�\@4@[�x@�!?����aa�@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@IS,��ٿS.�%A�@�m'�24@�d��!?Y`��@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@�/���ٿ��jr�@�����4@Q��m�!?/W`~ʕ@z�7�6�ٿ�lkB��@�^��4@S_�hj�!?6$;G��@z�7�6�ٿ�lkB��@�^��4@S_�hj�!?6$;G��@z�7�6�ٿ�lkB��@�^��4@S_�hj�!?6$;G��@z�7�6�ٿ�lkB��@�^��4@S_�hj�!?6$;G��@^�Нٿ�{X~Y��@�Wr��4@PXMd�!?V%=��@^�Нٿ�{X~Y��@�Wr��4@PXMd�!?V%=��@^�Нٿ�{X~Y��@�Wr��4@PXMd�!?V%=��@����A�ٿ�_��7�@aW��.4@�Zˏ��!?^�o�n��@����A�ٿ�_��7�@aW��.4@�Zˏ��!?^�o�n��@����A�ٿ�_��7�@aW��.4@�Zˏ��!?^�o�n��@����A�ٿ�_��7�@aW��.4@�Zˏ��!?^�o�n��@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@�� BХٿ�����@�~�Y�3@�s&b#�!?��UeMǕ@nq�Ǣٿ�ǟA'�@�����3@[.]�!?�ßP7�@nq�Ǣٿ�ǟA'�@�����3@[.]�!?�ßP7�@nq�Ǣٿ�ǟA'�@�����3@[.]�!?�ßP7�@��-fr�ٿ��`����@�,0��3@ÊZ�}�!?�oL���@��-fr�ٿ��`����@�,0��3@ÊZ�}�!?�oL���@��-fr�ٿ��`����@�,0��3@ÊZ�}�!?�oL���@��-fr�ٿ��`����@�,0��3@ÊZ�}�!?�oL���@B� �z�ٿ��;�@��Ly�3@�np�!?��*v�@�P�{.�ٿ�!M�9��@;��2��3@���А!?�c�}���@�P�{.�ٿ�!M�9��@;��2��3@���А!?�c�}���@汖=��ٿ������@c����3@��!2�!?~�	���@汖=��ٿ������@c����3@��!2�!?~�	���@汖=��ٿ������@c����3@��!2�!?~�	���@汖=��ٿ������@c����3@��!2�!?~�	���@汖=��ٿ������@c����3@��!2�!?~�	���@y\���ٿv5q���@���~%4@����!?T��'ƥ�@y\���ٿv5q���@���~%4@����!?T��'ƥ�@y\���ٿv5q���@���~%4@����!?T��'ƥ�@�F�9�ٿ���V��@����i|4@�	���!?{fs��:�@�F�9�ٿ���V��@����i|4@�	���!?{fs��:�@�F�9�ٿ���V��@����i|4@�	���!?{fs��:�@�F�9�ٿ���V��@����i|4@�	���!?{fs��:�@�XQ�1�ٿE\^}���@�+#��4@A����!?l��Ұ��@�XQ�1�ٿE\^}���@�+#��4@A����!?l��Ұ��@�XQ�1�ٿE\^}���@�+#��4@A����!?l��Ұ��@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@���h�ٿD��]�@�6J��I4@,$��4�!?��x�:'�@����ٿ8�)J?C�@!Sn6�@4@��$j`�!?<b��H�@����ٿ8�)J?C�@!Sn6�@4@��$j`�!?<b��H�@����ٿ8�)J?C�@!Sn6�@4@��$j`�!?<b��H�@����ٿ8�)J?C�@!Sn6�@4@��$j`�!?<b��H�@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@}��M�ٿ��X{��@� ��34@{n=�!?�q�ϕ@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@ӫ$�ٿ%��`L,�@[
 �4@RO�!?�����@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@��^D0�ٿE��篌�@B����3@�uef6�!?R�	(�a�@K����ٿ��YXI��@��X}��3@,��8�!?x#��6�@K����ٿ��YXI��@��X}��3@,��8�!?x#��6�@K����ٿ��YXI��@��X}��3@,��8�!?x#��6�@���\��ٿ���Ϛ��@�C#��3@�P8U�!?��c�6L�@���\��ٿ���Ϛ��@�C#��3@�P8U�!?��c�6L�@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@$�z�c�ٿ�T]Ţ�@��E���3@��>A�!?�P�n$��@R��1�ٿ��/]��@��Lv4@������!?,����r�@R��1�ٿ��/]��@��Lv4@������!?,����r�@{�y��ٿ$K�W�@�IA��4@P�~&�!?�N�Glݕ@{�y��ٿ$K�W�@�IA��4@P�~&�!?�N�Glݕ@{�y��ٿ$K�W�@�IA��4@P�~&�!?�N�Glݕ@{�y��ٿ$K�W�@�IA��4@P�~&�!?�N�Glݕ@�4~S�ٿ����"�@|��<�84@����E�!?e7C%�@�4~S�ٿ����"�@|��<�84@����E�!?e7C%�@�4~S�ٿ����"�@|��<�84@����E�!?e7C%�@�4~S�ٿ����"�@|��<�84@����E�!?e7C%�@a�x��ٿ{��P5��@��z� 4@%�qT�!?���7T�@a�x��ٿ{��P5��@��z� 4@%�qT�!?���7T�@a�x��ٿ{��P5��@��z� 4@%�qT�!?���7T�@a�x��ٿ{��P5��@��z� 4@%�qT�!?���7T�@a�x��ٿ{��P5��@��z� 4@%�qT�!?���7T�@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@���8�ٿv�Sp�R�@-�/4@�v}�r�!?�Z����@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@��fg��ٿ氪7���@��Դ��3@{݉�I�!?mz�W���@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@�rԐ�ٿ
zYj��@W�#VP4@��"E�!?+iٶ�U�@hPҒ��ٿs7P>C��@��r[k�3@�}��!?Lu�^:��@hPҒ��ٿs7P>C��@��r[k�3@�}��!?Lu�^:��@hPҒ��ٿs7P>C��@��r[k�3@�}��!?Lu�^:��@hPҒ��ٿs7P>C��@��r[k�3@�}��!?Lu�^:��@hPҒ��ٿs7P>C��@��r[k�3@�}��!?Lu�^:��@a��r�ٿ�pm`w��@6�X��3@'�<ɨ�!?�7��ҕ@a��r�ٿ�pm`w��@6�X��3@'�<ɨ�!?�7��ҕ@�Ie�˗ٿ�tS�4�@�V�/4@��"f�!?.�@)�@�Ie�˗ٿ�tS�4�@�V�/4@��"f�!?.�@)�@�Ie�˗ٿ�tS�4�@�V�/4@��"f�!?.�@)�@�Ie�˗ٿ�tS�4�@�V�/4@��"f�!?.�@)�@�Ie�˗ٿ�tS�4�@�V�/4@��"f�!?.�@)�@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@({����ٿ�l� ��@��])4@,�,A�!?N'�nߕ@{GdW7�ٿ� ޝ��@G;� 4@���I;�!?#��%4,�@{GdW7�ٿ� ޝ��@G;� 4@���I;�!?#��%4,�@{GdW7�ٿ� ޝ��@G;� 4@���I;�!?#��%4,�@��m�ٿ@J��5�@�T���3@�#@�l�!? ��7��@��m�ٿ@J��5�@�T���3@�#@�l�!? ��7��@��m�ٿ@J��5�@�T���3@�#@�l�!? ��7��@��56��ٿ]�?��@�eOϔ�3@9`�"�!?%@/cY"�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@<��ݟٿpA�?�t�@���}�3@"��2�!?\���0�@���e��ٿ����Ӽ�@r��"�3@-�>�!?Kc�;i�@���e��ٿ����Ӽ�@r��"�3@-�>�!?Kc�;i�@�L3��ٿ�^���<�@�2��4@�Fq��!?ľBG�t�@�����ٿ���6��@�B��B4@d�[�+�!?�x�@Y�@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@R$x�Ûٿd��TM�@s�u��-4@�0]�!?	�=�ŕ@�1�q��ٿ䲤�p�@)���w4@QB*ᗐ!?}���֕@�1�q��ٿ䲤�p�@)���w4@QB*ᗐ!?}���֕@�1�q��ٿ䲤�p�@)���w4@QB*ᗐ!?}���֕@�����ٿ%�P�@��OScO4@��6q�!?�K3K�a�@�����ٿ%�P�@��OScO4@��6q�!?�K3K�a�@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�6��ٿ��ݼ��@��.��h4@�~-�ؐ!?�����@�� �ٿͧ+%�@w-�'V4@ouϛ��!?��9)i�@�� �ٿͧ+%�@w-�'V4@ouϛ��!?��9)i�@j�,��ٿ�ZL���@��E�?4@�`Y.��!?�{� ��@j�,��ٿ�ZL���@��E�?4@�`Y.��!?�{� ��@j7[p֢ٿh�F��@��C�4@d-6��!?��t��@j7[p֢ٿh�F��@��C�4@d-6��!?��t��@�T�>�ٿ^q sۇ�@T���@4@��䮫�!?nu��@�T�>�ٿ^q sۇ�@T���@4@��䮫�!?nu��@���ٿE�7|��@5��K4@���IƐ!?�b��b�@���ٿE�7|��@5��K4@���IƐ!?�b��b�@���ٿE�7|��@5��K4@���IƐ!?�b��b�@���6s�ٿGס���@K;����3@�3���!?�礙X#�@���6s�ٿGס���@K;����3@�3���!?�礙X#�@���6s�ٿGס���@K;����3@�3���!?�礙X#�@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@� �ɐ�ٿ�.h�$��@�ߺ0��3@U����!?d/|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@9-!�ߤٿҗ �@�w��C4@�k��R�!?0��|��@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@����9�ٿt��5�@숼�dZ4@�R��;�!?��5�@)���ٿ�bu�o��@K�.L#:4@SȘ'�!?�yK<�Z�@)���ٿ�bu�o��@K�.L#:4@SȘ'�!?�yK<�Z�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@M�W�ٿ�����u�@dIn�G64@K�/��!?�k�)*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@L��{�ٿ��*�@�JؿH4@$
}�G�!?���;*�@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@�����ٿ��w���@^��z34@�W�g�!?K�����@󞀿p�ٿ\���2a�@�����4@���%K�!?��]����@}����ٿ �R��@��dtJ=4@%r��M�!?%�g��~�@}����ٿ �R��@��dtJ=4@%r��M�!?%�g��~�@V�r�W�ٿ�v�T��@v�1�x4@:z|]�!?�֍�M��@|u,���ٿ=o�!�g�@'00�4@�Ƚ�S�!?��M�`��@�4,��ٿf"���@Aݎ��l4@�$�"��!?���Q��@�4,��ٿf"���@Aݎ��l4@�$�"��!?���Q��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@����X�ٿ}���t��@=�F^_!4@e�Ʋ�!?`=�1��@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@y%	ǝٿu�SHb��@��vK94@{|���!?z3�����@�P�1H�ٿj�聯��@���&�4@1�'nÐ!?��`3�@�P�1H�ٿj�聯��@���&�4@1�'nÐ!?��`3�@�P�1H�ٿj�聯��@���&�4@1�'nÐ!?��`3�@�P�1H�ٿj�聯��@���&�4@1�'nÐ!?��`3�@�P�1H�ٿj�聯��@���&�4@1�'nÐ!?��`3�@�-&`�ٿ3M�C�@��	%4@��Զb�!?7���-��@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�s�8d�ٿ�~B윿�@��]hp4@�r�&o�!?������@�7�|B�ٿ�މ}|�@����|�3@���P�!?y.�ȡb�@�7�|B�ٿ�މ}|�@����|�3@���P�!?y.�ȡb�@�7�|B�ٿ�މ}|�@����|�3@���P�!?y.�ȡb�@�7�|B�ٿ�މ}|�@����|�3@���P�!?y.�ȡb�@m:��٣ٿ�meφ��@)!mI4@�Ĝ���!?k����ٕ@<p-�ƟٿWD�m���@��s�4@�Gv Ɛ!?֫��@<p-�ƟٿWD�m���@��s�4@�Gv Ɛ!?֫��@<p-�ƟٿWD�m���@��s�4@�Gv Ɛ!?֫��@E��!��ٿ�A����@����4@�$39o�!?��#���@E��!��ٿ�A����@����4@�$39o�!?��#���@E��!��ٿ�A����@����4@�$39o�!?��#���@��
%�ٿV��ƻ��@U���lQ4@JV�\�!?�]S'��@��
%�ٿV��ƻ��@U���lQ4@JV�\�!?�]S'��@��
%�ٿV��ƻ��@U���lQ4@JV�\�!?�]S'��@��
%�ٿV��ƻ��@U���lQ4@JV�\�!?�]S'��@��E>L�ٿ?�^���@�rv�B)4@X�&�e�!?�R�'�Ǖ@��E>L�ٿ?�^���@�rv�B)4@X�&�e�!?�R�'�Ǖ@��E>L�ٿ?�^���@�rv�B)4@X�&�e�!?�R�'�Ǖ@��E>L�ٿ?�^���@�rv�B)4@X�&�e�!?�R�'�Ǖ@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@?,y2��ٿP�x��@�a��3@i�Uk�!?�;N�ӡ�@�߶��ٿ�c���"�@�c����3@�j�'g�!?��k؜�@�߶��ٿ�c���"�@�c����3@�j�'g�!?��k؜�@�߶��ٿ�c���"�@�c����3@�j�'g�!?��k؜�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@��z��ٿ�U���Q�@����2&4@D�vz�!?�A$�K$�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@Hu��ٿ�8�ds��@��J>)4@:���!?�@*a�8�@���ٿ�6���j�@����34@"��8��!?Q��QO�@���ٿ�6���j�@����34@"��8��!?Q��QO�@���ٿ�6���j�@����34@"��8��!?Q��QO�@���ٿ�6���j�@����34@"��8��!?Q��QO�@���ٿ�6���j�@����34@"��8��!?Q��QO�@��_v�ٿ��̄��@`�!c��3@q%��s�!??�\@�@��_v�ٿ��̄��@`�!c��3@q%��s�!??�\@�@��H��ٿ����G��@��E��4@�Z�M��!?HJ�S�@��H��ٿ����G��@��E��4@�Z�M��!?HJ�S�@)=�-�ٿk�����@\p��4@���ژ�!?�
��D�@)=�-�ٿk�����@\p��4@���ژ�!?�
��D�@)=�-�ٿk�����@\p��4@���ژ�!?�
��D�@)=�-�ٿk�����@\p��4@���ژ�!?�
��D�@)=�-�ٿk�����@\p��4@���ژ�!?�
��D�@0�;�R�ٿwP�Q��@ߚ�K��3@����l�!?*;[澆�@0�;�R�ٿwP�Q��@ߚ�K��3@����l�!?*;[澆�@�����ٿ�'���/�@%�r"�3@Tq��~�!?ĳ���@�����ٿ�'���/�@%�r"�3@Tq��~�!?ĳ���@�����ٿ�'���/�@%�r"�3@Tq��~�!?ĳ���@�����ٿ�'���/�@%�r"�3@Tq��~�!?ĳ���@�����ٿ�'���/�@%�r"�3@Tq��~�!?ĳ���@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@���T�ٿ.G3����@f�^�2�3@w)���!?F��b�@%n���ٿ�Z���=�@0���3@H�}u�!?�
�?{��@%n���ٿ�Z���=�@0���3@H�}u�!?�
�?{��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@������ٿ�Ҽ��@�����3@v�ߨ��!?�G��@�����ٿ�N1Q��@>a�P�3@�����!?A��j"ʕ@�Fo�5�ٿ`�}"j��@�� �q4@��Л�!?l�/�	�@�Fo�5�ٿ`�}"j��@�� �q4@��Л�!?l�/�	�@�Fo�5�ٿ`�}"j��@�� �q4@��Л�!?l�/�	�@NT#��ٿ��%��@�+jjkE4@2V��:�!?Ot�Ȅӕ@NT#��ٿ��%��@�+jjkE4@2V��:�!?Ot�Ȅӕ@NT#��ٿ��%��@�+jjkE4@2V��:�!?Ot�Ȅӕ@NT#��ٿ��%��@�+jjkE4@2V��:�!?Ot�Ȅӕ@y����ٿ�vn�A �@�B3�B�3@5��B�!?r	[�w�@y����ٿ�vn�A �@�B3�B�3@5��B�!?r	[�w�@y����ٿ�vn�A �@�B3�B�3@5��B�!?r	[�w�@y����ٿ�vn�A �@�B3�B�3@5��B�!?r	[�w�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@�:���ٿk�_J ��@�S���%4@�hR�X�!?��E�݅�@0����ٿ���(��@a�
64@���l%�!?��U��@��Ÿ%�ٿ��`���@lqAؘF4@����!?n��I�@[C��ٿ݃�?֡�@:��"S4@Qe���!?�_<-�@?�
}�ٿ��<�@d����h4@Ⱥ:�Y�!?>�ݫe�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@�Õf�ٿ>}�X'*�@�H��e.4@h��V�!?QlV:r�@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@$�;��ٿ�Tl�e�@g��Mq&4@a��J�!?�f�ە@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@_-����ٿm�"�.�@��=4@����!?�ڬM=�@s�R~��ٿ�v��Ab�@��߆b4@���8��!?� ��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@�ja�ٿژ� ���@�����74@���8��!?��!��@c�r�ٿ���?��@#�0<\4@?Xc�u�!?�ժ'$ݕ@��j<�ٿA�f����@���r�$4@�^@�!?�V_���@��j<�ٿA�f����@���r�$4@�^@�!?�V_���@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�����ٿ�����@��#Y4@�ZP�!?'�)�.��@�3��ٿ��t��@��j;54@�A��|�!?o,���@F7,K�ٿ�O��1�@����04@�Ѳf�!?�P<}�o�@F7,K�ٿ�O��1�@����04@�Ѳf�!?�P<}�o�@F7,K�ٿ�O��1�@����04@�Ѳf�!?�P<}�o�@F7,K�ٿ�O��1�@����04@�Ѳf�!?�P<}�o�@F7,K�ٿ�O��1�@����04@�Ѳf�!?�P<}�o�@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@G�2a�ٿ��&����@Ǖ&��4@�MĠ�!?�n=���@�&���ٿ�/Y�@&<��4@����z�!?�į!���@�&���ٿ�/Y�@&<��4@����z�!?�į!���@�����ٿ�m�N{��@��!��M4@\Y=읐!?��	f��@�����ٿ�m�N{��@��!��M4@\Y=읐!?��	f��@�����ٿ�m�N{��@��!��M4@\Y=읐!?��	f��@�����ٿ�m�N{��@��!��M4@\Y=읐!?��	f��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@? �҇�ٿ����@��W4@(#bd<�!?%�d�n��@��ebѢٿ6.�X^y�@�	��?4@&�P�E�!?Y���R��@��ebѢٿ6.�X^y�@�	��?4@&�P�E�!?Y���R��@��ebѢٿ6.�X^y�@�	��?4@&�P�E�!?Y���R��@~�m ��ٿj�n?�l�@��$�(4@���&�!?��/?底@~�m ��ٿj�n?�l�@��$�(4@���&�!?��/?底@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@�����ٿ���͐��@��]u��3@�.O��!?�ڻЕ@eDq��ٿ/�8=��@�J�.�;4@u�-�!?iDA�@eDq��ٿ/�8=��@�J�.�;4@u�-�!?iDA�@eDq��ٿ/�8=��@�J�.�;4@u�-�!?iDA�@eDq��ٿ/�8=��@�J�.�;4@u�-�!?iDA�@eDq��ٿ/�8=��@�J�.�;4@u�-�!?iDA�@᫸���ٿ�Dj�@~�s��4@<�o�!?1��GU��@᫸���ٿ�Dj�@~�s��4@<�o�!?1��GU��@᫸���ٿ�Dj�@~�s��4@<�o�!?1��GU��@᫸���ٿ�Dj�@~�s��4@<�o�!?1��GU��@᫸���ٿ�Dj�@~�s��4@<�o�!?1��GU��@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@��l���ٿ}��!0��@��y�+4@��\�!?\�m���@�"���ٿ����}�@篜�4@S��R�!?}��*l�@�"���ٿ����}�@篜�4@S��R�!?}��*l�@�"���ٿ����}�@篜�4@S��R�!?}��*l�@�"���ٿ����}�@篜�4@S��R�!?}��*l�@�"���ٿ����}�@篜�4@S��R�!?}��*l�@�"���ٿ����}�@篜�4@S��R�!?}��*l�@���h�ٿ���j�@�d�4@��c�!?��R��J�@���h�ٿ���j�@�d�4@��c�!?��R��J�@���h�ٿ���j�@�d�4@��c�!?��R��J�@���h�ٿ���j�@�d�4@��c�!?��R��J�@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@�~ 餡ٿ��ku7�@�B���3@+�SN�!?�[�����@ �f��ٿ�{B���@�-�&#�3@صA�]�!?�}R�ƕ@ �f��ٿ�{B���@�-�&#�3@صA�]�!?�}R�ƕ@ �f��ٿ�{B���@�-�&#�3@صA�]�!?�}R�ƕ@ �f��ٿ�{B���@�-�&#�3@صA�]�!?�}R�ƕ@ �f��ٿ�{B���@�-�&#�3@صA�]�!?�}R�ƕ@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@*�#=��ٿ`E;��_�@���t�3@�߇0}�!?j%�߱�@�IƘ�ٿqGL���@��RV4@o��dJ�!?���7˒�@�IƘ�ٿqGL���@��RV4@o��dJ�!?���7˒�@�IƘ�ٿqGL���@��RV4@o��dJ�!?���7˒�@����ٿ��{P�M�@�����3@8��w�!?������@����ٿ��{P�M�@�����3@8��w�!?������@����ٿ��{P�M�@�����3@8��w�!?������@���(�ٿKw����@w��Y�4@?P�|�!?��s��@���(�ٿKw����@w��Y�4@?P�|�!?��s��@���(�ٿKw����@w��Y�4@?P�|�!?��s��@��c��ٿ�E�2Y|�@��=��-4@ĖBC�!?$��|�ٕ@��c��ٿ�E�2Y|�@��=��-4@ĖBC�!?$��|�ٕ@>S#ə�ٿ�C.{���@Q0 �4@�\>=i�!?3�WA���@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@vpA��ٿ4S�m��@��{���3@�z�5�!?�h��)9�@j�۟r�ٿ��G���@xt�.�3@Wߣ�J�!?���L���@�r��Ϣٿ�2E����@��5�3@���O�!?��u���@P~�,D�ٿyc	w�I�@����3@KՅ��!?�u?�@s4�A��ٿ���Ζ�@&1��4@�'r��!?p�D&C�@�4��ٿ�$a���@ϖ����3@��Ne��!?��8،��@�4��ٿ�$a���@ϖ����3@��Ne��!?��8،��@�4��ٿ�$a���@ϖ����3@��Ne��!?��8،��@�4��ٿ�$a���@ϖ����3@��Ne��!?��8،��@?m����ٿ�0���@�{����3@���!?\���@?m����ٿ�0���@�{����3@���!?\���@��٩9�ٿ�(K�0��@4ԙI4@m0���!?��E���@�r��ٿS��x�@�����<4@#�����!?Bf����@o,���ٿQ?f��@S��/5$4@�;.箐!?\?R���@o,���ٿQ?f��@S��/5$4@�;.箐!?\?R���@o,���ٿQ?f��@S��/5$4@�;.箐!?\?R���@o,���ٿQ?f��@S��/5$4@�;.箐!?\?R���@Uۤh��ٿ
R����@l�T��3@o�Ҕ�!?���;
�@Uۤh��ٿ
R����@l�T��3@o�Ҕ�!?���;
�@<����ٿyr*cY��@� ����3@�1���!?���
��@<����ٿyr*cY��@� ����3@�1���!?���
��@<����ٿyr*cY��@� ����3@�1���!?���
��@<����ٿyr*cY��@� ����3@�1���!?���
��@<����ٿyr*cY��@� ����3@�1���!?���
��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�.,ڛٿ�1�Yݞ�@h�4z��3@��EMe�!?G�9��@�"���ٿm>Py�@tújb�3@,N�Ce�!?&�:��@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@�5��ٿ#�OsL<�@d�]��3@�g��J�!?/ ]U�@����ٿ��(~a�@�i��G4@#q��D�!?��2��@����ٿ��(~a�@�i��G4@#q��D�!?��2��@N4��ٿEe��E��@Vx�c4@����!?�|?�z��@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@�2u�ٿ.2�J4�@���o�44@!3��!?_�d5먕@A��ɘٿ��a%Zr�@���&4@�wV�܏!?r+xӿ�@���N�ٿ?vә�@�����	4@�����!?I����@���N�ٿ?vә�@�����	4@�����!?I����@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@h��h�ٿ��f%p�@�IZ�4@���cO�!?��vC�N�@�����ٿ�E�3��@VA�s�3@�Hf�!?��.@Z�@�����ٿ�E�3��@VA�s�3@�Hf�!?��.@Z�@,l�C��ٿ�3��(��@�>Q�M4@h�7[N�!?�\�Pn�@,l�C��ٿ�3��(��@�>Q�M4@h�7[N�!?�\�Pn�@,l�C��ٿ�3��(��@�>Q�M4@h�7[N�!?�\�Pn�@ �"���ٿ���c"�@�����34@)���A�!?\���ʨ�@ �"���ٿ���c"�@�����34@)���A�!?\���ʨ�@ �"���ٿ���c"�@�����34@)���A�!?\���ʨ�@ �"���ٿ���c"�@�����34@)���A�!?\���ʨ�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@5K�E�ٿL�Q/��@bp��U4@���w@�!?�:�-�Y�@j�f���ٿ��T4	�@��u�G4@�'W�}�!?\��X�@j�f���ٿ��T4	�@��u�G4@�'W�}�!?\��X�@j�f���ٿ��T4	�@��u�G4@�'W�}�!?\��X�@��h�ٿ��CY��@�����@4@}?�zh�!?0d�S�a�@��h�ٿ��CY��@�����@4@}?�zh�!?0d�S�a�@��h�ٿ��CY��@�����@4@}?�zh�!?0d�S�a�@0t�ٿ�*����@�iG!h�3@���O�!?�ێʵ%�@0t�ٿ�*����@�iG!h�3@���O�!?�ێʵ%�@0t�ٿ�*����@�iG!h�3@���O�!?�ێʵ%�@0t�ٿ�*����@�iG!h�3@���O�!?�ێʵ%�@��J��ٿy��o��@�;�q~�3@G�w��!?�m�0n��@D�<;��ٿ �9�@;L�s��3@�x>52�!?�x���@e��1O�ٿ���V�z�@����z!4@����6�!?]�ҕ@e��1O�ٿ���V�z�@����z!4@����6�!?]�ҕ@e��1O�ٿ���V�z�@����z!4@����6�!?]�ҕ@e��1O�ٿ���V�z�@����z!4@����6�!?]�ҕ@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@�)Ǡٿ��-�@��I�L4@����9�!?�5g�|{�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@ް�=ޚٿl%�a�A�@SAN��)4@^j�3W�!?�T�@�j�@J���ٿ��I�O�@��T�N�3@���ܜ�!?%��ȕ@J���ٿ��I�O�@��T�N�3@���ܜ�!?%��ȕ@�:�ٗٿ���Mv�@%M���	4@���dr�!?Pi�p��@�:�ٗٿ���Mv�@%M���	4@���dr�!?Pi�p��@�:�ٗٿ���Mv�@%M���	4@���dr�!?Pi�p��@ݍ�}�ٿ���`�@P��ܕ'4@�ܮ���!?<:Q�ٕ@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@zq��ڡٿ'u+�4�@�v�n4@���LL�!?�b����@�鎳�ٿ������@Up((� 4@E� V�!?��,j��@�鎳�ٿ������@Up((� 4@E� V�!?��,j��@�鎳�ٿ������@Up((� 4@E� V�!?��,j��@�鎳�ٿ������@Up((� 4@E� V�!?��,j��@$�4�ٿ7�^:o?�@#S�J4@����N�!?���y6�@$�4�ٿ7�^:o?�@#S�J4@����N�!?���y6�@hu�Ə�ٿ�in;��@�����|4@V�7q�!?w��Y�K�@hu�Ə�ٿ�in;��@�����|4@V�7q�!?w��Y�K�@hu�Ə�ٿ�in;��@�����|4@V�7q�!?w��Y�K�@hu�Ə�ٿ�in;��@�����|4@V�7q�!?w��Y�K�@hu�Ə�ٿ�in;��@�����|4@V�7q�!?w��Y�K�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@�H��ɚٿ�O:fB�@!��Ŷ�4@sXzY�!?�HAtI5�@=��%��ٿ#qG���@�%Y�Xe4@<� ��!?���8�@=��%��ٿ#qG���@�%Y�Xe4@<� ��!?���8�@�Wn��ٿ������@'y@y�A4@�	��!?��;!�@�Wn��ٿ������@'y@y�A4@�	��!?��;!�@�Wn��ٿ������@'y@y�A4@�	��!?��;!�@�Wn��ٿ������@'y@y�A4@�	��!?��;!�@�Wn��ٿ������@'y@y�A4@�	��!?��;!�@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@_�.h�ٿ K �$�@���^�A4@��A��!?�`�@���@�xb�d�ٿ)�m �w�@�<L�4@���<�!?|�)����@�xb�d�ٿ)�m �w�@�<L�4@���<�!?|�)����@�xb�d�ٿ)�m �w�@�<L�4@���<�!?|�)����@�xb�d�ٿ)�m �w�@�<L�4@���<�!?|�)����@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@c4R�x�ٿ:��O��@3Koe�3@�&�jJ�!?(N$�`��@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�H�:��ٿW��k��@��}U�>4@r�(z�!?��t	ŀ�@�KyT]�ٿ3���V��@I�674@� ���!?隸�L��@�KyT]�ٿ3���V��@I�674@� ���!?隸�L��@�KyT]�ٿ3���V��@I�674@� ���!?隸�L��@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@}[dR�ٿ�����@rV
!w�3@���'�!?{�:(�ޕ@h�QGz�ٿ�b�)Go�@X���4@�P	�!?��o<Օ@h�QGz�ٿ�b�)Go�@X���4@�P	�!?��o<Օ@h�QGz�ٿ�b�)Go�@X���4@�P	�!?��o<Օ@h�QGz�ٿ�b�)Go�@X���4@�P	�!?��o<Օ@�}^,�ٿܥ�S���@L1��x?4@�|��!?]��9�z�@�}^,�ٿܥ�S���@L1��x?4@�|��!?]��9�z�@�}^,�ٿܥ�S���@L1��x?4@�|��!?]��9�z�@�}^,�ٿܥ�S���@L1��x?4@�|��!?]��9�z�@�}^,�ٿܥ�S���@L1��x?4@�|��!?]��9�z�@�I��l�ٿ�&6�}�@����"_4@�v�rq�!?�P���@�I��l�ٿ�&6�}�@����"_4@�v�rq�!?�P���@�Htt��ٿ_pH����@�<�nn/4@���!?E���@�Htt��ٿ_pH����@�<�nn/4@���!?E���@�^S���ٿ�uGd`�@�I��?4@�ʽ��!?��]���@�^S���ٿ�uGd`�@�I��?4@�ʽ��!?��]���@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@:.�K�ٿ�ԕ����@��9�n�3@\.�u�!?���߀��@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@뺝y��ٿ��w&�@�=AU�3@?���K�!?%�>�c�@�5��ٿaށ�X�@Q�j�4@ՙC8b�!?�JT�@��U
ɡٿ.��`0�@!��) 4@v�J�U�!?��H�cx�@��U
ɡٿ.��`0�@!��) 4@v�J�U�!?��H�cx�@��U
ɡٿ.��`0�@!��) 4@v�J�U�!?��H�cx�@��U
ɡٿ.��`0�@!��) 4@v�J�U�!?��H�cx�@��U
ɡٿ.��`0�@!��) 4@v�J�U�!?��H�cx�@OM���ٿ�w$
W�@!�B�X%4@l�$d�!?�*̸e�@OM���ٿ�w$
W�@!�B�X%4@l�$d�!?�*̸e�@OM���ٿ�w$
W�@!�B�X%4@l�$d�!?�*̸e�@OM���ٿ�w$
W�@!�B�X%4@l�$d�!?�*̸e�@���\I�ٿ�,��z�@؈#�54@���)��!?4��&���@�MF}�ٿs�4�P��@�8��[4@o�Vsy�!?Νļ��@�MF}�ٿs�4�P��@�8��[4@o�Vsy�!?Νļ��@�MF}�ٿs�4�P��@�8��[4@o�Vsy�!?Νļ��@�MF}�ٿs�4�P��@�8��[4@o�Vsy�!?Νļ��@�D����ٿ@�08_��@@7�AP4@�2�r
�!?4� P��@�D����ٿ@�08_��@@7�AP4@�2�r
�!?4� P��@�D����ٿ@�08_��@@7�AP4@�2�r
�!?4� P��@�D����ٿ@�08_��@@7�AP4@�2�r
�!?4� P��@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@w��}�ٿ|%M<\�@�Yt�&4@?{��!?x����@�wK>��ٿ� -��@]��d�4@Q��NL�!?�x�}��@�wK>��ٿ� -��@]��d�4@Q��NL�!?�x�}��@Q��-��ٿL	��9�@��u&4@�Qw1?�!?�����@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@�atݘٿ l�n���@N�/�54@�l.��!?�����ٕ@7�YG�ٿ;.tF���@gcߤoJ4@6p�!?y��Ė̕@7�YG�ٿ;.tF���@gcߤoJ4@6p�!?y��Ė̕@7�YG�ٿ;.tF���@gcߤoJ4@6p�!?y��Ė̕@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@��>Q�ٿjIh[��@�� ��04@j
�[�!?�އ��@�N�ٿ�r+���@�2�J;4@罰u�!?�Ѻ�o�@�N�ٿ�r+���@�2�J;4@罰u�!?�Ѻ�o�@�N�ٿ�r+���@�2�J;4@罰u�!?�Ѻ�o�@s�==M�ٿ�AX00��@�]�/4@�wL��!?i4��%�@s�==M�ٿ�AX00��@�]�/4@�wL��!?i4��%�@sX$�e�ٿd8A3��@�0�s4@�n��א!?��H��"�@sX$�e�ٿd8A3��@�0�s4@�n��א!?��H��"�@sX$�e�ٿd8A3��@�0�s4@�n��א!?��H��"�@sX$�e�ٿd8A3��@�0�s4@�n��א!?��H��"�@�yk���ٿ��7���@�9��<4@,l%]�!?ʕ�rTЕ@�yk���ٿ��7���@�9��<4@,l%]�!?ʕ�rTЕ@�yk���ٿ��7���@�9��<4@,l%]�!?ʕ�rTЕ@�yk���ٿ��7���@�9��<4@,l%]�!?ʕ�rTЕ@�yk���ٿ��7���@�9��<4@,l%]�!?ʕ�rTЕ@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@�����ٿ>����@�(1�y�3@a?{�!?��-"�@��Şٿ}V�t&�@k�f��3@+b�@m�!?����@��Şٿ}V�t&�@k�f��3@+b�@m�!?����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@&���R�ٿ���k��@��g���3@�ƻg�!?�����@��Չv�ٿ�'�b��@����3@�G�A��!?����ڕ@�n�,H�ٿ�sTh���@m�E�a�3@�}�q�!?�~fp��@���T�ٿ��r�@�Z�y��3@8�8O�!?�JLm@�@���T�ٿ��r�@�Z�y��3@8�8O�!?�JLm@�@�=v>y�ٿ
� ����@b�I��3@y��T�!?~��t�@:�#\�ٿ&op|�f�@Yu����3@S���C�!?5��Җ@�L�X�ٿ��4�sU�@���Hs�3@z87S=�!?	|��� �@�L�X�ٿ��4�sU�@���Hs�3@z87S=�!?	|��� �@�L�X�ٿ��4�sU�@���Hs�3@z87S=�!?	|��� �@�L�X�ٿ��4�sU�@���Hs�3@z87S=�!?	|��� �@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@������ٿ���a��@�(��q:4@c��N�!?����9�@sm��4�ٿ��fL��@5ɍ
�`4@Z�@s�!?Z��▕@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@'�x3�ٿK\wP�{�@ε/��%4@c�<��!?C�oD�@f��@��ٿA�Z�8�@��!u�D4@E"�Tn�!?��ʕ@f��@��ٿA�Z�8�@��!u�D4@E"�Tn�!?��ʕ@#� �c�ٿv׊brf�@�y�1j4@��� ��!?�%-���@#� �c�ٿv׊brf�@�y�1j4@��� ��!?�%-���@#� �c�ٿv׊brf�@�y�1j4@��� ��!?�%-���@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@NI�1֜ٿ��<4���@E��HX24@���ː!?:�&�@5�m/�ٿ_���$�@:-v4@����ɐ!?>k���M�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@�yk��ٿ�	��ch�@Eť5�D4@��"	А!?[��>�@���U˘ٿ%\�p�@T�	��P4@v�&��!?�v�	)@Ғ+5�ٿh�?��@w�H�f4@-B���!?�ƽ�5��@L~�	՝ٿ]ꂇ�l�@�I�G>S4@X�R�!?�֏Bu�@L~�	՝ٿ]ꂇ�l�@�I�G>S4@X�R�!?�֏Bu�@L~�	՝ٿ]ꂇ�l�@�I�G>S4@X�R�!?�֏Bu�@L~�	՝ٿ]ꂇ�l�@�I�G>S4@X�R�!?�֏Bu�@W�ĔјٿցKv��@�4@���!?�u�!ە@W�ĔјٿցKv��@�4@���!?�u�!ە@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@����ٿ#�>���@�#��/4@�Կ���!?@�C��p�@���D�ٿ�M� چ�@��ҧ��3@T5��!?�6��P�@���D�ٿ�M� چ�@��ҧ��3@T5��!?�6��P�@���D�ٿ�M� چ�@��ҧ��3@T5��!?�6��P�@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@�&N�ٿ��AE6�@~�+{	4@��O|�!?��bm���@R�g���ٿ��~�A�@7���3@*���!?�S�SǕ@R�g���ٿ��~�A�@7���3@*���!?�S�SǕ@R�g���ٿ��~�A�@7���3@*���!?�S�SǕ@R�g���ٿ��~�A�@7���3@*���!?�S�SǕ@(A�ʚٿ}����@�,��b�3@��/%��!?B ����@(A�ʚٿ}����@�,��b�3@��/%��!?B ����@(A�ʚٿ}����@�,��b�3@��/%��!?B ����@(A�ʚٿ}����@�,��b�3@��/%��!?B ����@a����ٿ�G����@��&�[�3@�퉡��!?A1{pӕ@a����ٿ�G����@��&�[�3@�퉡��!?A1{pӕ@a����ٿ�G����@��&�[�3@�퉡��!?A1{pӕ@��Ōߠٿς
�V��@��o9��3@4️�!?W�{ұ��@��Ōߠٿς
�V��@��o9��3@4️�!?W�{ұ��@��Ōߠٿς
�V��@��o9��3@4️�!?W�{ұ��@pjZ�ۙٿ$M�5��@Ⱦw�3@����!?܀�{$ܕ@pjZ�ۙٿ$M�5��@Ⱦw�3@����!?܀�{$ܕ@pjZ�ۙٿ$M�5��@Ⱦw�3@����!?܀�{$ܕ@�"7r.�ٿ������@��Z4@��_�!?*�Rm�+�@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@o�R��ٿ/�,n��@�l]���3@k���!?��/)��@��b;ܘٿ��>z�@,���4@0R��!?�o6rp��@��b;ܘٿ��>z�@,���4@0R��!?�o6rp��@Ʃ��T�ٿX0�p�d�@��W��(4@���!?�26����@Ʃ��T�ٿX0�p�d�@��W��(4@���!?�26����@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@(V�@W�ٿ[��
D��@����ڬ3@>>x%�!?�"y�3��@�7,���ٿ��H��P�@�V�,�3@��V�W�!?�ab��V�@�7,���ٿ��H��P�@�V�,�3@��V�W�!?�ab��V�@�7,���ٿ��H��P�@�V�,�3@��V�W�!?�ab��V�@�7,���ٿ��H��P�@�V�,�3@��V�W�!?�ab��V�@�L?sS�ٿ*�/�>��@/_<�4@0�Ag��!?��kZX�@�L?sS�ٿ*�/�>��@/_<�4@0�Ag��!?��kZX�@gH�[�ٿ}�����@���4@�}��!?�hŀŕ@gH�[�ٿ}�����@���4@�}��!?�hŀŕ@�@���ٿ�8�d���@�H�V44@�<'�4�!?�g2����@�@���ٿ�8�d���@�H�V44@�<'�4�!?�g2����@�@���ٿ�8�d���@�H�V44@�<'�4�!?�g2����@�@���ٿ�8�d���@�H�V44@�<'�4�!?�g2����@����ٿ��h���@�̜Du4@d\; ��!?u��ؕ@eF`���ٿ�g;��@L0�K�4@g��q�!?�JJ*�@eF`���ٿ�g;��@L0�K�4@g��q�!?�JJ*�@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@b����ٿ8��d[-�@����2#4@y��9��!?�>څ��@�u�H��ٿ��̌=g�@G�Q��4@T@�1v�!?���ځ�@�u�H��ٿ��̌=g�@G�Q��4@T@�1v�!?���ځ�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@I���0�ٿ3��$h��@Iך0�3@\E1ܐ!?�sT;�h�@fz��ѝٿ��k�R�@P��$�4@F���!?��ȑCM�@fz��ѝٿ��k�R�@P��$�4@F���!?��ȑCM�@fz��ѝٿ��k�R�@P��$�4@F���!?��ȑCM�@?U���ٿ�����@˙)$;04@k���Ð!?��ۑ���@?U���ٿ�����@˙)$;04@k���Ð!?��ۑ���@?U���ٿ�����@˙)$;04@k���Ð!?��ۑ���@drԘ�ٿ���^���@8��FS%4@ꄑ��!?��;�@drԘ�ٿ���^���@8��FS%4@ꄑ��!?��;�@D���ٿԡ�u���@����4�3@����!?�%M�@D���ٿԡ�u���@����4�3@����!?�%M�@d�d�ƛٿSЂq6��@]| f=�3@G���Ə!? �XLu/�@d�d�ƛٿSЂq6��@]| f=�3@G���Ə!? �XLu/�@�؈�ٿ`��z��@�	7o�3@����ޏ!?2奄��@�؈�ٿ`��z��@�	7o�3@����ޏ!?2奄��@�؈�ٿ`��z��@�	7o�3@����ޏ!?2奄��@�؈�ٿ`��z��@�	7o�3@����ޏ!?2奄��@�4��ٿ̈o&�@dI"	4@��?δ�!?G�5�ܕ@����ٿ'��)��@��ݤ��3@�F�s�!?�L�W���@����ٿ'��)��@��ݤ��3@�F�s�!?�L�W���@�~� ��ٿAwy��@�'��#4@Ns�S�!?���Ne�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@�ZA\�ٿ�}�:�@��=�644@�z��!?�Ui8�x�@��	hG�ٿ���U��@��Y4@o*T��!?|f�p��@��	hG�ٿ���U��@��Y4@o*T��!?|f�p��@�0�ᰝٿ�^D���@i~&�4@'��$k�!?�2i4餖@�0�ᰝٿ�^D���@i~&�4@'��$k�!?�2i4餖@�0�ᰝٿ�^D���@i~&�4@'��$k�!?�2i4餖@��YΞ�ٿ��v�_8�@[�Wb��3@���T�!?GZQV5ԕ@��YΞ�ٿ��v�_8�@[�Wb��3@���T�!?GZQV5ԕ@��YΞ�ٿ��v�_8�@[�Wb��3@���T�!?GZQV5ԕ@��YΞ�ٿ��v�_8�@[�Wb��3@���T�!?GZQV5ԕ@����ٿ��Sײ��@�TmAV4@��O���!?" �pZ�@����ٿ��Sײ��@�TmAV4@��O���!?" �pZ�@����ٿ��Sײ��@�TmAV4@��O���!?" �pZ�@����ٿ��Sײ��@�TmAV4@��O���!?" �pZ�@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@��{+�ٿ���Ǡ��@�;A�|04@!��cL�!?3�X���@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@�@��ٿ�1 #Ժ�@_���4@��9F�!?	3���v�@qWe1�ٿ𢭂9��@?Г�4@�H�>ڏ!?[�ѻi��@qWe1�ٿ𢭂9��@?Г�4@�H�>ڏ!?[�ѻi��@qWe1�ٿ𢭂9��@?Г�4@�H�>ڏ!?[�ѻi��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@mqⱖ�ٿ��N��@��F��4@Z[�n�!?��
��@ד�y�ٿ�UXp��@փ��B4@?�m�%�!?= D�]�@ד�y�ٿ�UXp��@փ��B4@?�m�%�!?= D�]�@ד�y�ٿ�UXp��@փ��B4@?�m�%�!?= D�]�@��r���ٿM.�a�@52�"4@֛<�!?��.z0�@��r���ٿM.�a�@52�"4@֛<�!?��.z0�@��r���ٿM.�a�@52�"4@֛<�!?��.z0�@��r���ٿM.�a�@52�"4@֛<�!?��.z0�@��r���ٿM.�a�@52�"4@֛<�!?��.z0�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�-��A�ٿҢB�R�@�6�+4@�hX�!?7��ۖp�@�P!̈́�ٿ7��{��@yY�<\4@�#S9�!?ab g��@�P!̈́�ٿ7��{��@yY�<\4@�#S9�!?ab g��@�P!̈́�ٿ7��{��@yY�<\4@�#S9�!?ab g��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@9V����ٿpc�x��@����4@=Z����!?���s��@�`:2�ٿ�T��Q��@�{޴��3@ƅ��؏!?́�v�ҕ@�`:2�ٿ�T��Q��@�{޴��3@ƅ��؏!?́�v�ҕ@�`:2�ٿ�T��Q��@�{޴��3@ƅ��؏!?́�v�ҕ@�`:2�ٿ�T��Q��@�{޴��3@ƅ��؏!?́�v�ҕ@������ٿE:�M�K�@�F�̜4@%Q�!?��+�^�@������ٿE:�M�K�@�F�̜4@%Q�!?��+�^�@������ٿE:�M�K�@�F�̜4@%Q�!?��+�^�@������ٿE:�M�K�@�F�̜4@%Q�!?��+�^�@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�63�~�ٿ}\i$Q�@C���'4@��e[�!?	!h=���@�}ŷ�ٿ�85j�@�e�j�4@����]�!?�l�LvC�@�}ŷ�ٿ�85j�@�e�j�4@����]�!?�l�LvC�@��Z�ٿ�񚸊C�@)�6�"4@'�o��!?��P���@��Z�ٿ�񚸊C�@)�6�"4@'�o��!?��P���@��Z�ٿ�񚸊C�@)�6�"4@'�o��!?��P���@B����ٿ�Z��V�@"�����3@;���a�!?DfΕ@B����ٿ�Z��V�@"�����3@;���a�!?DfΕ@��_�H�ٿmQ5����@�O��N 4@k�Ԅ��!? �Q���@��_�H�ٿmQ5����@�O��N 4@k�Ԅ��!? �Q���@��_�H�ٿmQ5����@�O��N 4@k�Ԅ��!? �Q���@��_�H�ٿmQ5����@�O��N 4@k�Ԅ��!? �Q���@j�T��ٿN�M�T��@^M�0�04@(.���!?
o�$�@ab[T�ٿ��p��{�@Lδg�+4@D/�^b�!?��.�B4�@�95�ٿ�_�jy�@�fr
s4@@�ȔD�!?\��v���@�95�ٿ�_�jy�@�fr
s4@@�ȔD�!?\��v���@�95�ٿ�_�jy�@�fr
s4@@�ȔD�!?\��v���@ڔG��ٿ]��ˢ�@M�w�&4@�>��J�!?4
t޵��@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@�/*���ٿC�����@�渂�4@�̔���!?"��ڻ�@w54R�ٿ]�N0�@��gNX4@�x����!?_6tM�b�@/���Y�ٿ��Z��@?Ȼ�k�3@W��Zr�!?̪��!Е@/���Y�ٿ��Z��@?Ȼ�k�3@W��Zr�!?̪��!Е@/���Y�ٿ��Z��@?Ȼ�k�3@W��Zr�!?̪��!Е@9W7@Ŗٿ7�M��@(��`4@�R_6ː!?m4�n%�@9W7@Ŗٿ7�M��@(��`4@�R_6ː!?m4�n%�@9W7@Ŗٿ7�M��@(��`4@�R_6ː!?m4�n%�@9W7@Ŗٿ7�M��@(��`4@�R_6ː!?m4�n%�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@��3vǛٿ�!�����@��3�3@�s�ǐ!?�M7�,a�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@7Anl��ٿ+���@�K���3@�"�QҐ!?��>tb�@P9�+5�ٿ�r���@ ��C4@OJw#��!?h2)})��@x1$�ٿ��ߞ��@�͟�R4@�*u�֐!?0L{F?r�@x1$�ٿ��ߞ��@�͟�R4@�*u�֐!?0L{F?r�@x1$�ٿ��ߞ��@�͟�R4@�*u�֐!?0L{F?r�@[2�kt�ٿ[�Qgw��@���:R4@� �?��!?[��%��@[2�kt�ٿ[�Qgw��@���:R4@� �?��!?[��%��@[2�kt�ٿ[�Qgw��@���:R4@� �?��!?[��%��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@:[�$�ٿ�r#ɕ�@��="�54@w�N��!?&�(8K��@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@�6��ٿ�����@��lё-4@�>PL�!?�kR����@un�ߙٿL�s�@�м%��3@���*�!?['1*���@4;3q�ٿ�hf����@��(�!4@�/���!?�խmnЕ@4;3q�ٿ�hf����@��(�!4@�/���!?�խmnЕ@4;3q�ٿ�hf����@��(�!4@�/���!?�խmnЕ@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@���ٿ��i�)F�@kax�74@�u2A�!?��U����@@}�
l�ٿ��Rn�@m%�m4@�U:W��!?�V�+��@@}�
l�ٿ��Rn�@m%�m4@�U:W��!?�V�+��@������ٿd�*��G�@;}�V�4@,���!?��͎@�@������ٿd�*��G�@;}�V�4@,���!?��͎@�@������ٿd�*��G�@;}�V�4@,���!?��͎@�@������ٿd�*��G�@;}�V�4@,���!?��͎@�@������ٿd�*��G�@;}�V�4@,���!?��͎@�@ʋ��S�ٿ�1Ad��@,_{\�3@�~^ꌐ!?��A��5�@ʋ��S�ٿ�1Ad��@,_{\�3@�~^ꌐ!?��A��5�@��P���ٿ�H��B�@QlV��3@���3�!?@.�p�@��P���ٿ�H��B�@QlV��3@���3�!?@.�p�@��P���ٿ�H��B�@QlV��3@���3�!?@.�p�@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@Hp����ٿ�ݫ�Vx�@�,�Gu�3@tm�} �!?�sR����@�d�ܡٿ$&�次�@X-���3@��k*�!?�����ە@�d�ܡٿ$&�次�@X-���3@��k*�!?�����ە@�d�ܡٿ$&�次�@X-���3@��k*�!?�����ە@�d�ܡٿ$&�次�@X-���3@��k*�!?�����ە@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@և`[ޝٿ�r���@5�����3@a#��!?X�teq��@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@lL�?ԗٿ����@�Bt���3@&z~�!?{+��D�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@3R�U+�ٿs��Eh
�@�B/�3@)/h�	�!?��#�'�@�"���ٿK�?3j��@�Hg���3@rZ}:�!?�z[��T�@�n;ha�ٿOӄ��@q��ò�3@!�&�l�!?p���U(�@�n;ha�ٿOӄ��@q��ò�3@!�&�l�!?p���U(�@�n;ha�ٿOӄ��@q��ò�3@!�&�l�!?p���U(�@	mI6"�ٿĥ�M�a�@�C���3@��4
�!?��Ld�@�����ٿ홫F��@sN�0�4@#bh�O�!?P�tVÕ@�����ٿ홫F��@sN�0�4@#bh�O�!?P�tVÕ@�fh�Ǟٿ�c|e�v�@	&"���3@C���!?��1k�@�fh�Ǟٿ�c|e�v�@	&"���3@C���!?��1k�@�fh�Ǟٿ�c|e�v�@	&"���3@C���!?��1k�@�JRF�ٿK�����@�M�/�)4@4��q-�!?%�"<�@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@�K�%�ٿӻ�oԯ�@o:T$�4@�V��!?�NU{��@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@XT���ٿ_�Fΰ�@BG��#4@@��B:�!?S�B�Y�@�CH���ٿ�ĳ��Y�@a�4)�44@|^:t�!?.X�~�@�CH���ٿ�ĳ��Y�@a�4)�44@|^:t�!?.X�~�@�CH���ٿ�ĳ��Y�@a�4)�44@|^:t�!?.X�~�@�CH���ٿ�ĳ��Y�@a�4)�44@|^:t�!?.X�~�@�CH���ٿ�ĳ��Y�@a�4)�44@|^:t�!?.X�~�@ƚ�U��ٿm��:��@B�H4@Vi�1�!?hb�n�0�@ƚ�U��ٿm��:��@B�H4@Vi�1�!?hb�n�0�@ƚ�U��ٿm��:��@B�H4@Vi�1�!?hb�n�0�@pq�@�ٿ ( ����@e�~b�I4@Mғ�!?�S�$d�@pq�@�ٿ ( ����@e�~b�I4@Mғ�!?�S�$d�@pq�@�ٿ ( ����@e�~b�I4@Mғ�!?�S�$d�@pq�@�ٿ ( ����@e�~b�I4@Mғ�!?�S�$d�@pq�@�ٿ ( ����@e�~b�I4@Mғ�!?�S�$d�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@�5W^�ٿ�z��C0�@l��4@5-���!?�5mr�$�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@����ٿ	��\0U�@�s��4@+�߇e�!?o�%ב�@pR��S�ٿ�2�ϛ9�@����3@���[�!?�C|��`�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�ޜ��ٿg>�PU��@�(�n;4@;ۃ6h�!?܍iC�@�-u���ٿs�Ta�@��\�;4@��t��!?{6��]v�@�-u���ٿs�Ta�@��\�;4@��t��!?{6��]v�@�-u���ٿs�Ta�@��\�;4@��t��!?{6��]v�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@4ݠ���ٿl�;��&�@	��G��3@�fC'<�!?f�$-�c�@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@��߇��ٿjf�d'��@%�j`!4@x\M��!?����@IWHқٿ��F�ȏ�@��ʚG4@���Qn�!?�6|�/!�@IWHқٿ��F�ȏ�@��ʚG4@���Qn�!?�6|�/!�@2h݃��ٿ��MN��@KBΟ�G4@,1�d�!?�ϳ+=B�@2h݃��ٿ��MN��@KBΟ�G4@,1�d�!?�ϳ+=B�@2h݃��ٿ��MN��@KBΟ�G4@,1�d�!?�ϳ+=B�@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@�IhBF�ٿ�޾&��@\_�BE4@�D��2�!?���ؕ@��y?��ٿ�v��G�@�j��hN4@�H|\�!?�{�ip�@��y?��ٿ�v��G�@�j��hN4@�H|\�!?�{�ip�@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@��;P�ٿwHS��@��ː4@!ѷ��!?c��5��@�1,h��ٿ��z�q�@���u0�3@�|��p�!?��� �@�1,h��ٿ��z�q�@���u0�3@�|��p�!?��� �@�r9t�ٿ)}�=�@��np�.4@�Kj��!?z�*�/�@��L��ٿ�4�m�J�@h�M��4@r��!f�!?B�Z��5�@��L��ٿ�4�m�J�@h�M��4@r��!f�!?B�Z��5�@��L��ٿ�4�m�J�@h�M��4@r��!f�!?B�Z��5�@��L��ٿ�4�m�J�@h�M��4@r��!f�!?B�Z��5�@	�	�%�ٿ#n��@�n�c�3@y�5]�!?WE�c(�@b��Q�ٿ��g���@JZ�(�4@�F�_}�!?Lÿ�ܕ@b��Q�ٿ��g���@JZ�(�4@�F�_}�!?Lÿ�ܕ@b��Q�ٿ��g���@JZ�(�4@�F�_}�!?Lÿ�ܕ@b��Q�ٿ��g���@JZ�(�4@�F�_}�!?Lÿ�ܕ@b��Q�ٿ��g���@JZ�(�4@�F�_}�!?Lÿ�ܕ@���悞ٿ���B��@�i0|34@~�uz_�!?,�g�>�@(�>W��ٿ�L`:��@�<R�C4@�qh��!?\ziiR�@�e�m�ٿ묅G��@�O��#4@M�*d�!?����h�@���T�ٿ�_���@��t4@���~�!?�m�y�@���T�ٿ�_���@��t4@���~�!?�m�y�@���T�ٿ�_���@��t4@���~�!?�m�y�@���T�ٿ�_���@��t4@���~�!?�m�y�@/����ٿ�3{��y�@c�sue�3@�gPM��!?h�[���@/����ٿ�3{��y�@c�sue�3@�gPM��!?h�[���@/����ٿ�3{��y�@c�sue�3@�gPM��!?h�[���@/����ٿ�3{��y�@c�sue�3@�gPM��!?h�[���@O�VĝٿU��L8��@�Re�4@��t'�!?Vå����@3����ٿ�������@ �c��3@h��j�!?��^�>��@3����ٿ�������@ �c��3@h��j�!?��^�>��@�Q�9��ٿY����@��/z�3@K��!?!�Y����@����ٿ	W5��@	Xȴ��3@�ZS"�!?�}�0`֕@����ٿ	W5��@	Xȴ��3@�ZS"�!?�}�0`֕@����ٿ	W5��@	Xȴ��3@�ZS"�!?�}�0`֕@XM���ٿK�����@��X>��3@%�PQ)�!?zF=TT�@:��tϣٿt-cd ��@aU˖@�3@����D�!??B��A�@:��tϣٿt-cd ��@aU˖@�3@����D�!??B��A�@:��tϣٿt-cd ��@aU˖@�3@����D�!??B��A�@:��tϣٿt-cd ��@aU˖@�3@����D�!??B��A�@"��|��ٿ\�	<Ϗ�@��5�4@�Yr�!?�U�Ou�@ xT��ٿ����@*uXp4@��!O�!?�8��U�@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@b\��ƞٿI+����@m�[�4@�g�\�!?m���@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@!��9ϗٿ���4�@��|m$4@���5�!?")v�@bbJ�r�ٿ��4��@aFy�4@�p
�A�!?F�|)x��@bbJ�r�ٿ��4��@aFy�4@�p
�A�!?F�|)x��@bbJ�r�ٿ��4��@aFy�4@�p
�A�!?F�|)x��@bbJ�r�ٿ��4��@aFy�4@�p
�A�!?F�|)x��@�H�}�ٿ�O�m�b�@�l�� W4@��\-��!?��K��@�H�}�ٿ�O�m�b�@�l�� W4@��\-��!?��K��@�H�}�ٿ�O�m�b�@�l�� W4@��\-��!?��K��@�H�}�ٿ�O�m�b�@�l�� W4@��\-��!?��K��@����Q�ٿb�'��v�@�����I4@N��e�!?���/h��@����Q�ٿb�'��v�@�����I4@N��e�!?���/h��@����Q�ٿb�'��v�@�����I4@N��e�!?���/h��@����Q�ٿb�'��v�@�����I4@N��e�!?���/h��@����Q�ٿb�'��v�@�����I4@N��e�!?���/h��@7�����ٿ�렰��@5k�$4@�/0:�!?C��ɨ��@7�����ٿ�렰��@5k�$4@�/0:�!?C��ɨ��@7�����ٿ�렰��@5k�$4@�/0:�!?C��ɨ��@�ƈO�ٿR燧׾�@X�-���3@�;3�!?�zEqѕ@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@�L�țٿl�OK��@Js1
�"4@m��Ő!?v(��o��@cF6���ٿ��4�~�@T�,�_ 4@��b�x�!?u�c���@cF6���ٿ��4�~�@T�,�_ 4@��b�x�!?u�c���@cF6���ٿ��4�~�@T�,�_ 4@��b�x�!?u�c���@cF6���ٿ��4�~�@T�,�_ 4@��b�x�!?u�c���@cF6���ٿ��4�~�@T�,�_ 4@��b�x�!?u�c���@5�$���ٿ�W���;�@�Es�C�3@f4[nl�!?���ko=�@5�$���ٿ�W���;�@�Es�C�3@f4[nl�!?���ko=�@�$x._�ٿ[:����@��Q�+�3@ۢ�r/�!?�\?���@�$x._�ٿ[:����@��Q�+�3@ۢ�r/�!?�\?���@[�.�ٿ�^_`�@j}c9�3@� Ă�!?�m�[�@[�.�ٿ�^_`�@j}c9�3@� Ă�!?�m�[�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@\U@�2�ٿ�۠���@5T9�3@̕
��!?�:�Έa�@��ã^�ٿj���s�@6�\� 4@;��/�!?JSt��@��ã^�ٿj���s�@6�\� 4@;��/�!?JSt��@��ã^�ٿj���s�@6�\� 4@;��/�!?JSt��@��ã^�ٿj���s�@6�\� 4@;��/�!?JSt��@�\�YٿP�����@����3@a���!?>��]N�@�\�YٿP�����@����3@a���!?>��]N�@�\�YٿP�����@����3@a���!?>��]N�@�\�YٿP�����@����3@a���!?>��]N�@�\�YٿP�����@����3@a���!?>��]N�@b<�T�ٿ��_�+��@�i�(1�3@ ��3�!?+�i��J�@b<�T�ٿ��_�+��@�i�(1�3@ ��3�!?+�i��J�@dO��l�ٿ=2Y�0��@��r.@4@=c{bD�!?�����@dO��l�ٿ=2Y�0��@��r.@4@=c{bD�!?�����@�n]�ٿ�����@���	4@0�l7�!?�I߀��@�n]�ٿ�����@���	4@0�l7�!?�I߀��@-��ҧٿGu�}Gs�@����U4@cV��0�!?1��Q�@-��ҧٿGu�}Gs�@����U4@cV��0�!?1��Q�@-��ҧٿGu�}Gs�@����U4@cV��0�!?1��Q�@��E�%�ٿ�J2m=�@3����4@�����!?���D"�@��E�%�ٿ�J2m=�@3����4@�����!?���D"�@��E�%�ٿ�J2m=�@3����4@�����!?���D"�@��t���ٿ�W�e��@kCg4@�VQI_�!?�.&���@��t���ٿ�W�e��@kCg4@�VQI_�!?�.&���@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@=�?:5�ٿHp�^p�@�����)4@�r� ��!?�Kq�@I|�sL�ٿ���i��@���m;4@@賁�!?9����@:tC��ٿ�ԛ-|��@j��@4@"��I�!?pQ��'�@&�ꑖٿEܵ����@��d"d4@D�`&U�!?���@�@&�ꑖٿEܵ����@��d"d4@D�`&U�!?���@�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@�e�"�ٿ�%{���@�2�?N4@F���!?�J{
�@W�;-��ٿ�� �:�@�8�� 4@jq�r��!?w�c/��@W�;-��ٿ�� �:�@�8�� 4@jq�r��!?w�c/��@W�;-��ٿ�� �:�@�8�� 4@jq�r��!?w�c/��@�*�x��ٿ�\}�dE�@����4@�D�KK�!?Ը�ƕ@�*�x��ٿ�\}�dE�@����4@�D�KK�!?Ը�ƕ@��4�Y�ٿ'�]����@����R4@�� B��!?Ck;W�@��q8o�ٿwHr����@@�
��84@K�u�{�!?����MЕ@��q8o�ٿwHr����@@�
��84@K�u�{�!?����MЕ@��q8o�ٿwHr����@@�
��84@K�u�{�!?����MЕ@��q8o�ٿwHr����@@�
��84@K�u�{�!?����MЕ@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@Oa��ٿ�U����@FCc�L4@ ���4�!?�Z���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@|�%���ٿÿ����@T�1�D4@�z�]�!?F�^(���@2�;ϜٿM"����@�K���4@#B�N�!?
R]V4�@2�;ϜٿM"����@�K���4@#B�N�!?
R]V4�@2�;ϜٿM"����@�K���4@#B�N�!?
R]V4�@�z�}��ٿ��uh5��@r��+&94@zu��p�!?�t��9�@�z�}��ٿ��uh5��@r��+&94@zu��p�!?�t��9�@�z�}��ٿ��uh5��@r��+&94@zu��p�!?�t��9�@�z�}��ٿ��uh5��@r��+&94@zu��p�!?�t��9�@�z�}��ٿ��uh5��@r��+&94@zu��p�!?�t��9�@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��*��ٿ�x8��.�@��E4@�% _L�!?`t����@��8��ٿc���M2�@`6��U4@�z;�!?�>6$�@��8��ٿc���M2�@`6��U4@�z;�!?�>6$�@��8��ٿc���M2�@`6��U4@�z;�!?�>6$�@��8��ٿc���M2�@`6��U4@�z;�!?�>6$�@��8��ٿc���M2�@`6��U4@�z;�!?�>6$�@�q�C�ٿ"������@��\,4@L�5���!?/��-�@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���x�ٿS5S�@p��j�H4@:#u��!?�_Sd���@���|��ٿ
\|���@�PɮD4@�V �M�!?2%�����@��p7ƚٿ��oQ�@/^�3@�u�#�!?��.Pͫ�@��p7ƚٿ��oQ�@/^�3@�u�#�!?��.Pͫ�@��p7ƚٿ��oQ�@/^�3@�u�#�!?��.Pͫ�@��p7ƚٿ��oQ�@/^�3@�u�#�!?��.Pͫ�@��p7ƚٿ��oQ�@/^�3@�u�#�!?��.Pͫ�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@�u���ٿ���!�@����3@�CfY�!?ė�.�@A�ٿ^h���@�@���m��3@T���N�!?+٘�G�@A�ٿ^h���@�@���m��3@T���N�!?+٘�G�@A�ٿ^h���@�@���m��3@T���N�!?+٘�G�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@����s�ٿx�"[��@�Y�_�84@�'�!?
��
�*�@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@��B�a�ٿנ߹�D�@�y#E4@a�w>�!?o>�����@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@���W�ٿ��}��@w/��*e4@:�YL�!?�Cr���@�@�ٿz
�o��@$�LY4@��+�!?�����@�@�ٿz
�o��@$�LY4@��+�!?�����@�@�ٿz
�o��@$�LY4@��+�!?�����@1���ٿT+u�{��@nz��H4@U�^|B�!?��v�%�@1���ٿT+u�{��@nz��H4@U�^|B�!?��v�%�@1���ٿT+u�{��@nz��H4@U�^|B�!?��v�%�@1���ٿT+u�{��@nz��H4@U�^|B�!?��v�%�@?p�$�ٿ����w�@�'q�04@z�O3�!?"�|Y�#�@?p�$�ٿ����w�@�'q�04@z�O3�!?"�|Y�#�@��\��ٿ%�QP!��@�����3@�M+U�!?�%�8jH�@��\��ٿ%�QP!��@�����3@�M+U�!?�%�8jH�@��E|�ٿ�E�lJ}�@��_\d;4@N����!?=r�(��@��E|�ٿ�E�lJ}�@��_\d;4@N����!?=r�(��@#K4�ٿ�F:��5�@[�̣74@)Vuӏ!?������@#K4�ٿ�F:��5�@[�̣74@)Vuӏ!?������@#K4�ٿ�F:��5�@[�̣74@)Vuӏ!?������@#K4�ٿ�F:��5�@[�̣74@)Vuӏ!?������@�'T�ٿ�y�b�@I痫)4@�R��!?�`���@�'T�ٿ�y�b�@I痫)4@�R��!?�`���@�'T�ٿ�y�b�@I痫)4@�R��!?�`���@@-�̬�ٿ�𒏤&�@�����'4@�⨏!?����@�����ٿ3ھ���@A9���4@'(�܏!?N$���@�����ٿ3ھ���@A9���4@'(�܏!?N$���@�����ٿ3ھ���@A9���4@'(�܏!?N$���@�����ٿ3ھ���@A9���4@'(�܏!?N$���@�����ٿ3ھ���@A9���4@'(�܏!?N$���@�����ٿ3ھ���@A9���4@'(�܏!?N$���@R �֖ٿ������@ih6�F$4@y6��!?ۥ��ʕ@R �֖ٿ������@ih6�F$4@y6��!?ۥ��ʕ@R �֖ٿ������@ih6�F$4@y6��!?ۥ��ʕ@R �֖ٿ������@ih6�F$4@y6��!?ۥ��ʕ@�ov^k�ٿA��{ �@��3��4@ˢB�!?�`vTV��@�ov^k�ٿA��{ �@��3��4@ˢB�!?�`vTV��@�o���ٿ��o�'�@���24@Tore5�!?����	�@�o���ٿ��o�'�@���24@Tore5�!?����	�@I��O�ٿ��0����@��-�4@�]�qk�!?���䤕@�8�ٿh�����@H�Q�	44@%��N�!?��e2���@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@f��@�ٿ�9�fK�@��(L`4@2���I�!?A鋃͛�@�ݻ5�ٿ���"���@���4@���o7�!?�����@sXsW�ٿ�uf��=�@&.�̺04@�Y�-�!?Ew�<��@dPi��ٿP;��x�@5R4z�H4@�浄�!?a��@Q�
@��ٿ�i%p>�@��^K@E4@ćo�K�!?����	�@Q�
@��ٿ�i%p>�@��^K@E4@ćo�K�!?����	�@Q�
@��ٿ�i%p>�@��^K@E4@ćo�K�!?����	�@Q�
@��ٿ�i%p>�@��^K@E4@ćo�K�!?����	�@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@�sb���ٿ-���hP�@"�R+)4@-%W�!?����Sϕ@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@��k1I�ٿ���,���@�u�Ij94@ ��պ�!?I$6���@_��6�ٿ��`9��@�A��54@���s�!?�P��@_��6�ٿ��`9��@�A��54@���s�!?�P��@_��6�ٿ��`9��@�A��54@���s�!?�P��@_��6�ٿ��`9��@�A��54@���s�!?�P��@_��6�ٿ��`9��@�A��54@���s�!?�P��@_��6�ٿ��`9��@�A��54@���s�!?�P��@�_��ٿp̙����@�����3@��},R�!?{"�nf�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@�ڗ*�ٿ?CIw��@�o�3@Q��f�!?��/Q�@����ɡٿ&ul?>��@s�f[�3@0��>H�!?����̕@����ɡٿ&ul?>��@s�f[�3@0��>H�!?����̕@v��.�ٿВ�s�&�@�(��4@��Z �!?Y��h��@�n�C�ٿU�ˇ�2�@׶�e�(4@,A)�F�!?{�����@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@h�|[~�ٿMG�8-�@�j�-4@�+K*_�!?_�r��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@���śٿh��@�t�}+4@��BMR�!?��u��@�7Y��ٿ�g�+L�@��F.�+4@ɽŊ|�!?J��-�ȕ@�7Y��ٿ�g�+L�@��F.�+4@ɽŊ|�!?J��-�ȕ@�7Y��ٿ�g�+L�@��F.�+4@ɽŊ|�!?J��-�ȕ@�7Y��ٿ�g�+L�@��F.�+4@ɽŊ|�!?J��-�ȕ@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�Cp�ٿ�H"C�X�@�zâ4@=���?�!?�S��z��@�n x��ٿ��ʹ��@rs���4@�&R��!?�l]��ɕ@�n x��ٿ��ʹ��@rs���4@�&R��!?�l]��ɕ@�n x��ٿ��ʹ��@rs���4@�&R��!?�l]��ɕ@�n x��ٿ��ʹ��@rs���4@�&R��!?�l]��ɕ@�n x��ٿ��ʹ��@rs���4@�&R��!?�l]��ɕ@\L�w�ٿ��:Vj�@Л�a4@���?q�!?�����@\L�w�ٿ��:Vj�@Л�a4@���?q�!?�����@\L�w�ٿ��:Vj�@Л�a4@���?q�!?�����@\L�w�ٿ��:Vj�@Л�a4@���?q�!?�����@J��+G�ٿ`v����@r� �>4@=�Γ!�!?�=�3e��@I����ٿ�e��@��I!�?4@���W�!?g��^|�@I����ٿ�e��@��I!�?4@���W�!?g��^|�@1�\��ٿ�����=�@��`Er34@��`1��!?Ȥ琞��@ʘ.�ٿ����j��@^Jr�c4@�c�!?��ݕ@�NMH-�ٿ��(�@=�p,#4@?oټ[�!?�+�w+�@��[7n�ٿTs��M��@���4@ ա|�!?	oCR��@��[7n�ٿTs��M��@���4@ ա|�!?	oCR��@��[7n�ٿTs��M��@���4@ ա|�!?	oCR��@;��	�ٿ�N|�p6�@'��6�#4@�`��o�!?�<й��@;��	�ٿ�N|�p6�@'��6�#4@�`��o�!?�<й��@� _�N�ٿr�p��@�����3@@N��4�!?]���\�@� _�N�ٿr�p��@�����3@@N��4�!?]���\�@N*�	/�ٿU�eqW�@6ē�O4@Zpz�a�!?�aj}�U�@R7n�ٿ;�e��@�I�IG4@��۩0�!?�r�ブ@�H��!�ٿ����j�@�a���3@������!?��,/^�@|��A�ٿ�r�t�@S`G� 4@Va�!a�!?���T�@|��A�ٿ�r�t�@S`G� 4@Va�!a�!?���T�@jԊV~�ٿ>�oߊ�@|��3@��R�!?���2��@jԊV~�ٿ>�oߊ�@|��3@��R�!?���2��@�Rv��ٿp�\���@8?��W;4@�&74V�!?X;s����@�Rv��ٿp�\���@8?��W;4@�&74V�!?X;s����@�Rv��ٿp�\���@8?��W;4@�&74V�!?X;s����@�:ͯq�ٿ{������@�����O4@�����!?T��\��@��Υ�ٿ��
`�j�@��|]�e4@��<K9�!?�3�"_�@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@{�R��ٿ�ekI���@��r��24@�Cj22�!?�5j��@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�~�w��ٿ�y�1�u�@�o5�U4@�l�t�!?S�E�_�@�n�{��ٿ�Z+^��@�"{G4@ެ"�<�!?]NM�U�@�n�{��ٿ�Z+^��@�"{G4@ެ"�<�!?]NM�U�@�n�{��ٿ�Z+^��@�"{G4@ެ"�<�!?]NM�U�@ǩs�~�ٿdG�f�@(>+N+4@�dL�!?�V����@ǩs�~�ٿdG�f�@(>+N+4@�dL�!?�V����@ˊ]rq�ٿ��v"��@~�2	4@ė�j;�!??�F�@ˊ]rq�ٿ��v"��@~�2	4@ė�j;�!??�F�@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@���|V�ٿ��YT���@&Y��4@��ۀ�!?�o:��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@�n���ٿ��Ĵ�Z�@nW���4@�f�G�!?�s��a��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@uR�{3�ٿ|�c`��@G��5�94@�;ID*�!?��?<��@:ڨ `�ٿ�=Dsv�@�!8E4@����8�!?H�*+�@:ڨ `�ٿ�=Dsv�@�!8E4@����8�!?H�*+�@:ڨ `�ٿ�=Dsv�@�!8E4@����8�!?H�*+�@:ڨ `�ٿ�=Dsv�@�!8E4@����8�!?H�*+�@:ڨ `�ٿ�=Dsv�@�!8E4@����8�!?H�*+�@`�����ٿv!�Ƞ�@�m��4@M[�	b�!?�u��f�@6�Cp�ٿGα����@�@�G�74@B��\�!?�!$���@6�Cp�ٿGα����@�@�G�74@B��\�!?�!$���@���U7�ٿ�<f���@�����v4@�] �b�!?3����@���U7�ٿ�<f���@�����v4@�] �b�!?3����@���U7�ٿ�<f���@�����v4@�] �b�!?3����@���U7�ٿ�<f���@�����v4@�] �b�!?3����@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@��
���ٿܯE-n��@Qt�_4@dI�x�!?^)b�WP�@4s��ɖٿ��A����@�s��_P4@�Z9��!?��B�:�@�"���ٿ��ҥ�.�@h�	4@�B� l�!?lHm3�5�@ ��\�ٿ�4�a��@V�n�v74@�z��n�!?x�Y�7��@ ��\�ٿ�4�a��@V�n�v74@�z��n�!?x�Y�7��@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@��$�ٿ-
ds�@�eC�4@�"�.�!?`,�Ҳ�@���R�ٿ"GD�̟�@�w�h� 4@>�K"c�!?_7�,k��@��3J�ٿ�������@5앹��3@R���w�!?�����@��<�ٿ�!0< ��@�
p�"?4@V~��o�!?��&��@��<�ٿ�!0< ��@�
p�"?4@V~��o�!?��&��@��<�ٿ�!0< ��@�
p�"?4@V~��o�!?��&��@��<�ٿ�!0< ��@�
p�"?4@V~��o�!?��&��@#Ekɘٿ�E+ξt�@A��bC4@��>�%�!?�0#{�̕@#Ekɘٿ�E+ξt�@A��bC4@��>�%�!?�0#{�̕@#Ekɘٿ�E+ξt�@A��bC4@��>�%�!?�0#{�̕@��9&�ٿ���6�S�@�LZ͘�3@��vu�!?*�Z���@��9&�ٿ���6�S�@�LZ͘�3@��vu�!?*�Z���@�HSM=�ٿ#�Θ�;�@�9�4@�
�v�!?������@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@x�(
�ٿ��D1\�@�D=*4@پ��!?
��喕@�У,�ٿPc;��(�@�a
A�4@� Q���!?	�V$��@�У,�ٿPc;��(�@�a
A�4@� Q���!?	�V$��@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@��+��ٿ �Uli �@�8��4@���?�!?�x��E�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@�q����ٿ��UUFe�@4��4@p��T�!?4��	_1�@��>$3�ٿ�]�����@�>pQ�4@�\I6L�!?�P7}4�@��>$3�ٿ�]�����@�>pQ�4@�\I6L�!?�P7}4�@�'	�ٿ��/� �@�y��74@�%T�\�!?Z��$
�@�'	�ٿ��/� �@�y��74@�%T�\�!?Z��$
�@�'	�ٿ��/� �@�y��74@�%T�\�!?Z��$
�@�'	�ٿ��/� �@�y��74@�%T�\�!?Z��$
�@�'	�ٿ��/� �@�y��74@�%T�\�!?Z��$
�@xˆ+U�ٿy�~��@�H.�[4@��b\�!?u���6�@儬�
�ٿ�Q���@
w���04@f�t�/�!?�0���b�@儬�
�ٿ�Q���@
w���04@f�t�/�!?�0���b�@儬�
�ٿ�Q���@
w���04@f�t�/�!?�0���b�@�)�ҙٿ��t	��@�HW4@�c��!?��Ѣ[�@����ٿ7���"��@��C��3@�7�r�!?�O�r��@����ٿ7���"��@��C��3@�7�r�!?�O�r��@�}~���ٿ��c�M�@�L�3�3@�����!?a���@�}~���ٿ��c�M�@�L�3�3@�����!?a���@�#�V�ٿ|��!Ն�@^�m�B44@r`��R�!?L���v�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�e��͚ٿ�����8�@��c24@\�Y8�!?,�2_0�@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@�V��ٿ���w�@G���==4@zsF]�!?y}|Õ@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@���E�ٿ�r8� �@�/��0P4@9�1�E�!?�E���@9�@ ��ٿ�/h`���@[�.e4@�vgW�!?��] �@9�@ ��ٿ�/h`���@[�.e4@�vgW�!?��] �@9�@ ��ٿ�/h`���@[�.e4@�vgW�!?��] �@9�@ ��ٿ�/h`���@[�.e4@�vgW�!?��] �@Ѻ�_��ٿ6z�e�f�@aw
W��3@����a�!?���	|/�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@��R���ٿ�]c�	�@ǠІ�3@Gб]�!?�"�3y�@ ����ٿ,�"g��@�`8�94@��o ��!?x��v8�@ ����ٿ,�"g��@�`8�94@��o ��!?x��v8�@MAې7�ٿ�����@���f�4@	򦌐!?K��A�@MAې7�ٿ�����@���f�4@	򦌐!?K��A�@���ٿd�dkf*�@@_n�4@/਄��!?�bM'��@���ٿd�dkf*�@@_n�4@/਄��!?�bM'��@���ٿd�dkf*�@@_n�4@/਄��!?�bM'��@���ٿd�dkf*�@@_n�4@/਄��!?�bM'��@���ٿd�dkf*�@@_n�4@/਄��!?�bM'��@��~�y�ٿ��<�4��@N4и 4@�)c��!?�7�ᎉ�@��~�y�ٿ��<�4��@N4и 4@�)c��!?�7�ᎉ�@��~�y�ٿ��<�4��@N4и 4@�)c��!?�7�ᎉ�@��~�y�ٿ��<�4��@N4и 4@�)c��!?�7�ᎉ�@@ ��ٿH;=��@�7ҿ64@+eB��!?�_O鬂�@@ ��ٿH;=��@�7ҿ64@+eB��!?�_O鬂�@@ ��ٿH;=��@�7ҿ64@+eB��!?�_O鬂�@�?�%�ٿ�Zk�>c�@TSJ4<4@��׼�!?p�껼�@�?�%�ٿ�Zk�>c�@TSJ4<4@��׼�!?p�껼�@���"��ٿ��9�m`�@���d�4@����!?ׁM���@���"��ٿ��9�m`�@���d�4@����!?ׁM���@���"��ٿ��9�m`�@���d�4@����!?ׁM���@���"��ٿ��9�m`�@���d�4@����!?ׁM���@0;�G�ٿBP֬���@���\%4@�&��r�!?��}�i�@0;�G�ٿBP֬���@���\%4@�&��r�!?��}�i�@��ȭ�ٿ��˽ �@�2�u�4@�Z�_`�!?*r�@]��O�ٿH3N�v/�@��S�4@��t��!?������@]��O�ٿH3N�v/�@��S�4@��t��!?������@����|�ٿsNݕ���@0EkA�4@��o��!?ݨ=g"j�@�H���ٿ�lV�U�@R�ǹ�3@L�߾ڐ!?��].~�@"�@P*�ٿ�Ė"���@ =�3*24@2���ݐ!?y	a0�1�@"�@P*�ٿ�Ė"���@ =�3*24@2���ݐ!?y	a0�1�@>��ɱ�ٿ=�bw��@��Շl4@���7��!?!9�b��@1�^�ٿm�$���@�^��"�3@�.!Đ!?e��۟S�@1�^�ٿm�$���@�^��"�3@�.!Đ!?e��۟S�@v��ٿ���͟��@��j��3@�$ӧ��!?�I��~��@-�\
S�ٿ$�CK�`�@�H���3@�VX]
�!?ti8N˕@-�\
S�ٿ$�CK�`�@�H���3@�VX]
�!?ti8N˕@-�\
S�ٿ$�CK�`�@�H���3@�VX]
�!?ti8N˕@� އ��ٿ ����@NKPR�3@CB�$`�!?��Y�ڹ�@� އ��ٿ ����@NKPR�3@CB�$`�!?��Y�ڹ�@�Gp_1�ٿ�B�c�@S��AT�3@`A�Q^�!?�0V��Е@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��Ҳ��ٿC)���x�@` R��3@ٓB�Z�!?R�]�h�@��ζ�ٿ�U����@���'��3@G,C�,�!?@��p��@��ζ�ٿ�U����@���'��3@G,C�,�!?@��p��@bq���ٿ>�����@M����4@�Vfu�!?�C��fJ�@�W��ٿ��E��@"p��4@'�QT�!?~������@�W��ٿ��E��@"p��4@'�QT�!?~������@�W��ٿ��E��@"p��4@'�QT�!?~������@�Y�@k�ٿɺ%�x�@Vl�3)4@� �Ph�!?�b�}Jԕ@�Y�@k�ٿɺ%�x�@Vl�3)4@� �Ph�!?�b�}Jԕ@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@����ٿ_���1��@\,v��4@����Z�!?�qI.���@��)�l�ٿ8:��L��@Q�deS4@��6�!?o�T:���@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@~�P*��ٿ>U�bz+�@�q]3<4@f�CNP�!?f����A�@'�[FЗٿ��� ��@<�`��M4@/�!?�퍮��@'�[FЗٿ��� ��@<�`��M4@/�!?�퍮��@'�[FЗٿ��� ��@<�`��M4@/�!?�퍮��@�E2r��ٿ�v"����@rK�V4@mz{A�!?�_6�BÕ@�E2r��ٿ�v"����@rK�V4@mz{A�!?�_6�BÕ@��]�_�ٿ�\��Z��@[���4@�g��!?Z�>���@�%vZ՞ٿ<8B�U�@f����3@>�L�B�!?)%�\8�@�%vZ՞ٿ<8B�U�@f����3@>�L�B�!?)%�\8�@*|%�ٿ!�+(��@sl�Im4@3�a�
�!?>�����@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@t�qq̝ٿ�n�$��@=��P�<4@+����!?q6�z��@��䢢ٿ[
Z	���@��x�I4@3D(�!?�wЏ��@��䢢ٿ[
Z	���@��x�I4@3D(�!?�wЏ��@��䢢ٿ[
Z	���@��x�I4@3D(�!?�wЏ��@��䢢ٿ[
Z	���@��x�I4@3D(�!?�wЏ��@=���5�ٿ`�dP)��@���JM-4@9z5Ӑ�!?��(�Qc�@=���5�ٿ`�dP)��@���JM-4@9z5Ӑ�!?��(�Qc�@=���5�ٿ`�dP)��@���JM-4@9z5Ӑ�!?��(�Qc�@=���5�ٿ`�dP)��@���JM-4@9z5Ӑ�!?��(�Qc�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@��6�Ɯٿ��Qzr��@�]_j*4@�JJ�!?{Ô&dj�@~Ul�ٿ���@��@��r9�64@�f7��!?�Q�V�@~Ul�ٿ���@��@��r9�64@�f7��!?�Q�V�@~Ul�ٿ���@��@��r9�64@�f7��!?�Q�V�@~Ul�ٿ���@��@��r9�64@�f7��!?�Q�V�@~Ul�ٿ���@��@��r9�64@�f7��!?�Q�V�@V#��ٿ���-�@T���4@π1b��!?��f��@�9��+�ٿ�Y��V�@�����K4@�h���!?��V���@�/��ٿd�CU��@���ǫG4@:4�P��!?7��+ڕ@�/��ٿd�CU��@���ǫG4@:4�P��!?7��+ڕ@�/��ٿd�CU��@���ǫG4@:4�P��!?7��+ڕ@�/��ٿd�CU��@���ǫG4@:4�P��!?7��+ڕ@�4��W�ٿIBmb��@��%��f4@mMdd�!?���y)��@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@�C勉�ٿ0�>b��@�.6C�>4@����5�!?�Y�5L�@B5����ٿ���R��@�K�@g4@KAGNC�!?�c��8a�@B5����ٿ���R��@�K�@g4@KAGNC�!?�c��8a�@B5����ٿ���R��@�K�@g4@KAGNC�!?�c��8a�@B5����ٿ���R��@�K�@g4@KAGNC�!?�c��8a�@B5����ٿ���R��@�K�@g4@KAGNC�!?�c��8a�@>�����ٿ��#��@ڭ?D�04@��d��!?h�Y�	�@>�����ٿ��#��@ڭ?D�04@��d��!?h�Y�	�@>�����ٿ��#��@ڭ?D�04@��d��!?h�Y�	�@>�����ٿ��#��@ڭ?D�04@��d��!?h�Y�	�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@��|q��ٿ���#���@ei�T�N4@/�D1�!?T�G�&�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���{��ٿ�;g���@Ör�V4@��<�4�!?�@��'�@���F3�ٿ~�%���@e�sq4@e�?x�!? �>��@"dA{�ٿ%{h��@; 9��,4@�?�D�!?53AG�@"dA{�ٿ%{h��@; 9��,4@�?�D�!?53AG�@"dA{�ٿ%{h��@; 9��,4@�?�D�!?53AG�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@}���ٿ�j�N�@���dB4@� ���!?1(;�C�@����ٿ\���E��@N�(�4@ٲ� �!?Зc���@����ٿ\���E��@N�(�4@ٲ� �!?Зc���@b��Ρٿ���N�@�$��3@�Pw��!?%��-�@���ρ�ٿ�]�D	�@���bu�3@�jQkj�!?��׫�,�@�W-��ٿ;�o�A��@n��U4@X(`r�!?�Y��+�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@g�Rm�ٿ>DO~���@9���3@4�h���!?�Z�h	x�@�g�ٿe},���@ �r���3@�4�
0�!?)�*���@�g�ٿe},���@ �r���3@�4�
0�!?)�*���@P/�>c�ٿDV4�4h�@�oJj�"4@���!?�3w$^�@P/�>c�ٿDV4�4h�@�oJj�"4@���!?�3w$^�@4���ٿ�����@<W5��4@�C�p�!?l}L�<S�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@�-L��ٿ��d?�@[���44@j�岌�!?���}�p�@3�ܖٿ4�,���@lR��3@��h�t�!?�^d#ʦ�@3�ܖٿ4�,���@lR��3@��h�t�!?�^d#ʦ�@3�ܖٿ4�,���@lR��3@��h�t�!?�^d#ʦ�@3�ܖٿ4�,���@lR��3@��h�t�!?�^d#ʦ�@3�ܖٿ4�,���@lR��3@��h�t�!?�^d#ʦ�@ƀ�gG�ٿZX� ��@�t})�3@b]�2ϐ!?�@W[��@~�X�G�ٿ�z�[]�@��lcg�3@V>�e��!?BǮQ �@~�X�G�ٿ�z�[]�@��lcg�3@V>�e��!?BǮQ �@~�X�G�ٿ�z�[]�@��lcg�3@V>�e��!?BǮQ �@~�X�G�ٿ�z�[]�@��lcg�3@V>�e��!?BǮQ �@E��~@�ٿc��]��@��P_�3@�_꣐!?��[ Z�@E��~@�ٿc��]��@��P_�3@�_꣐!?��[ Z�@E��~@�ٿc��]��@��P_�3@�_꣐!?��[ Z�@����ٿ�h3�-�@���X�3@��߬��!?(O�^�~�@�<�FN�ٿ�٨��7�@��g*�3@_�Pj}�!?N�5��`�@�<�FN�ٿ�٨��7�@��g*�3@_�Pj}�!?N�5��`�@�<�FN�ٿ�٨��7�@��g*�3@_�Pj}�!?N�5��`�@�<�FN�ٿ�٨��7�@��g*�3@_�Pj}�!?N�5��`�@�<�FN�ٿ�٨��7�@��g*�3@_�Pj}�!?N�5��`�@�#⶗ٿ- �����@����K4@���f��!?)�����@�#⶗ٿ- �����@����K4@���f��!?)�����@�#⶗ٿ- �����@����K4@���f��!?)�����@X�$Y��ٿ��Aa�A�@���-4@�LZ2X�!?D���N��@X�$Y��ٿ��Aa�A�@���-4@�LZ2X�!?D���N��@X�$Y��ٿ��Aa�A�@���-4@�LZ2X�!?D���N��@X�$Y��ٿ��Aa�A�@���-4@�LZ2X�!?D���N��@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�M�C�ٿ�ıЌ}�@���4@ h��C�!?/�kx�@�G����ٿw��~{�@����e-4@�SGp�!?��md��@�G����ٿw��~{�@����e-4@�SGp�!?��md��@�H����ٿƈ�zj?�@�eqހ�3@\؞�P�!?`�\�2�@'_���ٿ�R�����@%啙#4@�X�^=�!?{6�O|��@'_���ٿ�R�����@%啙#4@�X�^=�!?{6�O|��@'_���ٿ�R�����@%啙#4@�X�^=�!?{6�O|��@�u@ 6�ٿ�tZg��@�:u���3@lE�5�!?F���X�@?�~�ӟٿ&�4�Uc�@��c�s4@MŌ��!?�Q�3��@?�~�ӟٿ&�4�Uc�@��c�s4@MŌ��!?�Q�3��@?�~�ӟٿ&�4�Uc�@��c�s4@MŌ��!?�Q�3��@?�~�ӟٿ&�4�Uc�@��c�s4@MŌ��!?�Q�3��@?�~�ӟٿ&�4�Uc�@��c�s4@MŌ��!?�Q�3��@z��4�ٿ�mqm�5�@�/g s4@Ţ^K/�!?������@z��4�ٿ�mqm�5�@�/g s4@Ţ^K/�!?������@z��4�ٿ�mqm�5�@�/g s4@Ţ^K/�!?������@z��4�ٿ�mqm�5�@�/g s4@Ţ^K/�!?������@z��4�ٿ�mqm�5�@�/g s4@Ţ^K/�!?������@�[+	�ٿ��Ae�@s�!�^4@�7�N�!?1k|�~˕@�[+	�ٿ��Ae�@s�!�^4@�7�N�!?1k|�~˕@�[+	�ٿ��Ae�@s�!�^4@�7�N�!?1k|�~˕@�[+	�ٿ��Ae�@s�!�^4@�7�N�!?1k|�~˕@�[+	�ٿ��Ae�@s�!�^4@�7�N�!?1k|�~˕@e:����ٿ��l.!��@�8?��n4@3���!?��[�U�@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@!ޡ�Γٿ̾<X,�@��04@~e+��!?��(��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@��G��ٿm� ���@�!*��[4@��l9�!?l#�6��@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�_��S�ٿ'�(=l�@n�T�4@���r�!?��m�7�@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@�Q,Z1�ٿ�h?�I�@�#���3@��*��!?_Gr֥��@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@na���ٿ�R�ڔ�@�0� ��3@��4��!?g����{�@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@�Jo7�ٿ��S��@�F;%��3@O}�\�!?>LZ���@E= h=�ٿ\H�#z��@�8���3@�,���!?5v�n\��@N-^�ןٿ ?M51��@>�)$/~3@H ���!?�"�p�@N-^�ןٿ ?M51��@>�)$/~3@H ���!?�"�p�@N-^�ןٿ ?M51��@>�)$/~3@H ���!?�"�p�@�u�E�ٿ�Ů�B��@�=7��3@���!8�!?`:Z�4��@�u�E�ٿ�Ů�B��@�=7��3@���!8�!?`:Z�4��@9"'t��ٿ�u����@�L�r44@E���4�!?���	y��@9"'t��ٿ�u����@�L�r44@E���4�!?���	y��@� .�کٿR1����@��E4@{����!?�$���ٕ@� .�کٿR1����@��E4@{����!?�$���ٕ@� .�کٿR1����@��E4@{����!?�$���ٕ@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@���D\�ٿu��ǣ�@gر~N�3@Ov�&�!?�po�59�@�rNM�ٿ�⏴���@���S��3@t��tn�!?��/l�@�rNM�ٿ�⏴���@���S��3@t��tn�!?��/l�@�rNM�ٿ�⏴���@���S��3@t��tn�!?��/l�@�rNM�ٿ�⏴���@���S��3@t��tn�!?��/l�@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@+{!�ٿxR5��@0�7h�3@��i���!?`�S��@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@�	�J�ٿ}l�[�@7�ӏ94@*Z&,O�!?���Z�@>)@m�ٿϧ�5��@{�&4@����v�!?��ER�p�@�@;��ٿ]�%kE��@�����4@��8��!?�a�aU�@�@;��ٿ]�%kE��@�����4@��8��!?�a�aU�@�@;��ٿ]�%kE��@�����4@��8��!?�a�aU�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@%ⷘ��ٿ,�i9�@�ze`��3@��矣�!?���/a�@���ǝٿ�fj't�@�
�P�4@[{DP�!?�~����@���ǝٿ�fj't�@�
�P�4@[{DP�!?�~����@���ǝٿ�fj't�@�
�P�4@[{DP�!?�~����@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@�j
���ٿ�x�ީ��@�K�h4@�)Գ�!?�j�<9�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@���ٿRPkq<-�@7�k�,4@nU�Ð!?,/%�8�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@� 3��ٿ	&!x+�@p;�h�Y4@�έ��!?�a>>]�@���ٿ,�3�B�@����+4@Jul`p�!?�m }V��@���ٿ,�3�B�@����+4@Jul`p�!?�m }V��@���ٿ,�3�B�@����+4@Jul`p�!?�m }V��@���ٿ,�3�B�@����+4@Jul`p�!?�m }V��@���ٿ,�3�B�@����+4@Jul`p�!?�m }V��@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�@ɬ�ٿ{�ه��@i��0;4@�<�>�!?��P���@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@�7�ٿ�#a��E�@z�X��4@C<ɐ�!?�e��_Ε@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@���E��ٿ��g���@�i_�$4@@^�w�!?A�1ߕ@V"�ٿ�ɞ3��@�m� 4@��^T�!?�"�|w��@V"�ٿ�ɞ3��@�m� 4@��^T�!?�"�|w��@V"�ٿ�ɞ3��@�m� 4@��^T�!?�"�|w��@V"�ٿ�ɞ3��@�m� 4@��^T�!?�"�|w��@�2L��ٿd��٢��@�2��,.4@q`g��!?=���ϕ@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@�2�ٿ��$��U�@�����4@���T�!?��]�X�@-��ٿ����M�@��F=4@!��Q=�!?�VGD�1�@-��ٿ����M�@��F=4@!��Q=�!?�VGD�1�@�2��ٿ��f_,��@�%м�+4@����O�!?>^&��V�@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@k����ٿ�Qq��f�@��}�NW4@#���`�!?C+Bc��@h̕z�ٿ��/��@|��I4@@�G%��!?d�����@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@Kt	 
�ٿ�"����@[2�P�94@Y�� �!?���K˕@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@�`u�y�ٿ	�Z���@�L
�W4@^��]�!?`�;��@a�`E�ٿ�@�*�@�]7��24@؆�ҹ�!?� ���@a�`E�ٿ�@�*�@�]7��24@؆�ҹ�!?� ���@a�`E�ٿ�@�*�@�]7��24@؆�ҹ�!?� ���@a�`E�ٿ�@�*�@�]7��24@؆�ҹ�!?� ���@a�`E�ٿ�@�*�@�]7��24@؆�ҹ�!?� ���@`˫9�ٿ�����@�&�4@}��~��!?Y��FI��@`˫9�ٿ�����@�&�4@}��~��!?Y��FI��@`˫9�ٿ�����@�&�4@}��~��!?Y��FI��@`˫9�ٿ�����@�&�4@}��~��!?Y��FI��@h��w�ٿy#RȯP�@��X�)4@�C&{�!?�e���@h��w�ٿy#RȯP�@��X�)4@�C&{�!?�e���@h��w�ٿy#RȯP�@��X�)4@�C&{�!?�e���@h��w�ٿy#RȯP�@��X�)4@�C&{�!?�e���@h��w�ٿy#RȯP�@��X�)4@�C&{�!?�e���@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@`�����ٿ�R|	0��@ˑ �4@��~��!?���;7t�@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@��vȚٿ���d��@_a���3@�����!?|�h~��@f��mʛٿ�k���@Z�Fc��3@V	�7��!?@�m��ĕ@f��mʛٿ�k���@Z�Fc��3@V	�7��!?@�m��ĕ@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@l��6��ٿ��d����@�:��3@�<��h�!?G��|��@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@��$���ٿ�ٯ(
+�@|Q�	4@�B{�$�!?z�D]ȉ�@�|�Ξٿ���:���@ԣZm4@G��Y�!?WO�����@�|�Ξٿ���:���@ԣZm4@G��Y�!?WO�����@�֬A*�ٿ�#z}��@ �L�4@h'-Ӊ�!?2pob�@�֬A*�ٿ�#z}��@ �L�4@h'-Ӊ�!?2pob�@�֬A*�ٿ�#z}��@ �L�4@h'-Ӊ�!?2pob�@�֬A*�ٿ�#z}��@ �L�4@h'-Ӊ�!?2pob�@�t��c�ٿuY&C��@<�����3@K�n;T�!?l c���@�t��c�ٿuY&C��@<�����3@K�n;T�!?l c���@�t��c�ٿuY&C��@<�����3@K�n;T�!?l c���@�t��c�ٿuY&C��@<�����3@K�n;T�!?l c���@P��zբٿ�����Y�@�}n��*4@��+|��!?:�ɀ���@P��zբٿ�����Y�@�}n��*4@��+|��!?:�ɀ���@P��zբٿ�����Y�@�}n��*4@��+|��!?:�ɀ���@P��zբٿ�����Y�@�}n��*4@��+|��!?:�ɀ���@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���l�ٿl��O��@�T����3@l~�7q�!?	�J����@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@���סٿ����Q��@�� 4@����C�!?&:��y�@�#��̡ٿ�CB�\�@ɧ���3@c�a�!?�.k����@�#��̡ٿ�CB�\�@ɧ���3@c�a�!?�.k����@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@sSy���ٿ��ΰ��@�Vb�w&4@}����!?��݃�J�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�S7ݚٿ�:#3�@k�B��3@��>��!?�,�Ǭ�@�j�$�ٿ�	?�t�@	�2��4@ϲJ�ݐ!?D��0�ؕ@�j�$�ٿ�	?�t�@	�2��4@ϲJ�ݐ!?D��0�ؕ@�j�$�ٿ�	?�t�@	�2��4@ϲJ�ݐ!?D��0�ؕ@�{[�#�ٿ5��j½�@�_�$z�3@~R��i�!?F�upO�@�{[�#�ٿ5��j½�@�_�$z�3@~R��i�!?F�upO�@�{[�#�ٿ5��j½�@�_�$z�3@~R��i�!?F�upO�@�{[�#�ٿ5��j½�@�_�$z�3@~R��i�!?F�upO�@�{[�#�ٿ5��j½�@�_�$z�3@~R��i�!?F�upO�@�����ٿ7q�\�@�@��Rr4@��F�!?t�lf��@TcPc�ٿY�0.��@s֦��3@$�n�G�!?7�엶��@TcPc�ٿY�0.��@s֦��3@$�n�G�!?7�엶��@TcPc�ٿY�0.��@s֦��3@$�n�G�!?7�엶��@D�z�Þٿ�0Gr(�@{l���3@$�EN�!?�R�2�@�N<!b�ٿ�ih�Yn�@},�3@T�����!?��.!ԕ@�N<!b�ٿ�ih�Yn�@},�3@T�����!?��.!ԕ@�Ç�F�ٿ�_Q��=�@c�����3@���$�!?8��R|�@�Ç�F�ٿ�_Q��=�@c�����3@���$�!?8��R|�@i��Рٿ�o�,��@�`d�3@�s}>�!?�df��@)Ӻ�ٿ2A)y��@`2����3@����!?F���ȕ@)Ӻ�ٿ2A)y��@`2����3@����!?F���ȕ@)Ӻ�ٿ2A)y��@`2����3@����!?F���ȕ@)Ӻ�ٿ2A)y��@`2����3@����!?F���ȕ@)Ӻ�ٿ2A)y��@`2����3@����!?F���ȕ@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�dQ�ٿi��o�@��`�C�3@���!?��j=L��@�
����ٿvD�/�@���r�/4@�û�,�!?���4e��@�
����ٿvD�/�@���r�/4@�û�,�!?���4e��@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@?G&"��ٿ-F�iU��@v���4@���!Z�!?-�dA�ŕ@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@	Қ�U�ٿ�!a��F�@�R����3@�Z2��!?1�%�#�@Q�Q���ٿ-�&٥	�@,>���3@X����!?ſ$8��@Q�Q���ٿ-�&٥	�@,>���3@X����!?ſ$8��@��$!Q�ٿl�e�0�@X�KL,4@�3�J�!?喝�+�@��$!Q�ٿl�e�0�@X�KL,4@�3�J�!?喝�+�@�K�~�ٿ ��;�@�O�̟4@�8�=Q�!?7U����@�K�~�ٿ ��;�@�O�̟4@�8�=Q�!?7U����@�K�~�ٿ ��;�@�O�̟4@�8�=Q�!?7U����@����S�ٿ�.����@wo�4@~uWZ�!?� ��n(�@����S�ٿ�.����@wo�4@~uWZ�!?� ��n(�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@-����ٿ��#ɴ��@�lSn4@5@�ώ�!?��ml�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@ڪo��ٿ֫�go*�@�Oh�PX4@����Q�!?��,ʕa�@EǔYߞٿ^W?���@��� Y4@����!?��"XG�@EǔYߞٿ^W?���@��� Y4@����!?��"XG�@EǔYߞٿ^W?���@��� Y4@����!?��"XG�@EǔYߞٿ^W?���@��� Y4@����!?��"XG�@"��FJ�ٿh��R� �@Ge�'wK4@'b���!?lj
RG��@"��FJ�ٿh��R� �@Ge�'wK4@'b���!?lj
RG��@ML�p.�ٿ̯���@��D"n4@�_�N��!?SLbƖ�@ML�p.�ٿ̯���@��D"n4@�_�N��!?SLbƖ�@ML�p.�ٿ̯���@��D"n4@�_�N��!?SLbƖ�@ML�p.�ٿ̯���@��D"n4@�_�N��!?SLbƖ�@ ���R�ٿU��l�@ف�4@W=ƴ�!?Eo�S$ޕ@ؒę�ٿ�;Y��r�@�S_O34@i���!?��z����@ؒę�ٿ�;Y��r�@�S_O34@i���!?��z����@ؒę�ٿ�;Y��r�@�S_O34@i���!?��z����@D�����ٿ4<Fƞn�@��r�<4@b�Q�!?�
ہ˙�@D�����ٿ4<Fƞn�@��r�<4@b�Q�!?�
ہ˙�@l��Ϡٿ����r�@�OB��3@Ƌ]�o�!?��"�:�@l��Ϡٿ����r�@�OB��3@Ƌ]�o�!?��"�:�@l��Ϡٿ����r�@�OB��3@Ƌ]�o�!?��"�:�@l��Ϡٿ����r�@�OB��3@Ƌ]�o�!?��"�:�@l��Ϡٿ����r�@�OB��3@Ƌ]�o�!?��"�:�@N���ٿMSz����@�z�@!4@hVJo�!?��ù9�@N���ٿMSz����@�z�@!4@hVJo�!?��ù9�@N���ٿMSz����@�z�@!4@hVJo�!?��ù9�@���!W�ٿ�.�ކ�@{[*4@i�\ʸ�!?�ԉ��_�@���!W�ٿ�.�ކ�@{[*4@i�\ʸ�!?�ԉ��_�@4�b��ٿ�*ϋ���@��ݝ�4@�
(i��!?����ޕ@4�b��ٿ�*ϋ���@��ݝ�4@�
(i��!?����ޕ@j��Þٿ���T�@�z�4@[�����!?G��-�Օ@j��Þٿ���T�@�z�4@[�����!?G��-�Օ@j��Þٿ���T�@�z�4@[�����!?G��-�Օ@%!��ٿhg/�a�@��I�4@Т"�ǐ!?���Ez��@������ٿR��B>�@���U64@��>���!?��;���@������ٿR��B>�@���U64@��>���!?��;���@������ٿR��B>�@���U64@��>���!?��;���@E��ٔ�ٿ�������@u�,�}P4@�!/U��!?����@E��ٔ�ٿ�������@u�,�}P4@�!/U��!?����@bEzs�ٿ8��IF�@i
x�Ua4@��%��!?x��%��@bEzs�ٿ8��IF�@i
x�Ua4@��%��!?x��%��@bEzs�ٿ8��IF�@i
x�Ua4@��%��!?x��%��@�e��ٿ�p���e�@r_�FL4@��-"�!?��8��@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@���&ϖٿDl�ս��@�+�GId4@ �J�!?����+ �@�J�1)�ٿE�J���@�%�� 4@�٘�!?�#�3ٕ@��;;��ٿhn*E���@�zZ��`4@ڨt�Y�!?p���W�@��;;��ٿhn*E���@�zZ��`4@ڨt�Y�!?p���W�@?���u�ٿ�y�)F�@�JDk�h4@�RW��!?��q ��@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@��
Fk�ٿ��Q1�2�@W�_-�3@vi8H6�!?CL�yRl�@�yD�ٿ浆�{�@3�:�:�3@���7�!?m&����@�yD�ٿ浆�{�@3�:�:�3@���7�!?m&����@�yD�ٿ浆�{�@3�:�:�3@���7�!?m&����@�yD�ٿ浆�{�@3�:�:�3@���7�!?m&����@r>o*�ٿ������@�݀G�!4@�d���!?�vs�@r>o*�ٿ������@�݀G�!4@�d���!?�vs�@�k��ٿ�Dn ��@JS�4@��D��!?p�����@�k��ٿ�Dn ��@JS�4@��D��!?p�����@�k��ٿ�Dn ��@JS�4@��D��!?p�����@�{�e��ٿ'�<��@M���3@[�ݽ(�!?L�L���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@����ŜٿX?+i��@�Wxq�4@�Tmv�!?��*���@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@.�'�E�ٿZ$� gB�@���4�4@��˲%�!?������@����ٿ3��w��@�kM��64@5RB�!?��7�_#�@����ٿ3��w��@�kM��64@5RB�!?��7�_#�@�5��ٿå҉*�@�}�+�24@i�ꂐ!?���UE�@�5��ٿå҉*�@�}�+�24@i�ꂐ!?���UE�@$;��ٿ���Y��@N�ji
4@a����!?��R���@$;��ٿ���Y��@N�ji
4@a����!?��R���@$;��ٿ���Y��@N�ji
4@a����!?��R���@�T�ޘٿ�ʊ!�M�@�i4@7FB^�!?`��C��@�T�ޘٿ�ʊ!�M�@�i4@7FB^�!?`��C��@�T�ޘٿ�ʊ!�M�@�i4@7FB^�!?`��C��@����ٿg��AD0�@��x�K4@e����!?X��@����ٿg��AD0�@��x�K4@e����!?X��@����ٿg��AD0�@��x�K4@e����!?X��@�*o|�ٿ��)��T�@et��3@N;�ߛ�!?|�ꏋ��@�*o|�ٿ��)��T�@et��3@N;�ߛ�!?|�ꏋ��@�ZеL�ٿ=�z�{�@wo� ��3@���՛�!?�Ũ��ѕ@�ZеL�ٿ=�z�{�@wo� ��3@���՛�!?�Ũ��ѕ@�ZеL�ٿ=�z�{�@wo� ��3@���՛�!?�Ũ��ѕ@�Lq'X�ٿF-}U��@8��4@���刐!?Xf�ꘕ@�K���ٿi�AR�@ĳn��c4@�g��P�!?;����@�K���ٿi�AR�@ĳn��c4@�g��P�!?;����@KûV�ٿ��t�3��@�?Tk4@��̃g�!?��d���@KûV�ٿ��t�3��@�?Tk4@��̃g�!?��d���@KûV�ٿ��t�3��@�?Tk4@��̃g�!?��d���@b�̲��ٿ������@�����4@`��G�!?��J[��@b�̲��ٿ������@�����4@`��G�!?��J[��@b�̲��ٿ������@�����4@`��G�!?��J[��@b�̲��ٿ������@�����4@`��G�!?��J[��@b�̲��ٿ������@�����4@`��G�!?��J[��@g��IU�ٿɦ0P�@�0�64@����[�!?\��	��@g��IU�ٿɦ0P�@�0�64@����[�!?\��	��@�E�,+�ٿ�~�!�@�&�%�)4@���I�!?&n��o�@�E�,+�ٿ�~�!�@�&�%�)4@���I�!?&n��o�@�E�,+�ٿ�~�!�@�&�%�)4@���I�!?&n��o�@�E�,+�ٿ�~�!�@�&�%�)4@���I�!?&n��o�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�F�ٿ��W�}0�@���K4@9%��!?���UP�@�ɕ:b�ٿ���w5K�@�r{Om�3@�|��0�!?`�m��W�@�Բ���ٿ������@nh��4@T�&�z�!?)ֿ����@�Բ���ٿ������@nh��4@T�&�z�!?)ֿ����@�Բ���ٿ������@nh��4@T�&�z�!?)ֿ����@�Բ���ٿ������@nh��4@T�&�z�!?)ֿ����@�Բ���ٿ������@nh��4@T�&�z�!?)ֿ����@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@HwЬ��ٿ��b��t�@j�A94@��_���!?t���E�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@ӧ��ڛٿ|���Y�@1w�>��3@��ā��!?�6��(�@������ٿ.J��N��@m4�ת�3@a�h_x�!?��}��@^�0=M�ٿ�Շj��@q�d��"4@��#�w�!?�"?�@^�0=M�ٿ�Շj��@q�d��"4@��#�w�!?�"?�@;���=�ٿ���|71�@&�?4@��¯�!?Z���	ϕ@;���=�ٿ���|71�@&�?4@��¯�!?Z���	ϕ@;���=�ٿ���|71�@&�?4@��¯�!?Z���	ϕ@;���=�ٿ���|71�@&�?4@��¯�!?Z���	ϕ@���q̛ٿ�`s���@���l�A4@��/ɳ�!?ɱ-��@���q̛ٿ�`s���@���l�A4@��/ɳ�!?ɱ-��@�T~gݛٿ�vjy��@�s�s.4@�q7���!?��r�@�T~gݛٿ�vjy��@�s�s.4@�q7���!?��r�@�T~gݛٿ�vjy��@�s�s.4@�q7���!?��r�@�T~gݛٿ�vjy��@�s�s.4@�q7���!?��r�@�T~gݛٿ�vjy��@�s�s.4@�q7���!?��r�@F�:�ٿ�hY8M�@��3�EP4@���q�!?;��I���@F�:�ٿ�hY8M�@��3�EP4@���q�!?;��I���@+)���ٿ�'��@�2���=4@	AX��!?����ە@+)���ٿ�'��@�2���=4@	AX��!?����ە@+)���ٿ�'��@�2���=4@	AX��!?����ە@�,3ߤٿB����@G�����3@�
QD6�!?�mM٤�@�,3ߤٿB����@G�����3@�
QD6�!?�mM٤�@�,3ߤٿB����@G�����3@�
QD6�!?�mM٤�@���i%�ٿ�h~�U��@�q#]�$4@�F �!?����ھ�@���i%�ٿ�h~�U��@�q#]�$4@�F �!?����ھ�@���i%�ٿ�h~�U��@�q#]�$4@�F �!?����ھ�@���i%�ٿ�h~�U��@�q#]�$4@�F �!?����ھ�@���i%�ٿ�h~�U��@�q#]�$4@�F �!?����ھ�@!2��ٿ�O1��:�@��b4@�i�{��!?��l���@!2��ٿ�O1��:�@��b4@�i�{��!?��l���@��9t�ٿ-Y� :�@E�!h��3@u{w]��!?���/`�@��9t�ٿ-Y� :�@E�!h��3@u{w]��!?���/`�@��9t�ٿ-Y� :�@E�!h��3@u{w]��!?���/`�@^d�ܻ�ٿbS�,�@�@H1��*4@���Ő!?c9�Ak�@^d�ܻ�ٿbS�,�@�@H1��*4@���Ő!?c9�Ak�@����ٿz��e�@�(��S4@Fa�q��!?ǛǾ��@Ttaܦٿ�?�B��@�ɰ��3@oS�h�!?�Ix���@Ttaܦٿ�?�B��@�ɰ��3@oS�h�!?�Ix���@Ttaܦٿ�?�B��@�ɰ��3@oS�h�!?�Ix���@�2���ٿ�ܫ�]U�@����d�3@>�R8:�!?� �[��@�2���ٿ�ܫ�]U�@����d�3@>�R8:�!?� �[��@�2���ٿ�ܫ�]U�@����d�3@>�R8:�!?� �[��@�2���ٿ�ܫ�]U�@����d�3@>�R8:�!?� �[��@�2���ٿ�ܫ�]U�@����d�3@>�R8:�!?� �[��@�e=_s�ٿ'�Sq���@.�f�&�3@��7h�!?[q�@���ST�ٿӭ�3�@�=m��3@��
1�!?��. ��@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@-t���ٿcj���@d���]4@m�[}�!?hg��+5�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�߈Πٿ���o�@�B���*4@/�]�R�!?���+�@�)ι	�ٿ��f���@M�ܲ�4@)؀F��!?��Q�@�)ι	�ٿ��f���@M�ܲ�4@)؀F��!?��Q�@�ir���ٿ��u:�@\X��iL4@���]�!?���+d��@�ir���ٿ��u:�@\X��iL4@���]�!?���+d��@�ir���ٿ��u:�@\X��iL4@���]�!?���+d��@�ir���ٿ��u:�@\X��iL4@���]�!?���+d��@�ir���ٿ��u:�@\X��iL4@���]�!?���+d��@����ٿ�,���@&�w�,4@_ �JW�!?���7�|�@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�0R<<�ٿ�"^��J�@$�$4@��*?�!?��:!]��@�])�L�ٿ��L�P�@�%���4@�g����!?�	M���@�])�L�ٿ��L�P�@�%���4@�g����!?�	M���@�Us롞ٿE+���@����4@�a�6�!?Mu� F�@�Us롞ٿE+���@����4@�a�6�!?Mu� F�@�Us롞ٿE+���@����4@�a�6�!?Mu� F�@��p��ٿ�G"��v�@g�L�E84@��p�!?�0F���@��p��ٿ�G"��v�@g�L�E84@��p�!?�0F���@��p��ٿ�G"��v�@g�L�E84@��p�!?�0F���@������ٿ�sS���@�-��4@%�m��!?�����ɕ@������ٿ�sS���@�-��4@%�m��!?�����ɕ@������ٿ�sS���@�-��4@%�m��!?�����ɕ@������ٿ�sS���@�-��4@%�m��!?�����ɕ@������ٿ�sS���@�-��4@%�m��!?�����ɕ@� ��ٿ�=r��t�@Xn?l�;4@��f�!?�����@� ��ٿ�=r��t�@Xn?l�;4@��f�!?�����@�^��ٿ⹧�=�@��T~xS4@�:��q�!?�?�.vѕ@�^��ٿ⹧�=�@��T~xS4@�:��q�!?�?�.vѕ@�^��ٿ⹧�=�@��T~xS4@�:��q�!?�?�.vѕ@�^��ٿ⹧�=�@��T~xS4@�:��q�!?�?�.vѕ@���ً�ٿ��r��6�@V�F4@9t�"�!?�^�^���@;hw��ٿ��m��@��/�94@���X�!?tԎ�c�@;hw��ٿ��m��@��/�94@���X�!?tԎ�c�@����ٿ�p�>��@��D�E4@��I�!?���$��@����ٿ�p�>��@��D�E4@��I�!?���$��@�5 �$�ٿ���b�@~CYD�b4@����^�!?Td���R�@4�Aޡٿi6�;7��@F�t�3@(���ѐ!?����@�*����ٿ)�8�@���\7�3@qj�ؐ!?����ٕ@�*����ٿ)�8�@���\7�3@qj�ؐ!?����ٕ@_ 0��ٿ����R�@��|�U�3@y�cܐ!?Y�o�B�@_ 0��ٿ����R�@��|�U�3@y�cܐ!?Y�o�B�@_ 0��ٿ����R�@��|�U�3@y�cܐ!?Y�o�B�@��OES�ٿ�@�ce�@-'�/��3@pi��ΐ!?>�S���@/�9��ٿ�7�e��@��@�3@�����!?��kޣ�@�Y։�ٿ~�9>�{�@�o�G�3@2V�p�!?�]W�=��@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@�z�H�ٿ�V��a�@�|��4@k�%�!?�j0���@n�U��ٿl�}6�R�@��ZP<4@�b��!?����ň�@n�U��ٿl�}6�R�@��ZP<4@�b��!?����ň�@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@��褂�ٿ���c��@ܸ�b4@F)3Ɛ!?�[?����@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@)���Z�ٿ�*��@�F0�'4@}�T@E�!?���񽩕@�QQ�ٿh��u�@qi��(4@:2�Ǉ�!?���9�@�QQ�ٿh��u�@qi��(4@:2�Ǉ�!?���9�@�QQ�ٿh��u�@qi��(4@:2�Ǉ�!?���9�@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@�f����ٿF�&�m�@kg�z�4@��.�J�!?1�f���@c����ٿ/�j�1��@g'4@@E�#1�!?��&���@c����ٿ/�j�1��@g'4@@E�#1�!?��&���@c����ٿ/�j�1��@g'4@@E�#1�!?��&���@c����ٿ/�j�1��@g'4@@E�#1�!?��&���@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@/��P�ٿ���!��@���B4@Ǹ��[�!?wAt�鹕@_�נ#�ٿ��e$Zn�@;1J>4@ˆ��4�!?[:�%��@_�נ#�ٿ��e$Zn�@;1J>4@ˆ��4�!?[:�%��@_�נ#�ٿ��e$Zn�@;1J>4@ˆ��4�!?[:�%��@_�נ#�ٿ��e$Zn�@;1J>4@ˆ��4�!?[:�%��@_�נ#�ٿ��e$Zn�@;1J>4@ˆ��4�!?[:�%��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@����6�ٿ������@Rn	նC4@G�G�a�!?��(s��@܆n�ٿ�����)�@����04@��jڜ�!?&��J�@܆n�ٿ�����)�@����04@��jڜ�!?&��J�@܆n�ٿ�����)�@����04@��jڜ�!?&��J�@܆n�ٿ�����)�@����04@��jڜ�!?&��J�@܆n�ٿ�����)�@����04@��jڜ�!?&��J�@
�A줞ٿg}���@���u�4@,��s`�!?m>��]�@
�A줞ٿg}���@���u�4@,��s`�!?m>��]�@
�A줞ٿg}���@���u�4@,��s`�!?m>��]�@
�A줞ٿg}���@���u�4@,��s`�!?m>��]�@�2/c��ٿ�#):��@�*�
4@�c���!?���9��@�2/c��ٿ�#):��@�*�
4@�c���!?���9��@�2/c��ٿ�#):��@�*�
4@�c���!?���9��@�2/c��ٿ�#):��@�*�
4@�c���!?���9��@���gۣٿ��Q�	�@ ��4@�S��;�!?�� �dw�@M�%��ٿ�}���@����_$4@���/�!?���v�@M�%��ٿ�}���@����_$4@���/�!?���v�@M�%��ٿ�}���@����_$4@���/�!?���v�@M�%��ٿ�}���@����_$4@���/�!?���v�@M�%��ٿ�}���@����_$4@���/�!?���v�@M�%��ٿ�}���@����_$4@���/�!?���v�@��>hҠٿ��C���@Q�k�4@��b�0�!?S�Xr��@�D�n"�ٿ��_.��@�B�4@�@)��!?��O��@�D�n"�ٿ��_.��@�B�4@�@)��!?��O��@�D�n"�ٿ��_.��@�B�4@�@)��!?��O��@�D�n"�ٿ��_.��@�B�4@�@)��!?��O��@�D�n"�ٿ��_.��@�B�4@�@)��!?��O��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@K����ٿ���U��@�c��4@�]���!?�3%#��@=, ��ٿr��8��@IX��:�3@
���5�!?Z�^ǝ��@=, ��ٿr��8��@IX��:�3@
���5�!?Z�^ǝ��@=, ��ٿr��8��@IX��:�3@
���5�!?Z�^ǝ��@��d���ٿ�繪Lc�@s�+S4@��I�!?u��u�@��d���ٿ�繪Lc�@s�+S4@��I�!?u��u�@��d���ٿ�繪Lc�@s�+S4@��I�!?u��u�@�4W��ٿ�w]%��@ͨ|d�3@�Q�_S�!??���?�@�4W��ٿ�w]%��@ͨ|d�3@�Q�_S�!??���?�@�4W��ٿ�w]%��@ͨ|d�3@�Q�_S�!??���?�@�4W��ٿ�w]%��@ͨ|d�3@�Q�_S�!??���?�@�4��ٿ0�Ze�Q�@8ᱱ��3@���w�!?�u�<�@�4��ٿ0�Ze�Q�@8ᱱ��3@���w�!?�u�<�@�4��ٿ0�Ze�Q�@8ᱱ��3@���w�!?�u�<�@05T���ٿr}���,�@�R�ߏ4@�Wջ�!?�����@��ӳm�ٿ���V3�@��x��3@��Yɾ�!?`W�2i��@�p�7�ٿ���<��@�g�3@\��e�!?^)��8�@�p�7�ٿ���<��@�g�3@\��e�!?^)��8�@�p�7�ٿ���<��@�g�3@\��e�!?^)��8�@�/��ܜٿ���+0�@�����3@�R�G�!?����.�@�/��ܜٿ���+0�@�����3@�R�G�!?����.�@�/��ܜٿ���+0�@�����3@�R�G�!?����.�@�/��ܜٿ���+0�@�����3@�R�G�!?����.�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@P�G,��ٿ]�I����@ۍf���3@ �z�z�!?�j�)�A�@{ӱ�O�ٿ�����@�r~*�3@�^Ǥ�!?O����@{ӱ�O�ٿ�����@�r~*�3@�^Ǥ�!?O����@{ӱ�O�ٿ�����@�r~*�3@�^Ǥ�!?O����@�o\�B�ٿ���x��@�BNb4@)��ک�!?L|��� �@G���M�ٿ*`Ud��@��&4@xX�6��!?G����@Bɔ�ٿ&.�;�@��0u<4@��~��!?���P�&�@Bɔ�ٿ&.�;�@��0u<4@��~��!?���P�&�@C��Y�ٿ������@��
�T4@���Đ!?E��s���@C��Y�ٿ������@��
�T4@���Đ!?E��s���@�i$�\�ٿC�	�@��Ü4@-6��!?��8��ϕ@�i$�\�ٿC�	�@��Ü4@-6��!?��8��ϕ@�i$�\�ٿC�	�@��Ü4@-6��!?��8��ϕ@�i$�\�ٿC�	�@��Ü4@-6��!?��8��ϕ@2O�W��ٿlu ��p�@O�z�t'4@A\��:�!?f�U'L�@2O�W��ٿlu ��p�@O�z�t'4@A\��:�!?f�U'L�@2O�W��ٿlu ��p�@O�z�t'4@A\��:�!?f�U'L�@2O�W��ٿlu ��p�@O�z�t'4@A\��:�!?f�U'L�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@_�:[�ٿNm`ХC�@�+}n^4@,�3鉐!?�cC�ـ�@OǱ1��ٿ�G�K�@(���oB4@ȀfA�!?T�f�@����ٿ��T
l�@ �KɄ%4@7:q\�!?�͂"��@���@�ٿ���?��@���-4@L��&�!?��<-��@���@�ٿ���?��@���-4@L��&�!?��<-��@���@�ٿ���?��@���-4@L��&�!?��<-��@i)�9ӟٿY�UhNO�@��$���3@b:���!?��Yt��@AH`�v�ٿ��1����@Eͥx�4@��<�#�!?�G{ȕ@AH`�v�ٿ��1����@Eͥx�4@��<�#�!?�G{ȕ@AH`�v�ٿ��1����@Eͥx�4@��<�#�!?�G{ȕ@�6��ٿO,C?|�@���C4@���!?�1��f�@�6��ٿO,C?|�@���C4@���!?�1��f�@�6��ٿO,C?|�@���C4@���!?�1��f�@�6��ٿO,C?|�@���C4@���!?�1��f�@��>\�ٿ:gV��1�@@� I�3@����!?nK�|Ͽ�@��>\�ٿ:gV��1�@@� I�3@����!?nK�|Ͽ�@��>\�ٿ:gV��1�@@� I�3@����!?nK�|Ͽ�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@��J��ٿzz��5*�@���n�3@�6l�!?�S*��/�@���l�ٿ�{"�z�@��194@��Y=�!?��W�@���l�ٿ�{"�z�@��194@��Y=�!?��W�@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@��W�7�ٿ������@��U�d-4@(z\u�!?��J�ޕ@�4��?�ٿb!�H��@��^B.4@��B��!?j�e��7�@d[,�ٿ׫�@F3�k�4@2�2�f�!?]��Y�W�@d[,�ٿ׫�@F3�k�4@2�2�f�!?]��Y�W�@TB좛ٿV7�y�j�@���Y4@�񮒐!?��Z��@TB좛ٿV7�y�j�@���Y4@�񮒐!?��Z��@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@�@gs��ٿ��4��@�M���-4@4c7���!?���I�@��E�ٿ#NSX���@AD�]�84@)+�H�!?+�/��@��E�ٿ#NSX���@AD�]�84@)+�H�!?+�/��@��E�ٿ#NSX���@AD�]�84@)+�H�!?+�/��@��E�ٿ#NSX���@AD�]�84@)+�H�!?+�/��@lp��b�ٿ^Y���A�@	�m��B4@5�[i�!?���q�?�@lp��b�ٿ^Y���A�@	�m��B4@5�[i�!?���q�?�@lp��b�ٿ^Y���A�@	�m��B4@5�[i�!?���q�?�@lp��b�ٿ^Y���A�@	�m��B4@5�[i�!?���q�?�@��M���ٿrL6�q�@E�.�4@�^��;�!?Q-V�]�@��)b��ٿ�y[ij��@�h�l4@Umg9�!?ݻ��w�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@�.��ٿ�_78/d�@�l\��4@�A*$f�!?u�2�N�@j����ٿCMc���@l�l0�4@�R�!?��q�@Y�}q�ٿ8SN���@��4*4@�Џ{K�!?���VV�@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@�ЄOo�ٿ�2</��@���F�3@۱�<l�!?����@��L�ٿT�z/v�@-�ZU#4@0!���!?�S~��@Qa%��ٿI���&�@W�b�,4@0Bu�؏!?ݹ��ԍ�@|��D�ٿ�G	H��@)a�[@4@�I��!?{o36��@|��D�ٿ�G	H��@)a�[@4@�I��!?{o36��@|��D�ٿ�G	H��@)a�[@4@�I��!?{o36��@|��D�ٿ�G	H��@)a�[@4@�I��!?{o36��@%��H�ٿ�/Yf2��@ ���$4@ۀxm��!?�(a�@%��H�ٿ�/Yf2��@ ���$4@ۀxm��!?�(a�@%��H�ٿ�/Yf2��@ ���$4@ۀxm��!?�(a�@%��H�ٿ�/Yf2��@ ���$4@ۀxm��!?�(a�@%��H�ٿ�/Yf2��@ ���$4@ۀxm��!?�(a�@WY��ٿ����[�@��,804@o4����!?��#�<�@WY��ٿ����[�@��,804@o4����!?��#�<�@WY��ٿ����[�@��,804@o4����!?��#�<�@WY��ٿ����[�@��,804@o4����!?��#�<�@WY��ٿ����[�@��,804@o4����!?��#�<�@�ҧ��ٿ���E��@"fA�m>4@C.���!?��y�걕@x4��,�ٿ�m�^�@}���4@v܂hs�!?�3�~��@x4��,�ٿ�m�^�@}���4@v܂hs�!?�3�~��@x4��,�ٿ�m�^�@}���4@v܂hs�!?�3�~��@x4��,�ٿ�m�^�@}���4@v܂hs�!?�3�~��@֒��@�ٿP�$;<�@�J�W+4@�+Ts�!?��~��֕@֒��@�ٿP�$;<�@�J�W+4@�+Ts�!?��~��֕@֒��@�ٿP�$;<�@�J�W+4@�+Ts�!?��~��֕@֒��@�ٿP�$;<�@�J�W+4@�+Ts�!?��~��֕@֒��@�ٿP�$;<�@�J�W+4@�+Ts�!?��~��֕@���A	�ٿ����7�@���5h%4@Ct|L�!?W��V�@���A	�ٿ����7�@���5h%4@Ct|L�!?W��V�@���A	�ٿ����7�@���5h%4@Ct|L�!?W��V�@���A	�ٿ����7�@���5h%4@Ct|L�!?W��V�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@V�j2�ٿ��H����@�;�4@S��K��!?��.j�@�
��Ϝٿ�e���@3a�VV4@M{hF�!?�����˕@�
��Ϝٿ�e���@3a�VV4@M{hF�!?�����˕@�
��Ϝٿ�e���@3a�VV4@M{hF�!?�����˕@�
��Ϝٿ�e���@3a�VV4@M{hF�!?�����˕@�
��Ϝٿ�e���@3a�VV4@M{hF�!?�����˕@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@|:�ƍ�ٿ$󂈀�@�:}4@��`�!?�O3���@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@��V�ٿ�<�NX��@������3@��8���!?��!�@S�l�ٿy�E}|��@Y&S�i�3@�	m	<�!?=Y��;ȕ@��0�|�ٿ(����`�@<�T~�3@���X�!?�E��0�@-"�w�ٿ����2�@q���c�3@m��b�!?�g�%�\�@-"�w�ٿ����2�@q���c�3@m��b�!?�g�%�\�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@���4�ٿ����@�Z�»3@�t�!h�!?(/M�W�@��X6�ٿs���@PPGe�3@�u��:�!?����gZ�@�& '�ٿ ^pH��@be��g�3@Q
<�_�!?9�i/�q�@�^��ٿ� �Tܶ�@�ϢS�+4@nY �!?\����
�@��}al�ٿ��x+j�@m����4@V${�!?��"?'�@��}al�ٿ��x+j�@m����4@V${�!?��"?'�@��}al�ٿ��x+j�@m����4@V${�!?��"?'�@��}al�ٿ��x+j�@m����4@V${�!?��"?'�@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@*�&[O�ٿ�0�(���@)��΂;4@��
N�!?A����ݕ@��t�T�ٿ,��^��@V��_d�3@��xZ�!?�*�n�0�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@mL��H�ٿ�����@����3@�9�!?�HM-A�@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@���g��ٿ�� ʱ�@o�6j�3@����!?�7y���@�٣�ߣٿ7�=g@0�@�`��4@����)�!?^�\��c�@�٣�ߣٿ7�=g@0�@�`��4@����)�!?^�\��c�@�m!}�ٿ��i7��@��-Z��3@�1�8�!?��w�(�@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@
��ڡٿ�C8`��@�:�?h,4@}H�( �!?.li�ĕ@�����ٿ
5{,��@�����4@���-e�!?< �B�@�����ٿ
5{,��@�����4@���-e�!?< �B�@�����ٿ
5{,��@�����4@���-e�!?< �B�@�����ٿ
5{,��@�����4@���-e�!?< �B�@Α���ٿ/�q�e�@���J34@W�]�~�!?7�2�wc�@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@b|a6�ٿj���Z��@��k#4@���p@�!?�t�#��@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@���YC�ٿ(�! NC�@٣�(�4@ϙs�H�!??�G����@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@	q��ٿ�S��_��@ss�|� 4@#c�;�!?^��pݕ@1V��"�ٿ��kB�@�_�N~4@��r�%�!?�YB��@1V��"�ٿ��kB�@�_�N~4@��r�%�!?�YB��@1V��"�ٿ��kB�@�_�N~4@��r�%�!?�YB��@1V��"�ٿ��kB�@�_�N~4@��r�%�!?�YB��@��P��ٿ)��g��@U��U$4@���F�!?ܳI\d�@m� s�ٿ���5ܵ�@V�(�&4@�+g�!?W@	4��@m� s�ٿ���5ܵ�@V�(�&4@�+g�!?W@	4��@m� s�ٿ���5ܵ�@V�(�&4@�+g�!?W@	4��@V}ᨠٿ���O��@�ڦ�R
4@��.�n�!?�O���K�@V}ᨠٿ���O��@�ڦ�R
4@��.�n�!?�O���K�@�*Zv�ٿ�X�*ӎ�@sϸʁ 4@����!?�N7���@�*Zv�ٿ�X�*ӎ�@sϸʁ 4@����!?�N7���@�*Zv�ٿ�X�*ӎ�@sϸʁ 4@����!?�N7���@+���]�ٿS���@sЕ��,4@$�~�{�!?�ӗɢ�@+���]�ٿS���@sЕ��,4@$�~�{�!?�ӗɢ�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@Y��ٿsP;P���@�⫱�44@.̰<�!?���Q}�@���6�ٿ��,_��@�x_�A4@W��#�!?	a�T�@���6�ٿ��,_��@�x_�A4@W��#�!?	a�T�@l.���ٿ�7	�_��@YG��I4@��/"c�!?�72)$)�@�����ٿ9�����@�ý]:X4@1�׼p�!?£K����@�����ٿ9�����@�ý]:X4@1�׼p�!?£K����@��JtÜٿ	�}V���@,Ǻ��4@�^��!?�+��ە@��JtÜٿ	�}V���@,Ǻ��4@�^��!?�+��ە@��JtÜٿ	�}V���@,Ǻ��4@�^��!?�+��ە@]Q��ٿz�7�D��@�N_�*+4@g�,��!?6�xF�@]Q��ٿz�7�D��@�N_�*+4@g�,��!?6�xF�@]Q��ٿz�7�D��@�N_�*+4@g�,��!?6�xF�@j�a���ٿ�36��@�C�R�4@�j��^�!?{{��D-�@j�a���ٿ�36��@�C�R�4@�j��^�!?{{��D-�@j�a���ٿ�36��@�C�R�4@�j��^�!?{{��D-�@j�a���ٿ�36��@�C�R�4@�j��^�!?{{��D-�@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@���Ԙٿ@ ����@�����84@��lFT�!?��^��@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@wH�/}�ٿ}l�K+�@�S��4@\*��!?{,�eە@Zk��ٿ�v�E���@�4Z�E4@���z�!?����X�@Zk��ٿ�v�E���@�4Z�E4@���z�!?����X�@Zk��ٿ�v�E���@�4Z�E4@���z�!?����X�@Zk��ٿ�v�E���@�4Z�E4@���z�!?����X�@Zk��ٿ�v�E���@�4Z�E4@���z�!?����X�@�i��ٿx���@���m,�3@gH*�{�!?;�4��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@
���ٿ�]����@n�a+�4@O�Fz�!?��a�A��@<��e�ٿ��F���@<<|��3@��N`�!?^|֜���@<��e�ٿ��F���@<<|��3@��N`�!?^|֜���@<��e�ٿ��F���@<<|��3@��N`�!?^|֜���@�q���ٿ��q����@�Zy�4@n�;�b�!?|�PVP��@�q���ٿ��q����@�Zy�4@n�;�b�!?|�PVP��@�a�Wͪٿ(:`�H��@�ʰ7y!4@���X�!?x,�bډ�@ �M]�ٿ����c�@�/���3@o�q�!?����9�@���>W�ٿ|��B0��@u?o>�4@b�-WC�!?�uc�A�@���>W�ٿ|��B0��@u?o>�4@b�-WC�!?�uc�A�@����ٿ��MH�]�@��K{Ow4@�07�!�!?�1؇l��@����ٿ��MH�]�@��K{Ow4@�07�!�!?�1؇l��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�]�	�ٿxEy"��@��n�&4@�_�C�!?e�f\��@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@�iD��ٿs.��m��@��F��4@���V�!?Ɖ�cł�@��{�h�ٿ)%z��v�@�Aa�4@�B�+�!?����)�@_lޡ.�ٿ�	�5l�@�e�_4@K!`qj�!?W&摌-�@2�4�#�ٿ��J0�F�@�}���4@׾ː!?�t!��@2�4�#�ٿ��J0�F�@�}���4@׾ː!?�t!��@2�4�#�ٿ��J0�F�@�}���4@׾ː!?�t!��@2�4�#�ٿ��J0�F�@�}���4@׾ː!?�t!��@2�4�#�ٿ��J0�F�@�}���4@׾ː!?�t!��@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@%V�NE�ٿ�=o;2��@��BY*#4@��{���!?��@���@q�4�՛ٿ�����@/O�}'-4@f�o�,�!?ejy�!�@q�4�՛ٿ�����@/O�}'-4@f�o�,�!?ejy�!�@q�4�՛ٿ�����@/O�}'-4@f�o�,�!?ejy�!�@q�4�՛ٿ�����@/O�}'-4@f�o�,�!?ejy�!�@\6aΚٿ��}��.�@��14@�B���!?�\�Y~�@zy��D�ٿ0���و�@����R4@'�ͬb�!?�z�/f�@zy��D�ٿ0���و�@����R4@'�ͬb�!?�z�/f�@zy��D�ٿ0���و�@����R4@'�ͬb�!?�z�/f�@�@[�ٿAQ�����@Y6H>m4@p0�)v�!?�.g͑W�@FU�uQ�ٿ��`�I�@|�4�
+4@Y��j�!?_`��fs�@FU�uQ�ٿ��`�I�@|�4�
+4@Y��j�!?_`��fs�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@�Y�2k�ٿ����g�@��mF14@P7B��!?�ڇ�S�@t�U�4�ٿ�"t�ɰ�@�6��$4@����v�!?1������@t�U�4�ٿ�"t�ɰ�@�6��$4@����v�!?1������@t�U�4�ٿ�"t�ɰ�@�6��$4@����v�!?1������@t�U�4�ٿ�"t�ɰ�@�6��$4@����v�!?1������@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@��s�i�ٿ�u�j��@�,mV64@��I�X�!?9H���_�@�lki%�ٿ	�K^��@�D4@s��6�!?N>|���@�lki%�ٿ	�K^��@�D4@s��6�!?N>|���@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��ȱ�ٿN���Hx�@=�$P4@ʍ�Xr�!?���A�@��f�5�ٿ@T��@*�/�� 4@�I�!?���#�'�@��f�5�ٿ@T��@*�/�� 4@�I�!?���#�'�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@�r6�|�ٿ��ZS�@��q�24@.���!?O�Z@$�@O�r���ٿM�h
�z�@�tmo�Q4@=$���!?Ȅ�[�R�@�E3�9�ٿ�jXH� �@�+��54@�����!?�]U�Wؖ@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@��ɕٿޑf��@���)4@���X��!?⻿��1�@/�����ٿBaX�5��@bت�(4@��/��!?ؓEr�)�@xy<%_�ٿw�"�$�@��ŧ@4@q�o/O�!?_�Qٺ&�@xy<%_�ٿw�"�$�@��ŧ@4@q�o/O�!?_�Qٺ&�@����ٿ�MW<���@�F�)4@�1�@�!?��Y2tٖ@OA!FS�ٿ�]��۹�@�##�J4@�Am�?�!?zV�c~�@OA!FS�ٿ�]��۹�@�##�J4@�Am�?�!?zV�c~�@ޛ�ٿ�t,����@ly��E4@@$�H�!?0/���/�@G�
�ٿ2�!����@��%Cf4@�Z�Ð!?��Ǖ@G�
�ٿ2�!����@��%Cf4@�Z�Ð!?��Ǖ@t��)�ٿeD"��p�@43>Kp4@3�	ѐ!?��\@t��)�ٿeD"��p�@43>Kp4@3�	ѐ!?��\@t��)�ٿeD"��p�@43>Kp4@3�	ѐ!?��\@t��)�ٿeD"��p�@43>Kp4@3�	ѐ!?��\@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@��۷ �ٿ�s�	'��@vk�p�k4@e �ِ!?��mPv �@C��C��ٿ-J����@X��č�4@3��[��!?���*�ޕ@C��C��ٿ-J����@X��č�4@3��[��!?���*�ޕ@C��C��ٿ-J����@X��č�4@3��[��!?���*�ޕ@C��C��ٿ-J����@X��č�4@3��[��!?���*�ޕ@C��C��ٿ-J����@X��č�4@3��[��!?���*�ޕ@Y���w�ٿ$b���\�@�)�Q�\4@�E�P\�!?M�R5�@Y���w�ٿ$b���\�@�)�Q�\4@�E�P\�!?M�R5�@Y���w�ٿ$b���\�@�)�Q�\4@�E�P\�!?M�R5�@Y���w�ٿ$b���\�@�)�Q�\4@�E�P\�!?M�R5�@,\��C�ٿb���!�@��ڣ<4@}R��!?C	�γ�@_2����ٿ��N��&�@ +�'&4@���#��!?�Q�H��@_2����ٿ��N��&�@ +�'&4@���#��!?�Q�H��@_2����ٿ��N��&�@ +�'&4@���#��!?�Q�H��@y��H�ٿ���0��@��]�;4@�rPH�!?H�?��n�@i㠛ٿs+���@�SX��4@�����!?��!o��@i㠛ٿs+���@�SX��4@�����!?��!o��@i㠛ٿs+���@�SX��4@�����!?��!o��@i㠛ٿs+���@�SX��4@�����!?��!o��@i㠛ٿs+���@�SX��4@�����!?��!o��@i㠛ٿs+���@�SX��4@�����!?��!o��@�?
8�ٿ^���@��=o[\4@s���z�!?`�8���@����z�ٿ�С��@�K�*�.4@)�h�!?_z.��O�@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@T@�z"�ٿc:��g��@K�?+4@ �Ӥ��!?�T����@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�z�iw�ٿF�d���@����b14@�����!?�6�Si��@�7w �ٿ�[U����@s:�{34@ H{�t�!?S��КV�@�7w �ٿ�[U����@s:�{34@ H{�t�!?S��КV�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@�5���ٿD�,�q��@#?d[4@TrØ��!?V[B�*�@,�!�k�ٿ�]�Aa��@�1��4@���44�!?���D��@,�!�k�ٿ�]�Aa��@�1��4@���44�!?���D��@�WcJ��ٿ���%���@P��/��4@S��t�!?�}��=�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��|��ٿ{k��,5�@_�T=�4@?���S�!?��cbRs�@��4�3�ٿv�#s��@71Q�&�4@���'=�!?D�fM��@��4�3�ٿv�#s��@71Q�&�4@���'=�!?D�fM��@��4�3�ٿv�#s��@71Q�&�4@���'=�!?D�fM��@��4�3�ٿv�#s��@71Q�&�4@���'=�!?D�fM��@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@���X'�ٿY��?��@Q�!�>4@?m��!?�qS�Gȕ@RXl?�ٿ� 'UAl�@D��Đ4@(�,9�!?l�q{�3�@RXl?�ٿ� 'UAl�@D��Đ4@(�,9�!?l�q{�3�@RXl?�ٿ� 'UAl�@D��Đ4@(�,9�!?l�q{�3�@RXl?�ٿ� 'UAl�@D��Đ4@(�,9�!?l�q{�3�@RXl?�ٿ� 'UAl�@D��Đ4@(�,9�!?l�q{�3�@|v�V%�ٿ;^Z.h�@��l"4@fѵ
T�!?��� Q�@��[f�ٿ����@��k�,04@��@�1�!?����T��@��[f�ٿ����@��k�,04@��@�1�!?����T��@�_L�ٿd`��_�@x��)�3@��P��!?@�Xt��@�_L�ٿd`��_�@x��)�3@��P��!?@�Xt��@k�[oƙٿZ�X���@w�	�34@&����!?M:�p��@k�[oƙٿZ�X���@w�	�34@&����!?M:�p��@k�[oƙٿZ�X���@w�	�34@&����!?M:�p��@.`j�9�ٿ6gi�@��}%�N4@��R8y�!?������@.`j�9�ٿ6gi�@��}%�N4@��R8y�!?������@.`j�9�ٿ6gi�@��}%�N4@��R8y�!?������@.`j�9�ٿ6gi�@��}%�N4@��R8y�!?������@Gid���ٿ�wj�J^�@MsHǁ64@�e�=�!?1�z�@xTv���ٿU'�����@��o�/4@Qc����!?��a�ʫ�@xTv���ٿU'�����@��o�/4@Qc����!?��a�ʫ�@xTv���ٿU'�����@��o�/4@Qc����!?��a�ʫ�@xTv���ٿU'�����@��o�/4@Qc����!?��a�ʫ�@xTv���ٿU'�����@��o�/4@Qc����!?��a�ʫ�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��l�g�ٿ �U���@	[plI�3@�]1�!?q�k�@��ɪ�ٿ�88is?�@�&"���3@�d�%�!?��Vѕ@��ɪ�ٿ�88is?�@�&"���3@�d�%�!?��Vѕ@��ɪ�ٿ�88is?�@�&"���3@�d�%�!?��Vѕ@�-�
�ٿm����P�@�iwoM�3@U?�=j�!?��,ԭ��@�-�
�ٿm����P�@�iwoM�3@U?�=j�!?��,ԭ��@�-�
�ٿm����P�@�iwoM�3@U?�=j�!?��,ԭ��@�-�
�ٿm����P�@�iwoM�3@U?�=j�!?��,ԭ��@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@Z�~�ٿ�z�=���@V2s�3@g���R�!?Vi�̵�@C��g�ٿX�E���@�~͠?�3@(ء���!?�D�z��@C��g�ٿX�E���@�~͠?�3@(ء���!?�D�z��@C��g�ٿX�E���@�~͠?�3@(ء���!?�D�z��@C��g�ٿX�E���@�~͠?�3@(ء���!?�D�z��@0*�	�ٿ��ιώ�@i	�AO�3@�����!?�(�����@0*�	�ٿ��ιώ�@i	�AO�3@�����!?�(�����@0*�	�ٿ��ιώ�@i	�AO�3@�����!?�(�����@0*�	�ٿ��ιώ�@i	�AO�3@�����!?�(�����@0*�	�ٿ��ιώ�@i	�AO�3@�����!?�(�����@V��D�ٿ
�2��@�P(�|�3@Dg����!?m���.�@V��D�ٿ
�2��@�P(�|�3@Dg����!?m���.�@V��D�ٿ
�2��@�P(�|�3@Dg����!?m���.�@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@���ǜٿɨ�F�{�@�k���3@!���!?B����Օ@퓯�Ǜٿ��By�
�@��G�k�3@��+l�!?��;s�@퓯�Ǜٿ��By�
�@��G�k�3@��+l�!?��;s�@퓯�Ǜٿ��By�
�@��G�k�3@��+l�!?��;s�@����8�ٿ���+1�@��ũM24@���[P�!?�j����@����8�ٿ���+1�@��ũM24@���[P�!?�j����@����8�ٿ���+1�@��ũM24@���[P�!?�j����@�����ٿ���g�q�@��G�"$4@!�!tI�!?4)a��@�����ٿ���g�q�@��G�"$4@!�!tI�!?4)a��@�����ٿ���g�q�@��G�"$4@!�!tI�!?4)a��@�����ٿ���g�q�@��G�"$4@!�!tI�!?4)a��@���-^�ٿ�I�_��@���8J(4@d ���!?�s����@���-^�ٿ�I�_��@���8J(4@d ���!?�s����@���-^�ٿ�I�_��@���8J(4@d ���!?�s����@-���O�ٿ�[�Jj>�@��N4@3�V�!?���V�P�@-���O�ٿ�[�Jj>�@��N4@3�V�!?���V�P�@-���O�ٿ�[�Jj>�@��N4@3�V�!?���V�P�@-���O�ٿ�[�Jj>�@��N4@3�V�!?���V�P�@-���O�ٿ�[�Jj>�@��N4@3�V�!?���V�P�@�Si׍�ٿ��;}�w�@Z~��>4@��6�Z�!?H�usm�@�I׬s�ٿ�8�"���@��m��3@��[.\�!?jG^��|�@�I׬s�ٿ�8�"���@��m��3@��[.\�!?jG^��|�@�I׬s�ٿ�8�"���@��m��3@��[.\�!?jG^��|�@�I׬s�ٿ�8�"���@��m��3@��[.\�!?jG^��|�@�I׬s�ٿ�8�"���@��m��3@��[.\�!?jG^��|�@ �P��ٿ�[n���@T.��3@FV��d�!?��F�a�@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@%��9(�ٿ��?��@�(=��3@�\'瑐!?��fN��@�9����ٿ���8B��@&-+�3@�]��w�!?�|1�ŕ@�9����ٿ���8B��@&-+�3@�]��w�!?�|1�ŕ@�9����ٿ���8B��@&-+�3@�]��w�!?�|1�ŕ@�9����ٿ���8B��@&-+�3@�]��w�!?�|1�ŕ@�9����ٿ���8B��@&-+�3@�]��w�!?�|1�ŕ@�� ���ٿ��+Q}�@5&�@.�3@Kl��b�!?�N�tm��@�� ���ٿ��+Q}�@5&�@.�3@Kl��b�!?�N�tm��@�� ���ٿ��+Q}�@5&�@.�3@Kl��b�!?�N�tm��@�� ���ٿ��+Q}�@5&�@.�3@Kl��b�!?�N�tm��@�� ���ٿ��+Q}�@5&�@.�3@Kl��b�!?�N�tm��@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@��'�ٿ�Y�2��@�e���3@�^q�`�!?,�g!�@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@@��؞ٿFvк1�@�o��+�3@��5_�!?�-Ǖ@��W��ٿF�ӹ#�@�At�f�3@�G�
Z�!?!ˡk9�@��W��ٿF�ӹ#�@�At�f�3@�G�
Z�!?!ˡk9�@r���ٿ�̷g���@z����S4@� ��!?&Ҁ=B��@r���ٿ�̷g���@z����S4@� ��!?&Ҁ=B��@r���ٿ�̷g���@z����S4@� ��!?&Ҁ=B��@0񲲢ٿ��v��@��Q%p�3@�Y���!?�l��m֕@0񲲢ٿ��v��@��Q%p�3@�Y���!?�l��m֕@.WI��ٿ�tB���@�b���4@��h��!?���U��@.WI��ٿ�tB���@�b���4@��h��!?���U��@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@������ٿ�߯'��@��M"�3@'�V���!?�����Օ@�㺎��ٿ������@<H�Xc94@!G��m�!?���?ו@�e̹�ٿ��I�u�@C�em�34@�L35��!?l=�{��@�e̹�ٿ��I�u�@C�em�34@�L35��!?l=�{��@�e̹�ٿ��I�u�@C�em�34@�L35��!?l=�{��@m&�*ןٿ[��y��@T��e�4@ɇs��!?<��uy�@m&�*ןٿ[��y��@T��e�4@ɇs��!?<��uy�@m&�*ןٿ[��y��@T��e�4@ɇs��!?<��uy�@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@C�~޶�ٿ/+'�|�@�D�C�3@;i�ᩐ!?A��<���@V�*�ٿ\�V����@ˬ��:4@y����!?o ���@�M�ٿ�,�	��@���J5]4@�h�1^�!?�t5��1�@�:�!��ٿ��Z�E��@���M4@!��g�!?j�J7+��@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@v�^��ٿ�4����@��D�@4@�;Y�N�!?���w2�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@c��Y��ٿSۖJ�b�@>n��4@8��h�!?��u��6�@����ʓٿ��RF-�@��E4@��hӐ!?�-n2G�@����ʓٿ��RF-�@��E4@��hӐ!?�-n2G�@����ʓٿ��RF-�@��E4@��hӐ!?�-n2G�@����ʓٿ��RF-�@��E4@��hӐ!?�-n2G�@����ʓٿ��RF-�@��E4@��hӐ!?�-n2G�@>+���ٿ������@��vZ4@��f{�!?�u�1�R�@>+���ٿ������@��vZ4@��f{�!?�u�1�R�@>+���ٿ������@��vZ4@��f{�!?�u�1�R�@��w�|�ٿ��s7�J�@u3}��3@S���_�!?�nV��@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@:҉*�ٿG�֞pU�@FM���3@T��u�!?U����@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@Y���ٿ*>���@�#���4@�:r�a�!?�� �#�@ kr?��ٿx�'��@����94@��z�!?��Α'�@ kr?��ٿx�'��@����94@��z�!?��Α'�@���4�ٿ�rom��@/A]�>4@_=N���!?�d%o�-�@���4�ٿ�rom��@/A]�>4@_=N���!?�d%o�-�@���4�ٿ�rom��@/A]�>4@_=N���!?�d%o�-�@���4�ٿ�rom��@/A]�>4@_=N���!?�d%o�-�@��战�ٿ�f�;v��@�~�'�/4@Wd�]�!?�+���@��战�ٿ�f�;v��@�~�'�/4@Wd�]�!?�+���@��战�ٿ�f�;v��@�~�'�/4@Wd�]�!?�+���@9d+[S�ٿ�^St'��@��# 04@A��Rސ!?�6�߮ҕ@�;����ٿ!�H*��@#��2�t4@'�	���!?L>����@�;����ٿ!�H*��@#��2�t4@'�	���!?L>����@�;����ٿ!�H*��@#��2�t4@'�	���!?L>����@�;����ٿ!�H*��@#��2�t4@'�	���!?L>����@�u���ٿ+�&�Md�@Bo^�14@� ���!?uZ�A�@i�أ�ٿ��/��@�@���4@C���ѐ!?؏I�@i�أ�ٿ��/��@�@���4@C���ѐ!?؏I�@i�أ�ٿ��/��@�@���4@C���ѐ!?؏I�@z��R`�ٿ�=,�*��@݂q�O�3@�D�(�!?w�?�ӕ@��J���ٿ$���y�@��e�4@:�3�!?��{���@o!k�;�ٿ�M���@�Mwl��3@���w�!?����`�@o!k�;�ٿ�M���@�Mwl��3@���w�!?����`�@o!k�;�ٿ�M���@�Mwl��3@���w�!?����`�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@j����ٿM�q�?��@0����3@r.��`�!?��8~T�@���]�ٿ�V����@�9���3@�J��7�!?��E!.F�@V���ٿGh��hE�@B��4@��Ď�!?���huL�@V���ٿGh��hE�@B��4@��Ď�!?���huL�@V���ٿGh��hE�@B��4@��Ď�!?���huL�@V���ٿGh��hE�@B��4@��Ď�!?���huL�@V���ٿGh��hE�@B��4@��Ď�!?���huL�@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@W�/"�ٿ�d3�A�@�ExtC4@'&&ϐ!?���Օ@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@�m'��ٿ�{֙��@�,��U�3@t %��!?�k(Y�@ϩ2�,�ٿA[3U�@�	���3@�X���!?<�G[s�@犠��ٿ�qZ9�Y�@*x��*-4@���Q��!?�7_q��@犠��ٿ�qZ9�Y�@*x��*-4@���Q��!?�7_q��@犠��ٿ�qZ9�Y�@*x��*-4@���Q��!?�7_q��@犠��ٿ�qZ9�Y�@*x��*-4@���Q��!?�7_q��@�+hl��ٿ݄Yp*��@n�R;X4@o��|�!?�\�7��@��;D�ٿ<d�����@��<r�b4@[8�Bo�!?;h�9k�@,�8s�ٿ�e��o��@�:��54@+jG���!?�S���@,�8s�ٿ�e��o��@�:��54@+jG���!?�S���@,�8s�ٿ�e��o��@�:��54@+jG���!?�S���@��τ�ٿ4���3��@h��RkT4@�z��P�!?�W�`��@��τ�ٿ4���3��@h��RkT4@�z��P�!?�W�`��@����;�ٿ�aG $y�@p�x (4@������!?�������@����;�ٿ�aG $y�@p�x (4@������!?�������@�ԇO�ٿ��`^h�@(/;� T4@�p�!?Z��p�@�ԇO�ٿ��`^h�@(/;� T4@�p�!?Z��p�@�ԇO�ٿ��`^h�@(/;� T4@�p�!?Z��p�@��Q$�ٿ�KA���@�*��b4@�x�ڊ�!?��g��T�@��Q$�ٿ�KA���@�*��b4@�x�ڊ�!?��g��T�@��Q$�ٿ�KA���@�*��b4@�x�ڊ�!?��g��T�@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@�RSۥٿ2�Ǳ��@�/�y�4@�ƭ~�!?F��։ו@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@a�i�*�ٿ�9�c�@�K1%$4@@r�'��!?/�﹕@�S{<9�ٿ�'��v��@GV|�(4@���|�!?�ݕy-ʕ@޴3@.�ٿT�]Y�J�@��I�O}4@��z�!?~�'�h��@޴3@.�ٿT�]Y�J�@��I�O}4@��z�!?~�'�h��@޴3@.�ٿT�]Y�J�@��I�O}4@��z�!?~�'�h��@޴3@.�ٿT�]Y�J�@��I�O}4@��z�!?~�'�h��@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@9v���ٿ¯�6��@���X4@����r�!?B�(Ξ�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�#�_�ٿ���k�@���DE4@�M0�!?+u��L�@�]z��ٿݥ�u��@��ѭ�3@��9�!?	��?;�@A�~��ٿJN�=#�@�be�?54@$En��!?ML�=Ε@A�~��ٿJN�=#�@�be�?54@$En��!?ML�=Ε@A�~��ٿJN�=#�@�be�?54@$En��!?ML�=Ε@A�~��ٿJN�=#�@�be�?54@$En��!?ML�=Ε@]���ٿ�`C}��@H�B�
4@l��i�!? 6�~�@�P�n��ٿ���H��@�iP��4@���F�!?f�-)���@�P�n��ٿ���H��@�iP��4@���F�!?f�-)���@,m���ٿ��@�N��@�OYp�)4@�8զU�!?ՆЮ�j�@���@�ٿ�K���@�7�bB04@�I����!?1^�Kؖ@���@�ٿ�K���@�7�bB04@�I����!?1^�Kؖ@���@�ٿ�K���@�7�bB04@�I����!?1^�Kؖ@���ٿ�t���`�@�`��754@���q�!?�Hb�~�@F���g�ٿ,�\��@8�C�4@���9�!?)[�c��@F���g�ٿ,�\��@8�C�4@���9�!?)[�c��@F���g�ٿ,�\��@8�C�4@���9�!?)[�c��@���̖ٿ�)�K��@�ۉ9�A4@z�F~.�!?b�t�`s�@���̖ٿ�)�K��@�ۉ9�A4@z�F~.�!?b�t�`s�@���̖ٿ�)�K��@�ۉ9�A4@z�F~.�!?b�t�`s�@������ٿ�>��z��@�kd\Sc4@�]�b�!?��?�!^�@������ٿ�>��z��@�kd\Sc4@�]�b�!?��?�!^�@������ٿ�>��z��@�kd\Sc4@�]�b�!?��?�!^�@������ٿ�>��z��@�kd\Sc4@�]�b�!?��?�!^�@��q�ٿ����$��@?�4p<?4@�6Ҿ�!?O� ���@��q�ٿ����$��@?�4p<?4@�6Ҿ�!?O� ���@��q�ٿ����$��@?�4p<?4@�6Ҿ�!?O� ���@EÖn9�ٿ)�ЄZ��@��K�4@r+�(�!?,�Rҕ@e��B|�ٿ+�ѝ���@*�W@�3@��gg�!?������@e��B|�ٿ+�ѝ���@*�W@�3@��gg�!?������@e��B|�ٿ+�ѝ���@*�W@�3@��gg�!?������@,!	�ٿ׌��N�@�܈���3@8�<�p�!?O��8��@�J�;�ٿ-{|��@�\��&4@w��  �!?9���F�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@"^@eݝٿ�1iy���@"�:X�D4@գa�&�!?�H�%�B�@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�í^��ٿ�Qx4�g�@�b̫�O4@����O�!?��S�ߕ@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@�;�S�ٿ��'�.�@a�7F4@ADK�+�!?�U/��#�@7L��ٿ�ih��@m�0:4@_�Q�b�!?��8n��@7L��ٿ�ih��@m�0:4@_�Q�b�!?��8n��@7L��ٿ�ih��@m�0:4@_�Q�b�!?��8n��@7L��ٿ�ih��@m�0:4@_�Q�b�!?��8n��@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@8xjn��ٿ��ͼ��@���4@<��!?�m���#�@�Z��E�ٿj!�{��@�>d��64@��]@D�!?fNC�n�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@ky����ٿU�+��@�Þ�4@�8K��!?z:�lxD�@�Y�E��ٿh2A�j#�@=�W�G4@cq�>�!?6�h�(�@�Y�E��ٿh2A�j#�@=�W�G4@cq�>�!?6�h�(�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@���T�ٿ�A��f�@��L44@sNd�P�!?A�s$�;�@�����ٿ�z��L��@)���4@\Zl�!?׈���G�@�����ٿ�z��L��@)���4@\Zl�!?׈���G�@�����ٿ�z��L��@)���4@\Zl�!?׈���G�@�����ٿ�z��L��@)���4@\Zl�!?׈���G�@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@��dQ�ٿL�X�&�@�I#�J4@���9�!?�#w��@�Uz7�ٿ�;G��%�@څ��14@��%�!?�z��}�@�Uz7�ٿ�;G��%�@څ��14@��%�!?�z��}�@�Uz7�ٿ�;G��%�@څ��14@��%�!?�z��}�@�B��ߕٿJ��}�@"r�E54@�
]�!?����dڕ@�2*bg�ٿ(�5����@"�pYvk4@�nh&c�!?z+��}��@�2*bg�ٿ(�5����@"�pYvk4@�nh&c�!?z+��}��@�2*bg�ٿ(�5����@"�pYvk4@�nh&c�!?z+��}��@�2*bg�ٿ(�5����@"�pYvk4@�nh&c�!?z+��}��@�2*bg�ٿ(�5����@"�pYvk4@�nh&c�!?z+��}��@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@P]i?��ٿ�8�����@>z�x1'4@p�@]s�!? �R�A�@<I����ٿ�d'e2�@V=����3@��K&<�!?FV��N�@����ٿP����@\�U�=�3@Z>��L�!?��Iԕ@����ٿP����@\�U�=�3@Z>��L�!?��Iԕ@zfK��ٿ�0�N-�@17;�:�3@q���4�!?�B����@���͘ٿ8΋*z��@�<�\w�3@�R�;�!?+/5��ە@���͘ٿ8΋*z��@�<�\w�3@�R�;�!?+/5��ە@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@��!>�ٿ�.�n��@u�� 4@l���!?��n�ɕ@^a�.��ٿ��� b�@G�s�7�3@�h��F�!?d�����@^a�.��ٿ��� b�@G�s�7�3@�h��F�!?d�����@^a�.��ٿ��� b�@G�s�7�3@�h��F�!?d�����@^a�.��ٿ��� b�@G�s�7�3@�h��F�!?d�����@�����ٿ�q��Z
�@�1�,��3@[��!?f45.^�@ꍁͪ�ٿͤ2��@�9���3@9�4[��!?��Y�7�@ꍁͪ�ٿͤ2��@�9���3@9�4[��!?��Y�7�@ꍁͪ�ٿͤ2��@�9���3@9�4[��!?��Y�7�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@ڃKT��ٿ��W���@�� UY�3@&|��d�!?M^��;�@��3s;�ٿ�3=��W�@`�0L�3@S�y�!?
���O�@H7s��ٿT(�:�m�@��I�,4@��_��!?��2��@��J`�ٿ��|CA��@�C�(4@�1�o�!?�S=A���@��J`�ٿ��|CA��@�C�(4@�1�o�!?�S=A���@��J`�ٿ��|CA��@�C�(4@�1�o�!?�S=A���@�C��6�ٿ&�[R\��@�= )b4@/i���!?$+��<�@�C��6�ٿ&�[R\��@�= )b4@/i���!?$+��<�@G# ��ٿB��k�@$"�m��3@���e�!?�i��*�@G# ��ٿB��k�@$"�m��3@���e�!?�i��*�@G# ��ٿB��k�@$"�m��3@���e�!?�i��*�@G# ��ٿB��k�@$"�m��3@���e�!?�i��*�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@�#���ٿ�����9�@�,�S4@m~��}�!?w�|�+�@��@�ٿ�u�����@:���4@���R�!?e� 3s��@��@�ٿ�u�����@:���4@���R�!?e� 3s��@��@�ٿ�u�����@:���4@���R�!?e� 3s��@��@�ٿ�u�����@:���4@���R�!?e� 3s��@��@�ٿ�u�����@:���4@���R�!?e� 3s��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@�����ٿf��!���@=�[U�4@��ef�!?�d��@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@������ٿ��d��Z�@�(
<1�3@�	���!?
��~���@�8���ٿ_�����@O�2�4	4@�P��!?S}�r�Q�@�8���ٿ_�����@O�2�4	4@�P��!?S}�r�Q�@�2&D�ٿ�ذL.��@^�4@���2�!?*��)�@����̢ٿ8M����@�z���3@��x�l�!?�vXNr�@����̢ٿ8M����@�z���3@��x�l�!?�vXNr�@����̢ٿ8M����@�z���3@��x�l�!?�vXNr�@����̢ٿ8M����@�z���3@��x�l�!?�vXNr�@����̢ٿ8M����@�z���3@��x�l�!?�vXNr�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@�=|��ٿd2�U��@�����3@��p@�!?QT�n[�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@O��~��ٿ�־Tr�@�$n�G	4@f�2w�!?�~#d�D�@%��ٿn��s�@+�{ĝ'4@Z~�k�!?�#�ygÕ@%��ٿn��s�@+�{ĝ'4@Z~�k�!?�#�ygÕ@%��ٿn��s�@+�{ĝ'4@Z~�k�!?�#�ygÕ@%��ٿn��s�@+�{ĝ'4@Z~�k�!?�#�ygÕ@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@�7�x�ٿ~�L���@�ӥN4@��[@�!?,�,��@��7��ٿ�.:���@^���+4@$(�#�!?-/�W� �@��5ۜٿ���R�@�P���'4@]��>�!?)�å;��@��5ۜٿ���R�@�P���'4@]��>�!?)�å;��@E�LJ�ٿ|�M@��@T"s�'4@d�,on�!?(�? ��@E�LJ�ٿ|�M@��@T"s�'4@d�,on�!?(�? ��@E�LJ�ٿ|�M@��@T"s�'4@d�,on�!?(�? ��@E�LJ�ٿ|�M@��@T"s�'4@d�,on�!?(�? ��@����ٿ"� ��@�rM"�B4@���s]�!?٬��+ʕ@����ٿ"� ��@�rM"�B4@���s]�!?٬��+ʕ@����ٿ"� ��@�rM"�B4@���s]�!?٬��+ʕ@����ٿ"� ��@�rM"�B4@���s]�!?٬��+ʕ@����ٿ"� ��@�rM"�B4@���s]�!?٬��+ʕ@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@����ٿ_�V;ݿ�@����HE4@Ǭ����!?�S��f�@ݰ�p	�ٿ�O����@�_J��3@mMn�!?�pK����@ݰ�p	�ٿ�O����@�_J��3@mMn�!?�pK����@ݰ�p	�ٿ�O����@�_J��3@mMn�!?�pK����@ݰ�p	�ٿ�O����@�_J��3@mMn�!?�pK����@��,�ٿBگ�i��@���?4@�!
㡐!?!���9�@������ٿ��k���@� �]�4@�[t�Ȑ!?.ˤN��@������ٿ��k���@� �]�4@�[t�Ȑ!?.ˤN��@������ٿ��k���@� �]�4@�[t�Ȑ!?.ˤN��@������ٿ��k���@� �]�4@�[t�Ȑ!?.ˤN��@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@w��O�ٿ�"|k/�@�Z4��3@����v�!?�������@1۶�ěٿS�&��W�@]�� K4@{��p�!?�&/�ȕ@B�G�s�ٿt�J5�V�@���&�34@e��x�!?,�rS���@B�G�s�ٿt�J5�V�@���&�34@e��x�!?,�rS���@B�G�s�ٿt�J5�V�@���&�34@e��x�!?,�rS���@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@��|ٞٿ�4K8�@�� 74@qQ0���!?qT�R��@�8{�ٿ�(Ԋ��@��F�� 4@E�bថ!?L_:�s1�@�8{�ٿ�(Ԋ��@��F�� 4@E�bថ!?L_:�s1�@�8{�ٿ�(Ԋ��@��F�� 4@E�bថ!?L_:�s1�@rG�\��ٿ��zH
�@��\�A4@H��9�!?��.ݕ@rG�\��ٿ��zH
�@��\�A4@H��9�!?��.ݕ@ylu�ٿ��o���@O����+4@R.Z��!?�9?;0��@ylu�ٿ��o���@O����+4@R.Z��!?�9?;0��@ylu�ٿ��o���@O����+4@R.Z��!?�9?;0��@ylu�ٿ��o���@O����+4@R.Z��!?�9?;0��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@;�޻ �ٿ�I�3a��@祺+�4@8�qs�!?:�7��@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�;���ٿ��� ���@0��+L4@��rVd�!?�!�]X˕@�7��ٿ,R�8r�@��O�%4@�-���!?�����@�7��ٿ,R�8r�@��O�%4@�-���!?�����@�7��ٿ,R�8r�@��O�%4@�-���!?�����@�7��ٿ,R�8r�@��O�%4@�-���!?�����@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@t�X��ٿ��I>�@�}xO<4@�C�O�!?�kE��@�vT1��ٿ���Na�@Q�LY4@FAN�R�!?: K�ӕ@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@����ٿ�.�h��@Qc���4@:��X3�!?���w�@�}t��ٿܠ�".�@�32���3@��p�'�!?���Z�?�@�}t��ٿܠ�".�@�32���3@��p�'�!?���Z�?�@�& /*�ٿ�2q���@I�4�4@�!��!?����u-�@�w��̚ٿ�ۤ��@���_P4@����9�!?i�m��ϕ@�w��̚ٿ�ۤ��@���_P4@����9�!?i�m��ϕ@�w��̚ٿ�ۤ��@���_P4@����9�!?i�m��ϕ@�w��̚ٿ�ۤ��@���_P4@����9�!?i�m��ϕ@ϒ�^@�ٿP�#g ��@k2�.4@���G[�!?�� ��F�@ϒ�^@�ٿP�#g ��@k2�.4@���G[�!?�� ��F�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@<(bn�ٿ�=� +a�@*�e�>4@%��u]�!?|P�f�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@�����ٿ���d���@2��4@p�t�K�!?TWK.?�@C�QJ�ٿ$wϣ��@K~�,14@�n��P�!?B":�@���M�ٿ��`�w�@L|��+4@j�0?�!?�2
/@�@���M�ٿ��`�w�@L|��+4@j�0?�!?�2
/@�@�ٝٿ���<���@� :�z�3@�NqDR�!?)��1]W�@�G/�ٿ�D}�v;�@�G�J#(4@KVL�w�!?\��X`
�@�G/�ٿ�D}�v;�@�G�J#(4@KVL�w�!?\��X`
�@�Ĵ��ٿ�Z����@�-ݫ�4@�mݺM�!?����@�Ĵ��ٿ�Z����@�-ݫ�4@�mݺM�!?����@�Ĵ��ٿ�Z����@�-ݫ�4@�mݺM�!?����@�Ĵ��ٿ�Z����@�-ݫ�4@�mݺM�!?����@�Ĵ��ٿ�Z����@�-ݫ�4@�mݺM�!?����@�xI�>�ٿ'���w�@o��J�4@"�z�^�!??�lc^�@�xI�>�ٿ'���w�@o��J�4@"�z�^�!??�lc^�@y�/bJ�ٿ���h�@UH]�Z4@sIbE�!? ����H�@y�/bJ�ٿ���h�@UH]�Z4@sIbE�!? ����H�@�p�s?�ٿ?y�Z< �@���{%4@J�_��!?o�	��2�@�p�s?�ٿ?y�Z< �@���{%4@J�_��!?o�	��2�@�p�s?�ٿ?y�Z< �@���{%4@J�_��!?o�	��2�@�p�s?�ٿ?y�Z< �@���{%4@J�_��!?o�	��2�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�˸D�ٿ�x�0�@�S4@��B �!?�1b�@�Z��ٿ���Cx�@� ��4@7��!?����m�@�Z��ٿ���Cx�@� ��4@7��!?����m�@�u�E�ٿ �� ��@���	4@):�"�!?[S&Yb�@�u�E�ٿ �� ��@���	4@):�"�!?[S&Yb�@�u�E�ٿ �� ��@���	4@):�"�!?[S&Yb�@�u�E�ٿ �� ��@���	4@):�"�!?[S&Yb�@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@���Z�ٿ�Q�:E��@6<�Q�3@,�!?:���@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@m��㨣ٿ�����K�@��q�3@Jx�!?t�)��@%��>�ٿe�����@����3@����!�!?�o���#�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@��$V�ٿ�ۏ}r:�@�3H��4@f��!�!?Rg�#h�@i�0I�ٿ�e<| �@��S�)4@B�v\�!?%�ټ�U�@i�0I�ٿ�e<| �@��S�)4@B�v\�!?%�ټ�U�@i�0I�ٿ�e<| �@��S�)4@B�v\�!?%�ټ�U�@	����ٿ�}�*�@�Ɓ۫K4@/��G�!?�>���i�@	����ٿ�}�*�@�Ɓ۫K4@/��G�!?�>���i�@	����ٿ�}�*�@�Ɓ۫K4@/��G�!?�>���i�@	����ٿ�}�*�@�Ɓ۫K4@/��G�!?�>���i�@	����ٿ�}�*�@�Ɓ۫K4@/��G�!?�>���i�@���R�ٿs,,���@LY��M4@���{�!?�w(y�@���R�ٿs,,���@LY��M4@���{�!?�w(y�@���R�ٿs,,���@LY��M4@���{�!?�w(y�@������ٿ|c���@;,M<'4@f���!?Ű�g���@��rIV�ٿ�k��r��@�[&�4@��fji�!?�cS�EC�@��rIV�ٿ�k��r��@�[&�4@��fji�!?�cS�EC�@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@Ћ��؛ٿ��ڨ���@W�� m�3@��AON�!?��o��ϕ@��_���ٿ�1.6w��@��#�!4@򌐍\�!?׬jN��@��_���ٿ�1.6w��@��#�!4@򌐍\�!?׬jN��@�c�y�ٿ����{��@�שx��3@��]sW�!?NL�wLv�@�c�y�ٿ����{��@�שx��3@��]sW�!?NL�wLv�@@I�w�ٿ�C��_�@��c3s�3@&�H�!?�2�u��@@I�w�ٿ�C��_�@��c3s�3@&�H�!?�2�u��@@I�w�ٿ�C��_�@��c3s�3@&�H�!?�2�u��@�aȖ
�ٿ���S��@c��P4@��bX
�!?G*�m�p�@�aȖ
�ٿ���S��@c��P4@��bX
�!?G*�m�p�@�aȖ
�ٿ���S��@c��P4@��bX
�!?G*�m�p�@�aȖ
�ٿ���S��@c��P4@��bX
�!?G*�m�p�@�aȖ
�ٿ���S��@c��P4@��bX
�!?G*�m�p�@J���ٿ^�t>̍�@d���f4@}���!?ڍY�.̕@RM���ٿ|�sm �@�|k_4@t�ʌ��!?����B�@RM���ٿ|�sm �@�|k_4@t�ʌ��!?����B�@RM���ٿ|�sm �@�|k_4@t�ʌ��!?����B�@RM���ٿ|�sm �@�|k_4@t�ʌ��!?����B�@h�{��ٿ@P�s4�@��	�B4@�\P�!?B�a�҅�@h�{��ٿ@P�s4�@��	�B4@�\P�!?B�a�҅�@h�{��ٿ@P�s4�@��	�B4@�\P�!?B�a�҅�@h�{��ٿ@P�s4�@��	�B4@�\P�!?B�a�҅�@�3���ٿ� �� �@4=,�`4@��X<!�!?��/�ܑ�@@of�ڠٿ���^��@��T�3@X��u�!?!�2H�ƕ@@of�ڠٿ���^��@��T�3@X��u�!?!�2H�ƕ@R/ܢٿ�c�@��@C����4@���Y��!?$Hm���@R/ܢٿ�c�@��@C����4@���Y��!?$Hm���@�/K9�ٿ��>�R�@	!�� 4@Z�;��!?��<�v�@�/K9�ٿ��>�R�@	!�� 4@Z�;��!?��<�v�@��*ܜٿQ"����@/��'14@a����!?����@�@��*ܜٿQ"����@/��'14@a����!?����@�@��*ܜٿQ"����@/��'14@a����!?����@�@c�s��ٿۨ��9�@�r�<4@�h��!?p���eڕ@c�s��ٿۨ��9�@�r�<4@�h��!?p���eڕ@|{�y�ٿR��O���@��cs4@�s�~�!?i�?��2�@|{�y�ٿR��O���@��cs4@�s�~�!?i�?��2�@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@e�����ٿX.���@�$���3@�I^G�!?�"�ZZ��@p�����ٿ�"�A���@�����4@��E� �!?���Up�@Mz���ٿ��^��@��d.4@�x���!?&��=��@Mz���ٿ��^��@��d.4@�x���!?&��=��@7_M�0�ٿ�C�@!��[J4@��Z�?�!?�K�d�E�@7_M�0�ٿ�C�@!��[J4@��Z�?�!?�K�d�E�@7_M�0�ٿ�C�@!��[J4@��Z�?�!?�K�d�E�@7_M�0�ٿ�C�@!��[J4@��Z�?�!?�K�d�E�@��z�ٿc�U�_�@ħ��74@j�^�N�!?���U\�@��z�ٿc�U�_�@ħ��74@j�^�N�!?���U\�@H�<Нٿ3�p^Q�@/���3@��A��!?�zR2�B�@H�<Нٿ3�p^Q�@/���3@��A��!?�zR2�B�@H�<Нٿ3�p^Q�@/���3@��A��!?�zR2�B�@H�<Нٿ3�p^Q�@/���3@��A��!?�zR2�B�@�1���ٿI8U��@ ~I���3@�~�嫐!?{�͙�@�1���ٿI8U��@ ~I���3@�~�嫐!?{�͙�@�1���ٿI8U��@ ~I���3@�~�嫐!?{�͙�@�1���ٿI8U��@ ~I���3@�~�嫐!?{�͙�@�1���ٿI8U��@ ~I���3@�~�嫐!?{�͙�@�ZP�h�ٿy4Сr��@ƭ�>�3@�/�v�!?��|�^�@�ZP�h�ٿy4Сr��@ƭ�>�3@�/�v�!?��|�^�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@���W՘ٿ+�''���@�(�X4@�d�G��!?Ѭ�~�@i�S:g�ٿ�m��$��@���I�4@�@&P�!?`[�ҹ�@i�S:g�ٿ�m��$��@���I�4@�@&P�!?`[�ҹ�@i�S:g�ٿ�m��$��@���I�4@�@&P�!?`[�ҹ�@i�S:g�ٿ�m��$��@���I�4@�@&P�!?`[�ҹ�@D��|Ӝٿ�%����@��~&4@^�����!?Q�u?a�@D��|Ӝٿ�%����@��~&4@^�����!?Q�u?a�@D��|Ӝٿ�%����@��~&4@^�����!?Q�u?a�@�Ɣ:��ٿ�d����@-�v��_4@�>�n�!?
����k�@�Ɣ:��ٿ�d����@-�v��_4@�>�n�!?
����k�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@�R���ٿ�`B$�+�@X��ڞW4@� �О�!?q��BN�@خ�a�ٿ��0���@K�̥'4@��{2�!?��j���@خ�a�ٿ��0���@K�̥'4@��{2�!?��j���@خ�a�ٿ��0���@K�̥'4@��{2�!?��j���@خ�a�ٿ��0���@K�̥'4@��{2�!?��j���@ υ�2�ٿ8��X�@�v�,Y94@����,�!?��j�@2�E�ՠٿo~���@�+�F4@~�n�^�!?�j��@2�E�ՠٿo~���@�+�F4@~�n�^�!?�j��@2�E�ՠٿo~���@�+�F4@~�n�^�!?�j��@���Z��ٿ�^��{(�@��]�:4@5�)L�!?{8OO��@���Z��ٿ�^��{(�@��]�:4@5�)L�!?{8OO��@���Z��ٿ�^��{(�@��]�:4@5�)L�!?{8OO��@���Z��ٿ�^��{(�@��]�:4@5�)L�!?{8OO��@�#M4��ٿ�?�:<�@���4@���j�!?�r� �i�@�#M4��ٿ�?�:<�@���4@���j�!?�r� �i�@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@#���u�ٿs��1���@��dU��3@h�).R�!?ȹ'wh��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@U׿��ٿL���ɝ�@̍S�4@�{�!?�aɓ��@j��|�ٿ�Ay��-�@�����4@*�$�ݏ!?i��p'�@j��|�ٿ�Ay��-�@�����4@*�$�ݏ!?i��p'�@c�ݏ�ٿ���AG
�@<��.��3@���J�!?��m�@c�ݏ�ٿ���AG
�@<��.��3@���J�!?��m�@c�ݏ�ٿ���AG
�@<��.��3@���J�!?��m�@c�ݏ�ٿ���AG
�@<��.��3@���J�!?��m�@�����ٿ���%T�@�ن7��3@��{]�!?���?���@�����ٿ���%T�@�ن7��3@��{]�!?���?���@�����ٿ���%T�@�ن7��3@��{]�!?���?���@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@���^�ٿ��M�o�@W{���3@�ٚ�%�!?d8~y�@[�D�ݟٿf����"�@n��/��3@�4��!?#X�4�c�@[�D�ݟٿf����"�@n��/��3@�4��!?#X�4�c�@[�D�ݟٿf����"�@n��/��3@�4��!?#X�4�c�@՟��ٿCҍ��@�}a�Z4@9�"%�!?�1���8�@�s�2ՙٿ ���%�@ߛ��54@Κ_��!?�$@R�@�s�2ՙٿ ���%�@ߛ��54@Κ_��!?�$@R�@�AHq?�ٿT�w����@ը9I 4@���C�!?e��a��@�AHq?�ٿT�w����@ը9I 4@���C�!?e��a��@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@��#Б�ٿ���\��@��l4@�+�I&�!?M'6Z(�@�Z<ᶡٿKOk�O:�@��ƛc\4@��P��!?��L���@�Z<ᶡٿKOk�O:�@��ƛc\4@��P��!?��L���@,�産�ٿ}R�����@�d
gr94@
���!?l�B���@,�産�ٿ}R�����@�d
gr94@
���!?l�B���@,�産�ٿ}R�����@�d
gr94@
���!?l�B���@,�産�ٿ}R�����@�d
gr94@
���!?l�B���@{��B�ٿ���M�@b`YK�/4@��J �!?��E\4E�@{��B�ٿ���M�@b`YK�/4@��J �!?��E\4E�@{��B�ٿ���M�@b`YK�/4@��J �!?��E\4E�@{��B�ٿ���M�@b`YK�/4@��J �!?��E\4E�@]C����ٿ���e���@�4S��14@�8-�!�!?'�Ð��@]C����ٿ���e���@�4S��14@�8-�!�!?'�Ð��@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@+<�ٿR��o>8�@d@��4@&GN�@�!?H>�M=�@��ų�ٿib��@�+�Ʀ�3@��8�!?�#��C��@��ų�ٿib��@�+�Ʀ�3@��8�!?�#��C��@Qi��j�ٿ��	��@��A��3@Zd}�g�!?vU�ocѕ@̏A���ٿM�Ұ:�@������3@ɶ�7>�!?�y��ã�@̏A���ٿM�Ұ:�@������3@ɶ�7>�!?�y��ã�@̏A���ٿM�Ұ:�@������3@ɶ�7>�!?�y��ã�@̏A���ٿM�Ұ:�@������3@ɶ�7>�!?�y��ã�@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@ǒs|��ٿʷJ�P��@�7yr4@�VگE�!?�������@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@<iݑ�ٿ�6Lɫ�@�k��4@}���w�!?�Ќ�F�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@��m��ٿ� ��ާ�@����4@ՁX��!?zI&S0�@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@n�Dn��ٿ#��7��@kd:���3@Cē\�!?e$����@�Ta�s�ٿĳ/B�g�@Fz��3@Q��q�!?:P[�@�Ta�s�ٿĳ/B�g�@Fz��3@Q��q�!?:P[�@��k㳘ٿ��b��@~��u+D4@��QO�!?ݰ���@C�|�,�ٿ'"!�	�@�e�n4@�s'�P�!?!
�o��@C�|�,�ٿ'"!�	�@�e�n4@�s'�P�!?!
�o��@C�|�,�ٿ'"!�	�@�e�n4@�s'�P�!?!
�o��@C�|�,�ٿ'"!�	�@�e�n4@�s'�P�!?!
�o��@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@/�>.�ٿ�r~mX��@��Du�m4@�o�[�!?����⹕@aL�2C�ٿe7׆4�@:F�P44@�|!w�!?w�(��*�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@JH��]�ٿU;Ƨ\��@a��,�3@G��C�!?
�"�@��BJ؟ٿd_!|s��@�Q�&4@���lo�!?��;i�'�@GeD((�ٿ�$���@�ņq�(4@�)�]�!? ,b0ו@GeD((�ٿ�$���@�ņq�(4@�)�]�!? ,b0ו@GeD((�ٿ�$���@�ņq�(4@�)�]�!? ,b0ו@GeD((�ٿ�$���@�ņq�(4@�)�]�!? ,b0ו@GeD((�ٿ�$���@�ņq�(4@�)�]�!? ,b0ו@DWǉ�ٿ�G݂��@�q���94@���EY�!?�)|�婕@DWǉ�ٿ�G݂��@�q���94@���EY�!?�)|�婕@��\��ٿ9���B��@�.��44@#_o*�!?�lK��@��\��ٿ9���B��@�.��44@#_o*�!?�lK��@��\��ٿ9���B��@�.��44@#_o*�!?�lK��@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@M��b�ٿ&���&��@
�*�"4@�G���!?K*����@y�b9|�ٿh�%���@1���4@���E�!?�����e�@y�b9|�ٿh�%���@1���4@���E�!?�����e�@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@m곽 �ٿV����@��Em4@��hyY�!?pYM2ߕ@y�h�ןٿ��ҶF�@����;	4@�����!?�OI�u$�@y�h�ןٿ��ҶF�@����;	4@�����!?�OI�u$�@���Z�ٿ[��+�@Zf���3@�Q8C�!?��X���@���Z�ٿ[��+�@Zf���3@�Q8C�!?��X���@p����ٿR�zⴹ�@6�"$*�3@f��x�!?��5�F�@$�wU�ٿ?:����@�i��R�3@�g�b�!?�|f��a�@$�wU�ٿ?:����@�i��R�3@�g�b�!?�|f��a�@$�wU�ٿ?:����@�i��R�3@�g�b�!?�|f��a�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@^'�?��ٿ���8�}�@ǰX84@_v�#�!?��o�D�@�zqĻ�ٿwE�CS�@���ȝ4@��Tw�!?�\��}�@�zqĻ�ٿwE�CS�@���ȝ4@��Tw�!?�\��}�@�zqĻ�ٿwE�CS�@���ȝ4@��Tw�!?�\��}�@�zqĻ�ٿwE�CS�@���ȝ4@��Tw�!?�\��}�@/x�p�ٿ҆=-�@�$n�3@xrB�!?#�ݹq�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@����ٿ\�؋�P�@���4@ P��!?d���&�@��<�Ρٿ���7�@�7?�3@�V�Q�!?}��1�@��<�Ρٿ���7�@�7?�3@�V�Q�!?}��1�@��<�Ρٿ���7�@�7?�3@�V�Q�!?}��1�@��<�Ρٿ���7�@�7?�3@�V�Q�!?}��1�@��<�Ρٿ���7�@�7?�3@�V�Q�!?}��1�@t0�zn�ٿ���@P����3@}��~�!?�l҆�G�@���J�ٿ��w�͒�@�'8{@�3@*F���!?�R��@���J�ٿ��w�͒�@�'8{@�3@*F���!?�R��@���J�ٿ��w�͒�@�'8{@�3@*F���!?�R��@���J�ٿ��w�͒�@�'8{@�3@*F���!?�R��@���J�ٿ��w�͒�@�'8{@�3@*F���!?�R��@����ٿLZ��nt�@��=�4@tpF��!?�)���,�@����ٿLZ��nt�@��=�4@tpF��!?�)���,�@�t9o7�ٿo��93�@��[�J04@��o��!?���D}�@�t9o7�ٿo��93�@��[�J04@��o��!?���D}�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@
d�cV�ٿ�ú7���@7�:3M4@֔eGِ!?G�X袙�@�r�9]�ٿ�<�*ؾ�@o��w��3@�A���!?��eB�q�@�r�9]�ٿ�<�*ؾ�@o��w��3@�A���!?��eB�q�@��VZ�ٿ�GS�7�@P�V4@�$D!�!?����dN�@��VZ�ٿ�GS�7�@P�V4@�$D!�!?����dN�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@�$eC�ٿL^qp]��@�A�V/4@JdWj��!?����0O�@~���ٿWT+N=S�@�a�D�"4@�"8�!?+�ŕ��@~���ٿWT+N=S�@�a�D�"4@�"8�!?+�ŕ��@~���ٿWT+N=S�@�a�D�"4@�"8�!?+�ŕ��@~���ٿWT+N=S�@�a�D�"4@�"8�!?+�ŕ��@~���ٿWT+N=S�@�a�D�"4@�"8�!?+�ŕ��@l`ʊ�ٿi>R���@����04@�ϵF��!?������@U��C+�ٿ�o0�l��@$\EH*94@#�췅�!?�8Θ�,�@�:a���ٿ�^�8}��@�M�}�84@�S�(�!?n����@�:a���ٿ�^�8}��@�M�}�84@�S�(�!?n����@�:a���ٿ�^�8}��@�M�}�84@�S�(�!?n����@�����ٿ��п��@��c�{\4@�*^��!?H�Rҕ@�����ٿ��п��@��c�{\4@�*^��!?H�Rҕ@�����ٿ��п��@��c�{\4@�*^��!?H�Rҕ@�����ٿ��п��@��c�{\4@�*^��!?H�Rҕ@�����ٿ��п��@��c�{\4@�*^��!?H�Rҕ@qr�C�ٿg������@	�|�.t4@t``q�!?�?ƴ��@qr�C�ٿg������@	�|�.t4@t``q�!?�?ƴ��@qr�C�ٿg������@	�|�.t4@t``q�!?�?ƴ��@qr�C�ٿg������@	�|�.t4@t``q�!?�?ƴ��@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@u�7��ٿ�Z}.�S�@euF��34@C�2��!?֔����@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@0���ٿ��ú���@�����4@���5m�!?6!m㓰�@9���ٛٿ����+�@���4@{fF��!?m�aǉ`�@9���ٛٿ����+�@���4@{fF��!?m�aǉ`�@9���ٛٿ����+�@���4@{fF��!?m�aǉ`�@���Yٞٿ��?�]�@2Y:4@~qN�!?�*�kC�@���Yٞٿ��?�]�@2Y:4@~qN�!?�*�kC�@3{�ϕٿ��L���@̥���04@F�Ӭ��!?�~+����@3{�ϕٿ��L���@̥���04@F�Ӭ��!?�~+����@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@������ٿE{�֝��@���$4@�P��g�!?Ӳ��P�@(FcK�ٿG��g�@���4@\��!�!?п�kGW�@��ٿ�%GM���@Ǽ1O4@�Q�q�!?IW!�|��@I�0u �ٿ��<����@��[�5"4@�T�K��!?�D���@I�0u �ٿ��<����@��[�5"4@�T�K��!?�D���@���{�ٿ�6 ��@�d��#4@��!Ї�!?�ɕ@���{�ٿ�6 ��@�d��#4@��!Ї�!?�ɕ@���{�ٿ�6 ��@�d��#4@��!Ї�!?�ɕ@���{�ٿ�6 ��@�d��#4@��!Ї�!?�ɕ@���{�ٿ�6 ��@�d��#4@��!Ї�!?�ɕ@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�[񧾙ٿk��i���@��-�.4@ޢ�2�!?��KN��@�"�h�ٿ��
��=�@8 <��<4@Yl�D�!?�WÍ�@�"�h�ٿ��
��=�@8 <��<4@Yl�D�!?�WÍ�@�"�h�ٿ��
��=�@8 <��<4@Yl�D�!?�WÍ�@�"�h�ٿ��
��=�@8 <��<4@Yl�D�!?�WÍ�@u��ћٿ̀��e�@Jw���84@鑆�!?�
����@u��ћٿ̀��e�@Jw���84@鑆�!?�
����@u��ћٿ̀��e�@Jw���84@鑆�!?�
����@u��ћٿ̀��e�@Jw���84@鑆�!?�
����@u��ћٿ̀��e�@Jw���84@鑆�!?�
����@��n�ٿ�B~)���@Q0z���3@��$!?ك��#��@ז�Wϝٿ��M��6�@K��w��3@�"M�!?���^I�@ז�Wϝٿ��M��6�@K��w��3@�"M�!?���^I�@��Pٛٿ��J��@O��Z�3@��T�5�!?gS�7:�@��Pٛٿ��J��@O��Z�3@��T�5�!?gS�7:�@��Pٛٿ��J��@O��Z�3@��T�5�!?gS�7:�@��Pٛٿ��J��@O��Z�3@��T�5�!?gS�7:�@�0�Hٜٿk^����@:�HJ�3@��1�^�!?���z���@�0�Hٜٿk^����@:�HJ�3@��1�^�!?���z���@3	e���ٿ�\(F��@�0�Ŕ4@�@��!?�c�x�@����ٿ�eHq|5�@�����3@�}��!?/ٕ@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@B�u� �ٿd����@9IZ���3@�L:�2�!?b^�S�@�S��ٿ���ma��@@��~�4@��'LY�!?!)A�n+�@�P�48�ٿH�#�M�@�P�4� 4@ �<j�!?���᠕@�'�!�ٿ������@�@��=4@�&߶�!?��--���@�t/4��ٿ�tT{5C�@�͘%p`4@d}�ď!?�9�K�@�t/4��ٿ�tT{5C�@�͘%p`4@d}�ď!?�9�K�@�t/4��ٿ�tT{5C�@�͘%p`4@d}�ď!?�9�K�@�Cӆ��ٿ�������@��`�~p4@�m���!?��>��?�@�Cӆ��ٿ�������@��`�~p4@�m���!?��>��?�@�Cӆ��ٿ�������@��`�~p4@�m���!?��>��?�@����ٿ񣑡���@VaE|�4@�� �!?csf�T�@����ٿ񣑡���@VaE|�4@�� �!?csf�T�@n1�
�ٿ/��ȯ��@�'�ܒ4@%��8�!?\�3�y�@�"�u!�ٿޓ[�j��@Z*o� �3@��I5"�!?k�܇�ڕ@�"�u!�ٿޓ[�j��@Z*o� �3@��I5"�!?k�܇�ڕ@Xϵv��ٿ ����@<J%]��3@�y$Bs�!?-xZj�@+.�ڕ�ٿg$����@YB�c�	4@_��P�!?Vm��,�@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@0w�ET�ٿg1L���@=*ʏ�C4@�8=ze�!?]̩�5͕@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@/Z�!�ٿ�eN--�@��ȃ�4@�����!?�le!V8�@pFI�ٿs?捐�@��H4@� d���!?ђ��4�@eCES>�ٿVd]�!��@��M��4@�]���!?�̀�E�@:��[�ٿ��Kϸ��@5JW���3@9z���!?<Tn�(/�@:��[�ٿ��Kϸ��@5JW���3@9z���!?<Tn�(/�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@�[7+�ٿ�{�&M`�@^]t!j$4@� S�Z�!?DEr&ī�@6�9Bp�ٿ_�]N���@�07Z�3@h��!?���n�@6�9Bp�ٿ_�]N���@�07Z�3@h��!?���n�@6�9Bp�ٿ_�]N���@�07Z�3@h��!?���n�@6�9Bp�ٿ_�]N���@�07Z�3@h��!?���n�@6�9Bp�ٿ_�]N���@�07Z�3@h��!?���n�@�C�ϛٿ\�bSe�@p룾%4@���2�!?R�V��@�?}��ٿ�G�W��@U;�;�:4@Ȟ�O\�!?�B:ͥؕ@�?}��ٿ�G�W��@U;�;�:4@Ȟ�O\�!?�B:ͥؕ@u��d�ٿK�����@+�J�n74@Rx�㬐!?�E��ӽ�@u��d�ٿK�����@+�J�n74@Rx�㬐!?�E��ӽ�@u��d�ٿK�����@+�J�n74@Rx�㬐!?�E��ӽ�@u��d�ٿK�����@+�J�n74@Rx�㬐!?�E��ӽ�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@�^�|�ٿi�nd$�@C�4	:74@1Җun�!?܀��l,�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@	����ٿ��:͉��@m�	�@"4@4�3q�!?���Bk�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�� ��ٿz��?�C�@Ba��:4@!�hE]�!?��g�[Y�@�@88�ٿdlS�U/�@�oBFW64@�[����!?$�	��@�@88�ٿdlS�U/�@�oBFW64@�[����!?$�	��@d�3�)�ٿ#f��@�c=��J4@��x}�!?�-Z^��@d�3�)�ٿ#f��@�c=��J4@��x}�!?�-Z^��@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@���P�ٿ� ����@�,�|�4@�|�ԙ�!??���@f1�WP�ٿ����4/�@P�,��4@���n,�!?SP2�'�@f1�WP�ٿ����4/�@P�,��4@���n,�!?SP2�'�@΃{y��ٿ�,��@��B}K+4@�^3��!?8��Kѕ@΃{y��ٿ�,��@��B}K+4@�^3��!?8��Kѕ@΃{y��ٿ�,��@��B}K+4@�^3��!?8��Kѕ@΃{y��ٿ�,��@��B}K+4@�^3��!?8��Kѕ@B;��"�ٿ�c�[R�@~y�f4@+�J9�!?U����Õ@B;��"�ٿ�c�[R�@~y�f4@+�J9�!?U����Õ@�U�3�ٿ0WAYc�@�L�o`64@�L�s�!?����@�U�3�ٿ0WAYc�@�L�o`64@�L�s�!?����@@ �]�ٿ�2ڗ���@v�t�94@Z	X��!?��^8��@���U�ٿ"�r� ��@fl��44@�{[zz�!?B_��B�@���U�ٿ"�r� ��@fl��44@�{[zz�!?B_��B�@���U�ٿ"�r� ��@fl��44@�{[zz�!?B_��B�@�J�:��ٿ=��4��@����G4@:����!?��m��@�J�:��ٿ=��4��@����G4@:����!?��m��@�J�:��ٿ=��4��@����G4@:����!?��m��@�J�:��ٿ=��4��@����G4@:����!?��m��@�J�:��ٿ=��4��@����G4@:����!?��m��@�L�z)�ٿWR
1���@��Ԍ;:4@P�X��!?d��+�@�L�z)�ٿWR
1���@��Ԍ;:4@P�X��!?d��+�@�L�z)�ٿWR
1���@��Ԍ;:4@P�X��!?d��+�@&t༙ٿ��&+o�@����7G4@_J���!?���
'ӕ@&t༙ٿ��&+o�@����7G4@_J���!?���
'ӕ@C�:�ٿ��dL��@^��ѶT4@I3�!?c�5��@C�:�ٿ��dL��@^��ѶT4@I3�!?c�5��@C�:�ٿ��dL��@^��ѶT4@I3�!?c�5��@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@ �	�ܘٿVr�����@��B�Ub4@L��e�!?K>	E�ȕ@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@j��z��ٿ�������@39�ׁZ4@>.S�I�!?�r�ې@���r�ٿ��Gf]�@,΢� o4@�Bh���!?���@�@��;=��ٿnc���@^�c��Z4@o�(jv�!?l!ʨ]��@��;=��ٿnc���@^�c��Z4@o�(jv�!?l!ʨ]��@��;=��ٿnc���@^�c��Z4@o�(jv�!?l!ʨ]��@��;=��ٿnc���@^�c��Z4@o�(jv�!?l!ʨ]��@3�=Kf�ٿ]NT!��@�3�24@z�y�6�!? mv�ܦ�@��foןٿ��Y�C�@萂�4@p�[N �!?!�h
ӕ@倫o@�ٿ
�s^a�@�|�hF4@�U=�S�!?� M60�@倫o@�ٿ
�s^a�@�|�hF4@�U=�S�!?� M60�@倫o@�ٿ
�s^a�@�|�hF4@�U=�S�!?� M60�@倫o@�ٿ
�s^a�@�|�hF4@�U=�S�!?� M60�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@&��/�ٿ^����@*��0�m4@�Yӄ�!?g �;�i�@;X���ٿ:�n֭��@Rj�D?4@�LǤ��!?Uage��@�=��I�ٿ�U�A�@�_D#+X4@Е;���!?�B1ݕ@�=��I�ٿ�U�A�@�_D#+X4@Е;���!?�B1ݕ@��uy�ٿ�R�v�p�@}��N�f4@������!? �l�b�@��uy�ٿ�R�v�p�@}��N�f4@������!? �l�b�@��uy�ٿ�R�v�p�@}��N�f4@������!? �l�b�@��uy�ٿ�R�v�p�@}��N�f4@������!? �l�b�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@z�bC��ٿ{�@AZ�@{E�I�G4@��<.D�!?�D�I�@lB3E�ٿι[�]b�@��+�4@�r���!?<� 2���@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@Q2�ٿ8��Ч��@ꃺ�3@�lQ�C�!?�O���p�@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@�q_˱�ٿ��?-�O�@ -�4@�2Bv��!?T�R�Օ@w�����ٿ�����@��S^��3@�͚ɰ�!?� �n̕@w�����ٿ�����@��S^��3@�͚ɰ�!?� �n̕@�1c�ٿ%B�k��@�Z�L4@�Ȱ���!?���"��@�1c�ٿ%B�k��@�Z�L4@�Ȱ���!?���"��@�1c�ٿ%B�k��@�Z�L4@�Ȱ���!?���"��@�1c�ٿ%B�k��@�Z�L4@�Ȱ���!?���"��@�1c�ٿ%B�k��@�Z�L4@�Ȱ���!?���"��@f�v@w�ٿ�|�A�@��?�}(4@���Ő!?u�LϢ��@f�v@w�ٿ�|�A�@��?�}(4@���Ő!?u�LϢ��@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@�ɀ�ݛٿ��>"[e�@���4@�|Ȼj�!?�o���)�@���ç�ٿpT��Y�@����X4@>���!?\Md373�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@砫��ٿ''���@��-
�%4@�v~�!?`)��B�@��^?S�ٿUxB�_�@�`$M�,4@��(�Đ!?G<H:z0�@��^?S�ٿUxB�_�@�`$M�,4@��(�Đ!?G<H:z0�@��^?S�ٿUxB�_�@�`$M�,4@��(�Đ!?G<H:z0�@��^?S�ٿUxB�_�@�`$M�,4@��(�Đ!?G<H:z0�@	��C�ٿ�4C�H�@L**%r�3@�V#���!?u�N��@	��C�ٿ�4C�H�@L**%r�3@�V#���!?u�N��@	��C�ٿ�4C�H�@L**%r�3@�V#���!?u�N��@-�B���ٿ�Ib����@�%��h�3@[�=�ǐ!?3�S-�@-�B���ٿ�Ib����@�%��h�3@[�=�ǐ!?3�S-�@��TrȠٿU������@�n�
A4@�JB	��!?��:
��@��TrȠٿU������@�n�
A4@�JB	��!?��:
��@��TrȠٿU������@�n�
A4@�JB	��!?��:
��@��TrȠٿU������@�n�
A4@�JB	��!?��:
��@��TrȠٿU������@�n�
A4@�JB	��!?��:
��@A���ǡٿ$r(	���@d���	4@=����!?�����@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@J�zs�ٿ1�v�J�@�Ւ~�3@����!?��h}�@$��ʠٿ�	�����@�N��a�3@\�e��!?��s����@$��ʠٿ�	�����@�N��a�3@\�e��!?��s����@$��ʠٿ�	�����@�N��a�3@\�e��!?��s����@R�L"^�ٿ�/�7��@�sy\)�3@�{��z�!?���v�~�@R�L"^�ٿ�/�7��@�sy\)�3@�{��z�!?���v�~�@ܼ[;��ٿ�f�G���@�x���3@��mM��!?6PCa)�@ܼ[;��ٿ�f�G���@�x���3@��mM��!?6PCa)�@ܼ[;��ٿ�f�G���@�x���3@��mM��!?6PCa)�@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@=L�ٚٿ�姬Lm�@��eR	 4@!�eqv�!?�N���@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@a1-F̜ٿRC�����@�|~ɺ4@h;*y�!? �8Ԇ��@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@7S��ٿ��O���@?�� b4@�k�Vz�!?ke�{�@d�=Cߖٿ���h�@}���`4@4�o�e�!?�9���@d�=Cߖٿ���h�@}���`4@4�o�e�!?�9���@d�=Cߖٿ���h�@}���`4@4�o�e�!?�9���@���6�ٿd�7���@~bl��4@�Ž���!?L���6�@���6�ٿd�7���@~bl��4@�Ž���!?L���6�@���6�ٿd�7���@~bl��4@�Ž���!?L���6�@H��T9�ٿ��Gp�@�-�v�C4@?�����!?�{�_Õ@H��T9�ٿ��Gp�@�-�v�C4@?�����!?�{�_Õ@H��T9�ٿ��Gp�@�-�v�C4@?�����!?�{�_Õ@H��T9�ٿ��Gp�@�-�v�C4@?�����!?�{�_Õ@�`Ȕ��ٿj�?�,�@�����(4@Tq�j�!?;q8
Ε@�`Ȕ��ٿj�?�,�@�����(4@Tq�j�!?;q8
Ε@�`Ȕ��ٿj�?�,�@�����(4@Tq�j�!?;q8
Ε@Y���	�ٿ�q3XI�@a�;��=4@666�!?/Jˆ�Օ@Y���	�ٿ�q3XI�@a�;��=4@666�!?/Jˆ�Օ@Y���	�ٿ�q3XI�@a�;��=4@666�!?/Jˆ�Օ@Y���	�ٿ�q3XI�@a�;��=4@666�!?/Jˆ�Օ@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@jL��(�ٿ|�K!{��@��m�>4@`M��A�!?[K⮾��@ޢ�nz�ٿ޾�gp��@����4@��0�}�!?��S�p�@ޢ�nz�ٿ޾�gp��@����4@��0�}�!?��S�p�@ޢ�nz�ٿ޾�gp��@����4@��0�}�!?��S�p�@Г�|��ٿ널�p�@n���54@#��v�!?�".�ە@Г�|��ٿ널�p�@n���54@#��v�!?�".�ە@Г�|��ٿ널�p�@n���54@#��v�!?�".�ە@��qG�ٿ6��a��@˷*0��3@����2�!?��4>:��@��qG�ٿ6��a��@˷*0��3@����2�!?��4>:��@��qG�ٿ6��a��@˷*0��3@����2�!?��4>:��@��qG�ٿ6��a��@˷*0��3@����2�!?��4>:��@�飈��ٿ�=�d]b�@O�#c4@�s;��!?H�4��@�飈��ٿ�=�d]b�@O�#c4@�s;��!?H�4��@�飈��ٿ�=�d]b�@O�#c4@�s;��!?H�4��@�飈��ٿ�=�d]b�@O�#c4@�s;��!?H�4��@�飈��ٿ�=�d]b�@O�#c4@�s;��!?H�4��@�nǎ*�ٿ����-�@�pN94@��g@�!?ph9�;�@�W�ʞ�ٿ�q��h�@�֛�3@��Y}_�!?�uH�ff�@�*�۳�ٿ���4��@튏Ax�3@Y>X��!?�`H��@�*�۳�ٿ���4��@튏Ax�3@Y>X��!?�`H��@�*�۳�ٿ���4��@튏Ax�3@Y>X��!?�`H��@(;ſ�ٿ)���*��@�g�(�3@	�`?2�!?AO0���@*�EK$�ٿ�}`�3��@ �\r�24@�^<��!?���ys�@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@������ٿ     ��@      4@�t><K�!?��=��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@ ;��ٿq�����@�M� 4@0i��l�!?5Ƒ3��@qD��ٿ��b����@��( 4@��Ɲ�!?�;����@qD��ٿ��b����@��( 4@��Ɲ�!?�;����@qD��ٿ��b����@��( 4@��Ɲ�!?�;����@qD��ٿ��b����@��( 4@��Ɲ�!?�;����@qD��ٿ��b����@��( 4@��Ɲ�!?�;����@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@����ٿC������@ŕr9 4@�>���!?��h���@\5��ٿ>�Q����@��Vk 4@�;2Ox�!?��cZ��@\5��ٿ>�Q����@��Vk 4@�;2Ox�!?��cZ��@���&�ٿxq�����@j�3i 4@	s~���!?�~ǃ��@���&�ٿxq�����@j�3i 4@	s~���!?�~ǃ��@���&�ٿxq�����@j�3i 4@	s~���!?�~ǃ��@���&�ٿxq�����@j�3i 4@	s~���!?�~ǃ��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@��I��ٿJ�����@wo7� 4@h�1es�!?�n+��@����ٿ�g�����@!;�Q 4@���Z�!?\�f��@����ٿ�g�����@!;�Q 4@���Z�!?\�f��@����ٿ�g�����@!;�Q 4@���Z�!?\�f��@��C8�ٿ�������@�
 4@�t� P�!?�(���@��C8�ٿ�������@�
 4@�t� P�!?�(���@��C8�ٿ�������@�
 4@�t� P�!?�(���@��C8�ٿ�������@�
 4@�t� P�!?�(���@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@��	\�ٿ=�~����@��q
 4@�2(���!?AWq ��@_����ٿD�����@<
/�	 4@ӡp���!?_����@_����ٿD�����@<
/�	 4@ӡp���!?_����@_����ٿD�����@<
/�	 4@ӡp���!?_����@�G}f�ٿ/������@��Q
 4@틳���!?�����@���ٿ�������@g5O
 4@�}��Y�!?�Z���@���ٿ�������@g5O
 4@�}��Y�!?�Z���@���ٿ�������@g5O
 4@�}��Y�!?�Z���@���ٿ�������@g5O
 4@�}��Y�!?�Z���@�_�c�ٿP7�����@_n
 4@�;�W�!?�K����@�_�c�ٿP7�����@_n
 4@�;�W�!?�K����@ҷ�ٿf������@��ǣ
 4@�;`Ԇ�!?>͔���@�n8�ٿu�(����@�*� 4@��v�!?Kr����@�n8�ٿu�(����@�*� 4@��v�!?Kr����@�n8�ٿu�(����@�*� 4@��v�!?Kr����@��L�ٿR�y����@z���
 4@g��ő�!?�p����@���d�ٿ�ѿ����@i&v- 4@j]�?��!?\m����@���d�ٿ�ѿ����@i&v- 4@j]�?��!?\m����@V��ٿ�[�����@@��g 4@;��C��!?y����@�F�1�ٿ;tW����@�v�0 4@=�c��!?�l����@�ԋ��ٿO������@
PR> 4@a��P�!?UE����@�ԋ��ٿO������@
PR> 4@a��P�!?UE����@ֵi�ٿ�������@�B�� 4@9rPn�!?���	��@�&��ٿi�!����@[{L1 4@��_�j�!?R����@�&��ٿi�!����@[{L1 4@��_�j�!?R����@����ٿl�����@�ö� 4@L�8��!?�<���@����ٿl�����@�ö� 4@L�8��!?�<���@����ٿl�����@�ö� 4@L�8��!?�<���@dCF��ٿ8����@p��� 4@�%�D��!?�p����@ ����ٿؑ����@��~� 4@Y�`l�!?�O=���@u�u� �ٿ簮����@�A�4 4@�HIe�!?@����@.��ٿ��>����@�l7� 4@ qY��!?Xq����@.��ٿ��>����@�l7� 4@ qY��!?Xq����@���ٿ~�����@���� 4@���NL�!?��1���@���ٿ~�����@���� 4@���NL�!?��1���@cS� �ٿ��p����@u� 4@U��l�!?$�����@cS� �ٿ��p����@u� 4@U��l�!?$�����@cS� �ٿ��p����@u� 4@U��l�!?$�����@cS� �ٿ��p����@u� 4@U��l�!?$�����@cS� �ٿ��p����@u� 4@U��l�!?$�����@X6���ٿ@�>����@]&C_ 4@�f�T�!?(�_���@�5O��ٿ�G�����@��K 4@khU�r�!?�����@@b�x �ٿ������@
͎� 4@�ԻZǐ!?��X���@@b�x �ٿ������@
͎� 4@�ԻZǐ!?��X���@@b�x �ٿ������@
͎� 4@�ԻZǐ!?��X���@/�8"�ٿ;>�����@>��" 4@��%@Ɛ!? �^���@���A%�ٿ),y����@��[) 4@�Wp�!?C�&���@���A%�ٿ),y����@��[) 4@�Wp�!?C�&���@��*�!�ٿ�fI����@��� 4@Y��2��!?NH���@`�b�$�ٿ�������@
ڬ  4@h��V<�!?;�����@.Zb7#�ٿ������@��� 4@7�N�o�!?�Ʋ���@:��>'�ٿ�f�����@�� 4@F�`�!?�Fs���@:��>'�ٿ�f�����@�� 4@F�`�!?�Fs���@��p,�ٿZ������@"p� 4@m,�q`�!?|�M���@��>(�ٿ-�����@��X 4@��H�!?*����@>�0'�ٿ�<,����@��Xv 4@;���h�!?�����@>�0'�ٿ�<,����@��Xv 4@;���h�!?�����@��u�#�ٿ52�����@T��� 4@ �苐!?NDu���@��u�#�ٿ52�����@T��� 4@ �苐!?NDu���@�cd$�ٿye�����@]�ֽ 4@|wEb�!?�  ���@�cd$�ٿye�����@]�ֽ 4@|wEb�!?�  ���@���"�ٿ������@n��  4@v�ah��!??�����@�Me"�ٿ� M����@c��� 4@��H���!?�5����@K�q�ٿ�<�����@	|Z 4@W�&.��!?�����@Ȧ��ٿ7�����@O	p% 4@s��Y�!?ݽ���@-o3��ٿuF�����@�� � 4@��<���!?�@���@|�p��ٿ�+�����@R#� 4@T��!?+B ���@|�p��ٿ�+�����@R#� 4@T��!?+B ���@vgLp �ٿv&R����@Qcv 4@~�{B��!?�w����@vgLp �ٿv&R����@Qcv 4@~�{B��!?�w����@��C!�ٿ6�����@m=� 4@Mys��!?�z��@�ZL��ٿ�������@)�# 4@ߞ]�t�!?~?���@!B�P�ٿ$������@��� 4@`��9��!?CӁ���@����ٿ� ����@�#Q� 4@��m�Ő!?q�o���@"��ٿ��T����@N�G� 4@��/�'�!?��Ԩ��@;���ٿR����@�ޟ 4@��� �!?�R����@\=K��ٿ��t����@p*)� 4@[#!e�!?�{����@\=K��ٿ��t����@p*)� 4@[#!e�!?�{����@(��S�ٿ'~�����@�A'I 4@�f#i�!?��:���@(��S�ٿ'~�����@�A'I 4@�f#i�!?��:���@�G���ٿ�~�����@��P 4@��Ր!?�d6���@�G���ٿ�~�����@��P 4@��Ր!?�d6���@jށ �ٿ������@"�QF 4@�f�!?{^���@��e�ٿ�������@��� 4@?"i�C�!?��D���@)�V+�ٿ������@L%E: 4@y���}�!?yoΎ��@)�V+�ٿ������@L%E: 4@y���}�!?yoΎ��@�m)�ٿ�������@��o> 4@��ǀb�!?Cٗ��@�m)�ٿ�������@��o> 4@��ǀb�!?Cٗ��@����ٿ|������@��<� 4@7Pru]�!?�Q���@ö$�!�ٿFP����@P<L� 4@�:"�!?�V���@���$�ٿ-����@�Z� 4@h�E�A�!?�����@���$�ٿ-����@�Z� 4@h�E�A�!?�����@<�#"�ٿ�������@c�� 4@�D6�U�!?+2�{��@Vt��ٿ�N�����@o�J
 4@�ds���!?��c���@��[w#�ٿ�a`����@,�� 4@��/N��!?��T���@��[w#�ٿ�a`����@,�� 4@��/N��!?��T���@�I�#�ٿ>Y�����@4�� 4@��M���!?w(���@Stq��ٿ0>�����@�� 4@8�)Dx�!?p�[���@����ٿ'������@|D� 4@� V��!?�����@�z��!�ٿC������@&��� 4@�9�6��!?3�����@
��V$�ٿ�%����@��� 4@���dĐ!?_����@ٓ�.$�ٿD������@/!� 4@N�@|��!?:q���@�O�"�ٿUpj����@���� 4@=%F�]�!?zE����@�3#>"�ٿ&������@���� 4@!0L�!?��[���@wL!� �ٿ�������@���� 4@��^%T�!?79���@|����ٿ������@8-~� 4@��j�!?
����@yc���ٿ������@�K} 4@�N�B�!?(�]���@�#z��ٿwo�����@&�< 4@�����!?$r����@�#z��ٿwo�����@&�< 4@�����!?$r����@s��R�ٿ�%�����@S��
 4@6�S�!?��.���@���d�ٿ������@����
 4@���uQ�!?��P���@+ �ٿ⿧����@Ƥ0�
 4@�A/�!?�6Ř��@�w���ٿNGH����@2#��
 4@"ݯ+�!?Y2����@���ٿ]�7����@��
 4@��d�
�!?�j���@`"��ٿ�������@�pZs
 4@=
��.�!?�N܏��@#����ٿ�G*����@�U
 4@�X�2'�!?O����@#����ٿ�G*����@�U
 4@�X�2'�!?O����@#����ٿ�G*����@�U
 4@�X�2'�!?O����@#����ٿ�G*����@�U
 4@�X�2'�!?O����@H7���ٿ������@>m��
 4@&�z$�!?�ێc��@�\{�ٿ������@s~��
 4@x�l���!?>�vh��@2���ٿ
x����@@ˀv
 4@���!?��M��@r|k��ٿ�ya����@�Q�B
 4@�xz0�!?O��1��@��Ԍ�ٿ�������@P�
 4@�F�j�!?n��e��@ۧ�#"�ٿ�.����@�|.�
 4@�J�\��!?=��_��@h n$�ٿr:����@�u�
 4@�!�J��!?���E��@��Q�'�ٿ�E�����@WQ4� 4@��٩��!?��g��@��Q�'�ٿ�E�����@WQ4� 4@��٩��!?��g��@4��(�ٿ�I����@�]�� 4@��ސ�!?qҡ���@��<&�ٿ��5����@�E0 4@��␐!?�}����@��<&�ٿ��5����@�E0 4@��␐!?�}����@5�+�%�ٿ������@pù  4@A����!?^@]v��@m�V!�ٿ�g�����@��w 4@�~�ǐ!?��j��@m�V!�ٿ�g�����@��w 4@�~�ǐ!?��j��@�KFq �ٿ�����@Gea�
 4@K�͐!?�%uh��@�rbM�ٿ�E�����@xD�3
 4@�[���!??)�b��@�o�b�ٿL ����@�B�	 4@��c�!?{Y��@״���ٿ��U����@@3z�	 4@=z��k�!?�,�X��@״���ٿ��U����@@3z�	 4@=z��k�!?�,�X��@�zm�ٿy)T����@+2� 4@�{N�F�!?�!*��@!�Y�ٿ�	f����@�r 4@E3'�Y�!?F׳5��@�j�u#�ٿ�9�����@�G�<	 4@��؈d�!?�7:��@�j�u#�ٿ�9�����@�G�<	 4@��؈d�!?�7:��@�N[� �ٿ�������@�ob(	 4@T eN�!?�|F��@�N[� �ٿ�������@�ob(	 4@T eN�!?�|F��@�N[� �ٿ�������@�ob(	 4@T eN�!?�|F��@�N[� �ٿ�������@�ob(	 4@T eN�!?�|F��@]�e�"�ٿ������@y�ks 4@��MW�!?(��,��@��G!$�ٿ�����@,sQ� 4@�+� �!?�ϖ��@��m�'�ٿ������@�F2	 4@�P�Q�!?�9��@& ��$�ٿ *����@&t��	 4@����X�!?�G��@�.��%�ٿ�*�����@B��
 4@���CT�!? b�M��@�d��+�ٿ:�����@�!T! 4@���::�!?��C��@��'�&�ٿ�����@�䷁ 4@�]��b�!?3�Um��@��*;$�ٿ��h����@�-�& 4@� \�!?���}��@�ӣ�!�ٿ������@�q� 4@R#��!�!?�@���@�ӣ�!�ٿ������@�q� 4@R#��!�!?�@���@�ӣ�!�ٿ������@�q� 4@R#��!�!?�@���@K��%�ٿ��l����@AʰJ 4@�ƾ��!?�l����@ع?q(�ٿ�8�����@R�BC 4@z~��Ð!?
K���@ع?q(�ٿ�8�����@R�BC 4@z~��Ð!?
K���@��@]'�ٿ�����@QgY 4@��/��!?�Mh���@��@]'�ٿ�����@QgY 4@��/��!?�Mh���@����ٿRâ����@�D׋ 4@£����!?l26���@����ٿRâ����@�D׋ 4@£����!?l26���@sT�"�ٿ~?�����@v*2� 4@��o��!?�˟��@�	��$�ٿ�B����@���j 4@���&_�!?+�w��@ o��"�ٿ�������@�.�� 4@�1��|�!?�_~��@�D��ٿ������@��Zl 4@x�E�Y�!?�-�~��@\'И!�ٿ�-e����@�d� 4@�m�0N�!?�e�S��@~L�(�ٿ3������@���
 4@&Q�|�!?��@��@�.�)�ٿYj����@��/
 4@V3�CM�!?`'����@�/a1�ٿ.�U����@��2	 4@��k`�!?̧v���@l4��.�ٿ�c�����@Dhi: 4@�ј��!?;Hʵ��@l4��.�ٿ�c�����@Dhi: 4@�ј��!?;Hʵ��@l4��.�ٿ�c�����@Dhi: 4@�ј��!?;Hʵ��@�}l�3�ٿ��ʪ���@���	 4@^�����!?�*���@�}l�3�ٿ��ʪ���@���	 4@^�����!?�*���@�[��2�ٿ�������@�@� 4@Ht\���!?�,}��@cSl5�ٿKټ����@�Q�g 4@?�8���!?�����@*��1�ٿ�������@w�xb 4@��P��!?�����@*��1�ٿ�������@w�xb 4@��P��!?�����@��ZR.�ٿAx�����@�^Q� 4@�5+^�!?G8=��@ȩ&�ٿ�3K����@r`. 4@Ze9���!?�&N��@�-;��ٿl�t����@ol�0 4@���<�!?r����@����ٿQH����@�ޠ 4@��eW�!?6����@����ٿQH����@�ޠ 4@��eW�!?6����@$���ٿ�&� ��@3`�� 4@�Ƹj<�!?��2��@fX��ٿ[~�	 ��@�Y 4@b��.g�!?�	?8��@(mZ��ٿ��A ��@(��7 4@�At\�!?���:��@��ٿ�q=����@��� 4@(��=��!?3����@]�� �ٿH�����@媇� 4@��~Hb�!?J�����@]�� �ٿH�����@媇� 4@��~Hb�!?J�����@�;�(�ٿ�,*����@��! 4@�3����!?iC���@9��/�ٿY�6����@��V� 4@����]�!?��%��@Y��-0�ٿ�C����@W�? 4@~g�x�!?=L��@T��:�ٿ�Ŏ����@'A�� 4@�Ѝ!?��*��@mWۭA�ٿ�����@�M�� 4@�p�[�!?K����@mWۭA�ٿ�����@�M�� 4@�p�[�!?K����@U_�H=�ٿH�S����@�,�� 4@��:R�!?T��]��@�%�L�ٿ��� ��@���= 4@�
��U�!?.����@QCȑ[�ٿ��C ��@5�2� 4@/8a�!?+��v��@Q"i�ٿ�� ��@��r 4@&z/���!?�e���@Q"i�ٿ�� ��@��r 4@&z/���!?�e���@ɳ�Nk�ٿu� ��@ܾ�� 4@4NBJ�!?��Hb��@[���q�ٿ�� ��@�`ڌ 4@�J�^�!?e���@|�\�o�ٿ��%# ��@Ӥ��  4@`8x�!?���*��@B֖0��ٿF��( ��@S[�& 4@�)q�j�!?i�>���@�� &��ٿ���8 ��@	Mj/ 4@��jh�!?@`���@̮K���ٿfz�J ��@�!^- 4@81k@T�!?)�[���@̮K���ٿfz�J ��@�!^- 4@81k@T�!?)�[���@̮K���ٿfz�J ��@�!^- 4@81k@T�!?)�[���@�U� ��ٿ΢�j ��@��(2 4@60N2�!?�E
��@Hc��ٿn�	� ��@�e�K 4@ w�:�!?���G��@6���G�ٿ��6� ��@!���Y 4@�r")!�!?���O��@6���G�ٿ��6� ��@!���Y 4@�r")!�!?���O��@6���G�ٿ��6� ��@!���Y 4@�r")!�!?���O��@l>P>�ٿ�9���@;� � 4@F�)i�!?�S����@�Q�$O�ٿ�^����@�X8 � 4@1)���!?��3v��@@Sl���ٿnV�\��@��&� 4@g����!?�LO���@��s�ٿS�?��@��.k 4@�r���!?}�����@a@P+əٿv�� ��@1�&]; 4@�`qL�!?�L��@a@P+əٿv�� ��@1�&]; 4@�`qL�!?�L��@$#��ٿΙ�����@�\[���3@'�Ǥ9�!?��vl��@$#��ٿΙ�����@�\[���3@'�Ǥ9�!?��vl��@-�]��ٿ&!�J���@nڦ��3@��mRW�!?��kE��@5�i^&�ٿ�����@�G�p
 4@��H�!?"(R)��@�򻋘ٿPe����@��5��3@?����!?0��-��@����ٿΕ;���@g�����3@�����!?7�p ��@�|^'��ٿ�[Op���@3�!��3@�+f_�!?hO1���@�*aŃ�ٿ�T>���@��F��3@s��i�!?b����@*��8T�ٿ��c����@mQ)� 4@3!���!?���	��@�̊@Ԙٿ�VwG���@�����3@�zٺ�!?K_���@Z��>�ٿ�	�����@̣r| 4@�χĹ�!?��$��@m@[��ٿ�HYL���@A����3@�FP7�!?��|��@aᅙٿ>s����@�0* 4@Kh:��!?Z����@Ƽ�
�ٿH����@�YN� 4@M�_׊�!?^S]��@Ƽ�
�ٿH����@�YN� 4@M�_׊�!?^S]��@�D����ٿ���6��@W>4�r 4@f�>6��!?������@W��M�ٿa]����@��Rp� 4@�F��q�!?j��	��@^����ٿ�D� ��@�!Lg 4@uM���!?)��p��@^����ٿ�D� ��@�!Lg 4@uM���!?)��p��@^����ٿ�D� ��@�!Lg 4@uM���!?)��p��@� ^t��ٿ������@�CK��3@�f�X�!?Sd����@� ^t��ٿ������@�CK��3@�f�X�!?Sd����@� ^t��ٿ������@�CK��3@�f�X�!?Sd����@�@B�/�ٿIꊆ ��@s~p�L 4@ ��*�!?PKĤ��@� D���ٿ�Aw ��@�:.�3 4@`%�_	�!?W�gg��@� D���ٿ�Aw ��@�:.�3 4@`%�_	�!?W�gg��@�/F�:�ٿ������@�y_u 4@3��g��!?�Q���@�/F�:�ٿ������@�y_u 4@3��g��!?�Q���@��0��ٿ9������@���
 4@<��b_�!?��f��@@);%�ٿ����@K� �� 4@:��Xb�!?mݪF��@@);%�ٿ����@K� �� 4@:��Xb�!?mݪF��@@);%�ٿ����@K� �� 4@:��Xb�!?mݪF��@�>�k�ٿ��*���@�}�1� 4@DR�u�!?�A����@g�ͳI�ٿ8|���@� �� 4@=�|�R�!?�eW��@���j6�ٿ9����@b@��'4@�P{�!?��A��@;Ȉ;�ٿ�Y���@����� 4@r��cv�!?�S���@��
�ٿ�n����@�G��� 4@�O���!?�����@�?�?�ٿu�����@�����3@(��p�!?�i���@Pr����ٿ�����@G�h4@�Vz@�!?ȸѨ��@ �X=�ٿ�G^���@Z��� 4@jy;�d�!?�ݵ?��@������ٿ$�#��@�-�E4@���o�!?��7���@���lm�ٿ��D���@�(�-� 4@d�͋K�!?pg��@���lm�ٿ��D���@�(�-� 4@d�͋K�!?pg��@2y(B�ٿ��L���@��sb� 4@Y_q?�!?=����@߀�%�ٿi,���@�x� 4@
1h�i�!?Ec1S��@X����ٿr�����@�v	���3@��V�!?���-��@tz��v�ٿ��#b���@1Y�u*�3@i�Om�!?`ҕv��@tz��v�ٿ��#b���@1Y�u*�3@i�Om�!?`ҕv��@tz��v�ٿ��#b���@1Y�u*�3@i�Om�!?`ҕv��@tz��v�ٿ��#b���@1Y�u*�3@i�Om�!?`ҕv��@tz��v�ٿ��#b���@1Y�u*�3@i�Om�!?`ҕv��@�&ʚٿ��V���@a/3�� 4@��d�!?
�����@�b͡$�ٿ�M.���@|j�y04@��|2�!?��n��@�b͡$�ٿ�M.���@|j�y04@��|2�!?��n��@�)�t��ٿ�G����@0��T�4@��B�V�!?�Q:���@�)�t��ٿ�G����@0��T�4@��B�V�!?�Q:���@�)�t��ٿ�G����@0��T�4@��B�V�!?�Q:���@:n����ٿ�G����@Z�=&84@:����!?�ao��@:n����ٿ�G����@Z�=&84@:����!?�ao��@�p�%�ٿu���@���z 4@M��!?�v��@ԍ���ٿWBJ��@�A��!4@���t�!?N����@ԍ���ٿWBJ��@�A��!4@���t�!?N����@�>ߗٿecTO���@x^i��3@P�:p��!?ʲ�&��@�>ߗٿecTO���@x^i��3@P�:p��!?ʲ�&��@�>ߗٿecTO���@x^i��3@P�:p��!?ʲ�&��@��e���ٿNj�y��@��� 4@P�M�d�!?K���@o��.��ٿ��;���@�`�f 4@�f�$�!?A�b��@o��.��ٿ��;���@�`�f 4@�f�$�!?A�b��@���
D�ٿN���@�jG�( 4@���S�!?M���@�m	��ٿΜ�:��@��e�� 4@��h��!?yK�;��@�m	��ٿΜ�:��@��e�� 4@��h��!?yK�;��@�m	��ٿΜ�:��@��e�� 4@��h��!?yK�;��@�m	��ٿΜ�:��@��e�� 4@��h��!?yK�;��@��ٿ	7Y	��@H����4@TR����!?�����@�<�Q��ٿC%���@ܝ��4@�g�F�!?�(�|��@S0����ٿ�VL���@�B�� 4@Fs��c�!?�!
f��@S0����ٿ�VL���@�B�� 4@Fs��c�!?�!
f��@S0����ٿ�VL���@�B�� 4@Fs��c�!?�!
f��@�꥜ŞٿiO����@�O@,�4@�b��4�!?�k�~��@�D�wĞٿ�&n��@�t���4@Sy����!?�wR��@�D�wĞٿ�&n��@�t���4@Sy����!?�wR��@�D�wĞٿ�&n��@�t���4@Sy����!?�wR��@��JיٿU�p ��@aA�5 4@�h���!?�2����@��JיٿU�p ��@aA�5 4@�h���!?�2����@#u��ٿ�[��@, ~�4@��[�!?�K���@�	�S��ٿ�|�����@�ġ�g�3@r�$�-�!?�2�E��@��d-��ٿU'����@3�+&��3@�����!?_�����@=�ZI_�ٿ�{ә ��@�����3@ή�mԐ!?��t���@=�ZI_�ٿ�{ә ��@�����3@ή�mԐ!?��t���@=�ZI_�ٿ�{ә ��@�����3@ή�mԐ!?��t���@=�ZI_�ٿ�{ә ��@�����3@ή�mԐ!?��t���@��7���ٿ|[� ��@+�=�� 4@k2�{��!?�����@���M�ٿ�-���@B�!X\4@��e���!?��A��@���M�ٿ�-���@B�!X\4@��e���!?��A��@2O����ٿH]����@�ʧ�z4@�L���!?�l���@��:ԝٿuM�����@~���� 4@ǅ�N[�!?V1��@��:ԝٿuM�����@~���� 4@ǅ�N[�!?V1��@��:ԝٿuM�����@~���� 4@ǅ�N[�!?V1��@�I�SA�ٿ2R���@�s>r  4@��%5�!?܂T��@����ٿQ�s���@  ��� 4@�޷�!?p�e���@(#����ٿ������@�V��4@+�Lޏ!?�bX��@TK:�¡ٿȪ����@��Â�4@5�n͏!?������@��1���ٿ��2����@���� 4@T����!?\j%+��@�dM��ٿ] ����@��Y�D 4@�Ё�!?�}w^��@˛�N�ٿ@������@�爐��3@jI���!?�jy��@˛�N�ٿ@������@�爐��3@jI���!?�jy��@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@�e5���ٿ������@�$KB��3@�<H���!?�����@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@jiF<�ٿ(�'��@4��64@��ξ�!?��/��@���ge�ٿ��F��@[� �4@�߬��!?|�w���@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@)|�l�ٿ� x���@RQEY�4@H�F7��!?qX����@%Q�9�ٿ�/��@�֨|%4@�􍡋�!? 3���@��f$��ٿ�%6Q��@��x�j4@�����!? Խ)��@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@4�m�ٿDv����@�V�0E 4@�k��L�!?	0���@����b�ٿ���	��@�Z*�4@x�/��!?7�i��@����b�ٿ���	��@�Z*�4@x�/��!?7�i��@��8q�ٿIP����@#����3@��8��!?��(��@��8q�ٿIP����@#����3@��8��!?��(��@��8q�ٿIP����@#����3@��8��!?��(��@��8q�ٿIP����@#����3@��8��!?��(��@"���ٿ��EQ܇�@)xg�(�3@6H{��!?���in�@�CB��ٿG�ه�@+�����3@��U"��!?��c}�@�CB��ٿG�ه�@+�����3@��U"��!?��c}�@�CB��ٿG�ه�@+�����3@��U"��!?��c}�@�CB��ٿG�ه�@+�����3@��U"��!?��c}�@�CB��ٿG�ه�@+�����3@��U"��!?��c}�@�#b^�ٿ�6_�Ƈ�@\�F �3@4�;&X�!?�k�^S�@�k�y_�ٿ�V)���@3t�d��3@Bp���!?}V誦�@�k�y_�ٿ�V)���@3t�d��3@Bp���!?}V誦�@����r�ٿ���=��@s�;H�3@h�h�ʐ!?�>���@����r�ٿ���=��@s�;H�3@h�h�ʐ!?�>���@�Im���ٿ���}ԇ�@�����3@�>��!?��뛎�@�Im���ٿ���}ԇ�@�����3@�>��!?��뛎�@Ty2�ٿ4*���@�Z3>u�3@�[�]�!?"*Љ��@�w�=��ٿ�ˣ���@�j��7�3@�	��!?� ,U��@�w�=��ٿ�ˣ���@�j��7�3@�	��!?� ,U��@,��pp�ٿD�>އ�@C{�%�3@XK�{�!?FyUy�@9e��ġٿqP�(ʇ�@I�{o*�3@G�D)��!?Bx��L�@9e��ġٿqP�(ʇ�@I�{o*�3@G�D)��!?Bx��L�@9e��ġٿqP�(ʇ�@I�{o*�3@G�D)��!?Bx��L�@9e��ġٿqP�(ʇ�@I�{o*�3@G�D)��!?Bx��L�@�Ȏ�D�ٿݩ�ч�@�9����3@j�J ��!?�vb.e�@�Ȏ�D�ٿݩ�ч�@�9����3@j�J ��!?�vb.e�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@C~F��ٿ�0f����@�~D��3@p���h�!?CJG�.�@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@3���2�ٿ������@�"
��3@yG��`�!?þÓ��@	��Νٿ����G��@k��q_�3@��u�[�!?�(�u�@�F��؟ٿR��h��@��R���3@f{��m�!?����@�՚f�ٿB�����@~�6��3@�흇��!?�����@�՚f�ٿB�����@~�6��3@�흇��!?�����@�՚f�ٿB�����@~�6��3@�흇��!?�����@�՚f�ٿB�����@~�6��3@�흇��!?�����@�՚f�ٿB�����@~�6��3@�흇��!?�����@�՚f�ٿB�����@~�6��3@�흇��!?�����@���M�ٿc��@��@����;�3@#E)�b�!?g����@����ٿ�5f��@XtS��3@�W��!?U������@����ٿ�5f��@XtS��3@�W��!?U������@ ��GO�ٿ^JK���@��zj�3@��*q�!?�j6>��@ ��GO�ٿ^JK���@��zj�3@��*q�!?�j6>��@ ��GO�ٿ^JK���@��zj�3@��*q�!?�j6>��@�C8U�ٿ�>�'/��@�L��֡3@�*w@P�!?|�����@�C8U�ٿ�>�'/��@�L��֡3@�*w@P�!?|�����@�C8U�ٿ�>�'/��@�L��֡3@�*w@P�!?|�����@˒+��ٿ�`#;��@�*���3@��HD�!?���}��@˒+��ٿ�`#;��@�*���3@��HD�!?���}��@˒+��ٿ�`#;��@�*���3@��HD�!?���}��@˒+��ٿ�`#;��@�*���3@��HD�!?���}��@˒+��ٿ�`#;��@�*���3@��HD�!?���}��@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@#8�p�ٿ,��fˆ�@`�
��3@V}P�!?�Q��� �@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@�l��ٿ安{C��@�GB���3@dt���!?A����@����Y�ٿ��>/,��@,$���3@؛Gx��!?����@x���ĕٿ��Y힇�@������3@�f.}��!?���@KN�4��ٿ�X�����@1_~5� 4@��U�!? ��nl�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@GC5���ٿ��Mb��@�����3@��J�*�!?©G�U�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@� G��ٿ"�a�ɇ�@������3@Y�#^�!?���CW�@"J	p�ٿuå���@�J�z��3@��Fy�!?����@"J	p�ٿuå���@�J�z��3@��Fy�!?����@"J	p�ٿuå���@�J�z��3@��Fy�!?����@"J	p�ٿuå���@�J�z��3@��Fy�!?����@"J	p�ٿuå���@�J�z��3@��Fy�!?����@"J	p�ٿuå���@�J�z��3@��Fy�!?����@�n�M��ٿw��Έ�@*�c�O4@iz}�!?~|<���@��<]^�ٿ?���އ�@x�����3@��͸P�!?���f�@��<]^�ٿ?���އ�@x�����3@��͸P�!?���f�@��<]^�ٿ?���އ�@x�����3@��͸P�!?���f�@��<]^�ٿ?���އ�@x�����3@��͸P�!?���f�@��<]^�ٿ?���އ�@x�����3@��͸P�!?���f�@�g�y�ٿ+_�����@�̃� 4@�~�y�!?K.��V�@�g�y�ٿ+_�����@�̃� 4@�~�y�!?K.��V�@�g�y�ٿ+_�����@�̃� 4@�~�y�!?K.��V�@�$/��ٿ"��?6��@�v���3@.~�Wk�!?cj&X��@�$/��ٿ"��?6��@�v���3@.~�Wk�!?cj&X��@e�~%�ٿ���Ɉ�@�K���4@���l�!?�U���@ƕ ��ٿ�u�Q��@7k*�H4@Q�o��!?�N�v	�@ƕ ��ٿ�u�Q��@7k*�H4@Q�o��!?�N�v	�@ƕ ��ٿ�u�Q��@7k*�H4@Q�o��!?�N�v	�@ƕ ��ٿ�u�Q��@7k*�H4@Q�o��!?�N�v	�@ƕ ��ٿ�u�Q��@7k*�H4@Q�o��!?�N�v	�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@C�'!Q�ٿ�Ñ%@��@��#@
4@�P���!?N�t�l�@���_`�ٿ�Ěc���@HY`��3@��u�P�!?����K�@���_`�ٿ�Ěc���@HY`��3@��u�P�!?����K�@���_`�ٿ�Ěc���@HY`��3@��u�P�!?����K�@���_`�ٿ�Ěc���@HY`��3@��u�P�!?����K�@�ı��ٿ��W����@@g��44@%=�<�!?ؖ�ժ�@�M�W�ٿחhL��@,��	O4@�l��֏!?X+�Y�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@��C.�ٿvw��R��@�ے��N4@��O��!?�>�N�	�@�.���ٿӵ!_`��@_sy2R4@]�~��!?��"�	�@�.���ٿӵ!_`��@_sy2R4@]�~��!?��"�	�@=b��L�ٿ�r�ʕ��@��י��3@�'��!?�&��e �@p=�a�ٿ���1~��@��~�(�3@�Y뗐!?;g	10 �@p=�a�ٿ���1~��@��~�(�3@�Y뗐!?;g	10 �@G��CҙٿA)�BA��@����f�3@L.!�{�!?Dܔ)�@�����ٿ��p�e��@&ON��Q4@a�93�!?j��:�	�@1�t�أٿD8g>p��@�M���3@���n�!?i|��d�@1�t�أٿD8g>p��@�M���3@���n�!?i|��d�@1�t�أٿD8g>p��@�M���3@���n�!?i|��d�@h��3��ٿ��[ꊇ�@O�[s.�3@�.s��!?S�ś�@h��3��ٿ��[ꊇ�@O�[s.�3@�.s��!?S�ś�@k���ٿ��2!��@������3@'̷���!?To���@k���ٿ��2!��@������3@'̷���!?To���@k���ٿ��2!��@������3@'̷���!?To���@k���ٿ��2!��@������3@'̷���!?To���@k���ٿ��2!��@������3@'̷���!?To���@a��^h�ٿ�k���@�|�r/E4@��_���!?����@a��^h�ٿ�k���@�|�r/E4@��_���!?����@a��^h�ٿ�k���@�|�r/E4@��_���!?����@�6��ٿ�����@��84@��7Ԥ�!?�0h���@�6��ٿ�����@��84@��7Ԥ�!?�0h���@�6��ٿ�����@��84@��7Ԥ�!?�0h���@�6��ٿ�����@��84@��7Ԥ�!?�0h���@�6��ٿ�����@��84@��7Ԥ�!?�0h���@�(� �ٿ=���ى�@���'@4@ ����!?��Dp�@�(� �ٿ=���ى�@���'@4@ ����!?��Dp�@�(� �ٿ=���ى�@���'@4@ ����!?��Dp�@�(� �ٿ=���ى�@���'@4@ ����!?��Dp�@���U�ٿ���q���@Ƨ��1�3@i���H�!?�~<��@���U�ٿ���q���@Ƨ��1�3@i���H�!?�~<��@���U�ٿ���q���@Ƨ��1�3@i���H�!?�~<��@���U�ٿ���q���@Ƨ��1�3@i���H�!?�~<��@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@?���ٿ�N���@'E��) 4@/_���!?�0hٝ�@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@�]W��ٿ�d�e���@�_Ӡ�4@���(q�!?�{���@��6��ٿ�B��Ƈ�@��7��3@0�Oni�!?�ͦ>[�@��6��ٿ�B��Ƈ�@��7��3@0�Oni�!?�ͦ>[�@��6��ٿ�B��Ƈ�@��7��3@0�Oni�!?�ͦ>[�@��6��ٿ�B��Ƈ�@��7��3@0�Oni�!?�ͦ>[�@��6��ٿ�B��Ƈ�@��7��3@0�Oni�!?�ͦ>[�@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@]��X�ٿ�k����@���$�3@��p�!?��[��@Hs*���ٿx�˚Ƈ�@�ۖTf�3@�_b���!?R�#�@Hs*���ٿx�˚Ƈ�@�ۖTf�3@�_b���!?R�#�@Hs*���ٿx�˚Ƈ�@�ۖTf�3@�_b���!?R�#�@Hs*���ٿx�˚Ƈ�@�ۖTf�3@�_b���!?R�#�@Hs*���ٿx�˚Ƈ�@�ۖTf�3@�_b���!?R�#�@��!+�ٿ1Nsb��@Zӽ �3@���W��!?��X� �@��!+�ٿ1Nsb��@Zӽ �3@���W��!?��X� �@�z꜖ٿӂ�6���@���3@��1;�!?:�Pj �@�z꜖ٿӂ�6���@���3@��1;�!?:�Pj �@�z꜖ٿӂ�6���@���3@��1;�!?:�Pj �@�z꜖ٿӂ�6���@���3@��1;�!?:�Pj �@��>��ٿc�Sܣ��@Q˧Oi�3@|�ז�!?m�#[ �@��>��ٿc�Sܣ��@Q˧Oi�3@|�ז�!?m�#[ �@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@E���}�ٿ��,�W��@��R��	4@V(�v�!?n*m��@����F�ٿ�=#t6��@E��F��3@�ZE���!?���Ö�@�@���ٿo�2��@����14@ezސ!?��\���@΁���ٿ9@��@�|���3@E;'�t�!?�#��*�@΁���ٿ9@��@�|���3@E;'�t�!?�#��*�@9��sŠٿJG�I��@���4�3@��^���!?�֦���@ܟh}�ٿ�?잆�@,�dW�3@զT�0�!?:e���@ܟh}�ٿ�?잆�@,�dW�3@զT�0�!?:e���@%�+ٗٿy|R���@�zR��3@�K_�!?%�iL��@�IϽ�ٿˮ��l��@X#q{��3@�A��V�!?�w���@�IϽ�ٿˮ��l��@X#q{��3@�A��V�!?�w���@�IϽ�ٿˮ��l��@X#q{��3@�A��V�!?�w���@6��+��ٿN]��?��@끴Z�3@�x�v�!?/!FX��@6��+��ٿN]��?��@끴Z�3@�x�v�!?/!FX��@6��+��ٿN]��?��@끴Z�3@�x�v�!?/!FX��@6��+��ٿN]��?��@끴Z�3@�x�v�!?/!FX��@6��+��ٿN]��?��@끴Z�3@�x�v�!?/!FX��@�_X��ٿ��al'��@cq�g��3@���h�!?J���@�_X��ٿ��al'��@cq�g��3@���h�!?J���@�_X��ٿ��al'��@cq�g��3@���h�!?J���@�_X��ٿ��al'��@cq�g��3@���h�!?J���@�_X��ٿ��al'��@cq�g��3@���h�!?J���@��z�̕ٿʋuL%��@��%
�=4@'�yސ!?D��՞	�@�'��ٿ��G��@�`�EnP4@��́��!?��I|	�@�'��ٿ��G��@�`�EnP4@��́��!?��I|	�@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@ŀb�ٿO5}�7��@9��|��3@&�c��!?�!�)��@����G�ٿ��	gE��@0����'4@��Ƞ��!?���6�@9�ٿgx�P���@�	��4@5�lbg�!?���xq�@9�ٿgx�P���@�	��4@5�lbg�!?���xq�@#��Z�ٿD����@Ι��3@��X�!?�q����@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�Lb��ٿ�/�E��@���4@�,��$�!?@T���@�hߋ��ٿ�6���@��3�,X4@���ѐ!?�Xb��@�hߋ��ٿ�6���@��3�,X4@���ѐ!?�Xb��@�hߋ��ٿ�6���@��3�,X4@���ѐ!?�Xb��@�hߋ��ٿ�6���@��3�,X4@���ѐ!?�Xb��@� Н�ٿi����@��}M4@`#FvƐ!?�L����@� Н�ٿi����@��}M4@`#FvƐ!?�L����@� Н�ٿi����@��}M4@`#FvƐ!?�L����@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@Kϊ�ٿ�*�Ѫ��@磁m�4@����*�!?������@����ٿ��ZB���@
�7��4@*�_�^�!?���a�@����ٿ��ZB���@
�7��4@*�_�^�!?���a�@����ٿ��ZB���@
�7��4@*�_�^�!?���a�@����ٿ��ZB���@
�7��4@*�_�^�!?���a�@����ٿ��ZB���@
�7��4@*�_�^�!?���a�@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@��
��ٿ�ys�ň�@���Z4@��صD�!?�f� �@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@���&��ٿ'��QV��@Zn���3@�o��]�!?A����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@�]���ٿ���ۇ�@����3@�� ��!?�����@>1�z��ٿ�Pɂ{��@�E[�4@���u�!?��	�S�@>1�z��ٿ�Pɂ{��@�E[�4@���u�!?��	�S�@>1�z��ٿ�Pɂ{��@�E[�4@���u�!?��	�S�@>1�z��ٿ�Pɂ{��@�E[�4@���u�!?��	�S�@$��¦ٿ��|���@-z�3@��k�1�!?0{j�7�@G�)��ٿ1:D(���@mLp�3@7�JG�!?��Ly� �@G�)��ٿ1:D(���@mLp�3@7�JG�!?��Ly� �@5�4A�ٿ�g^��@F49j4@�د�!?��g �@�=�ڛٿܚ@y���@xҍ=i4@��!?;2Gs	�@�=�ڛٿܚ@y���@xҍ=i4@��!?;2Gs	�@�=�ڛٿܚ@y���@xҍ=i4@��!?;2Gs	�@�=�ڛٿܚ@y���@xҍ=i4@��!?;2Gs	�@�=�ڛٿܚ@y���@xҍ=i4@��!?;2Gs	�@��gŠٿ��y��@�]&f�3@#�o� �!?O��@��gŠٿ��y��@�]&f�3@#�o� �!?O��@��gŠٿ��y��@�]&f�3@#�o� �!?O��@��gŠٿ��y��@�]&f�3@#�o� �!?O��@X2�E]�ٿ/���$��@��Ո��3@�[��O�!?��y�Z�@X2�E]�ٿ/���$��@��Ո��3@�[��O�!?��y�Z�@X2�E]�ٿ/���$��@��Ո��3@�[��O�!?��y�Z�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@o���ٿ->��=��@!fߢ4@����d�!?�,�:�@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@@�Q���ٿǮ�����@�2�n�4@\F��!?�M4��@Em�/�ٿ�k�i��@t5h�k�3@&�i�&�!?�?PD��@��Ɋ�ٿh�m#�@UF	4@�<}�!?  \���@��Ɋ�ٿh�m#�@UF	4@�<}�!?  \���@��"��ٿ��;��y�@�/��-�3@~��OF�!?c�ځ�Ԗ@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@�\��ٿ�_�e3��@[���4@���g�!?�|8���@#�rq�ٿ��f��@��7���3@MFM��!?d	����@#�rq�ٿ��f��@��7���3@MFM��!?d	����@#�rq�ٿ��f��@��7���3@MFM��!?d	����@#�rq�ٿ��f��@��7���3@MFM��!?d	����@��S�ٿ[V��u�@��,��3@����p�!?�-��Ɩ@��S�ٿ[V��u�@��,��3@����p�!?�-��Ɩ@X.�M�ٿ�����|�@���jT4@�v�s�!?�Bָݖ@D�M2�ٿ���y�@��>��3@b%�]�!?~c��gі@D�M2�ٿ���y�@��>��3@b%�]�!?~c��gі@+�֚͒ٿ,[��Mz�@�)]�54@B���+�!?o�	k�Ӗ@�#�ޛٿ��I2^�@@�{�3@QuK��!?l����v�@�#�ޛٿ��I2^�@@�{�3@QuK��!?l����v�@�#�ޛٿ��I2^�@@�{�3@QuK��!?l����v�@���ٿh���uw�@|c;��3@͆�JZ�!?��!t̖@�m�.הٿ���N�h�@�rEy�4@�Юt�!?ϟ����@�ѯ��ٿ�{�%zo�@��<��4@�2$d�!?T�$R���@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@��Ú��ٿC��\[�@qGI��3@��L���!?m��V�j�@�����ٿ�CX��[�@����4�3@VCCÐ!?�[�	n�@�����ٿ�CX��[�@����4�3@VCCÐ!?�[�	n�@�����ٿ�CX��[�@����4�3@VCCÐ!?�[�	n�@�����ٿ�CX��[�@����4�3@VCCÐ!?�[�	n�@�����ٿ�CX��[�@����4�3@VCCÐ!?�[�	n�@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@g���Țٿ�O�d�@�o��4@�z)a��!?)��`u��@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@�	��k�ٿ��TH�W�@}}{S�3@�z���!?sT5��_�@JO��ٿd"�D�@g�����3@�Z�z�!?���>�@JO��ٿd"�D�@g�����3@�Z�z�!?���>�@JO��ٿd"�D�@g�����3@�Z�z�!?���>�@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�{�WКٿB� �C�@!ܭ7d�3@�0�fj�!?n3E��@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@�؁Ζٿ0�	+9�@�9�!�#4@����̐!?��X���@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@nβ͛ٿ��S!�@�~}��3@�@��L�!?�U��Q��@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@#��mz�ٿ^��5i@�@�Wob�3@���N�!?D�e4�@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@}�~*�ٿ�x{�<�@���G/4@���l�!?]�f�V��@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@��:��ٿ� E�>�@����	4@8#�f�!?�F	D	�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@ X���ٿ��ę�C�@\B{$4@�i8�~�!?�kŵ�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@�a6�ٿ�%��D�@�����4@��̙�!?E�[�@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@���ٿ��f�T;�@ߥG���3@@��R��!?[�����@��X蕢ٿ�_���8�@ʂ�3y�3@�M�Vi�!?�D����@��X蕢ٿ�_���8�@ʂ�3y�3@�M�Vi�!?�D����@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@���'�ٿ<��@4�@�2�]��3@7�~��!?���ݤ�@]pc���ٿa� 1�V�@��~,�3@��L�e�!?��']�@]pc���ٿa� 1�V�@��~,�3@��L�e�!?��']�@]pc���ٿa� 1�V�@��~,�3@��L�e�!?��']�@]pc���ٿa� 1�V�@��~,�3@��L�e�!?��']�@��J}�ٿ%�s�NT�@�^�Nv"4@om�'@�!?'p�]R�@��J}�ٿ%�s�NT�@�^�Nv"4@om�'@�!?'p�]R�@[�8q^�ٿ܏��IW�@g���D/4@�|6E�!?��s^\�@[�8q^�ٿ܏��IW�@g���D/4@�|6E�!?��s^\�@`�j�ٿg���O�@�K�(�-4@ޖUz�!?:�[�B�@;L�Ėٿ��t�(�@w�b�M4@���*B�!?��?s��@;L�Ėٿ��t�(�@w�b�M4@���*B�!?��?s��@���ٿ(|L��S�@���'&4@�kԤ?�!?���JoP�@���ٿ(|L��S�@���'&4@�kԤ?�!?���JoP�@�=1�ٿ����F�@�-�:�Z4@<_�X�!?�-2�"�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@
 ~0�ٿzm3�P�@��i�74@��ᄐ!?���}E�@]�aϙٿԜVhY%�@H��4@	�C��!?�;��M��@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@���c^�ٿ���D�@��� 4@X�54��!?4zw�@4���Q�ٿĂ�&K=�@j�(A4@�e1Ň�!?$�����@4���Q�ٿĂ�&K=�@j�(A4@�e1Ň�!?$�����@4���Q�ٿĂ�&K=�@j�(A4@�e1Ň�!?$�����@4���Q�ٿĂ�&K=�@j�(A4@�e1Ň�!?$�����@4���Q�ٿĂ�&K=�@j�(A4@�e1Ň�!?$�����@���ٿ2�� +�@i��[=@4@mA��Y�!?�%"M�ĕ@���ٿ2�� +�@i��[=@4@mA��Y�!?�%"M�ĕ@���ٿ2�� +�@i��[=@4@mA��Y�!?�%"M�ĕ@+?@�ٿB���1�@��s��3@ܙ(1�!?}�[�ܕ@}Gswĝٿf�p�I�@��J.��3@�a�n�!?��$,1�@}Gswĝٿf�p�I�@��J.��3@�a�n�!?��$,1�@}Gswĝٿf�p�I�@��J.��3@�a�n�!?��$,1�@}Gswĝٿf�p�I�@��J.��3@�a�n�!?��$,1�@�z-�ٿ�uA�4>�@�h�h4@�.'�!?�x�d�@�z-�ٿ�uA�4>�@�h�h4@�.'�!?�x�d�@�z-�ٿ�uA�4>�@�h�h4@�.'�!?�x�d�@�z-�ٿ�uA�4>�@�h�h4@�.'�!?�x�d�@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@}�R��ٿCN���:�@7x���3@�(�M��!?i�,A��@!vAРٿ*�A�c�@8��7�O4@x5����!?YLϥ��@!vAРٿ*�A�c�@8��7�O4@x5����!?YLϥ��@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@5I���ٿ��|r�\�@�g/%8;4@�Yxb��!?K	�8n�@H#�!�ٿS�b�@���7B"4@e�rn�!?�������@H#�!�ٿS�b�@���7B"4@e�rn�!?�������@H#�!�ٿS�b�@���7B"4@e�rn�!?�������@H#�!�ٿS�b�@���7B"4@e�rn�!?�������@H#�!�ٿS�b�@���7B"4@e�rn�!?�������@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@D��{�ٿ��[MH[�@���W�4@���tz�!?�����i�@�wΕٿ��@!^�@ԡ3���3@X�Y�!?p�eљu�@�wΕٿ��@!^�@ԡ3���3@X�Y�!?p�eљu�@�wΕٿ��@!^�@ԡ3���3@X�Y�!?p�eљu�@�wΕٿ��@!^�@ԡ3���3@X�Y�!?p�eљu�@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@n�݃��ٿǄ�e�0�@���
4@b�Q��!?���~ڕ@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@U�5��ٿ�8�_�@)L	ŗ4@V�P��!?�H�m|z�@S*��h�ٿۆ��r-�@��L*�3@,&D�s�!?�{XRRϕ@�2pi�ٿ� �E�@�AI4��3@.�?7�!?3T;L)"�@�2pi�ٿ� �E�@�AI4��3@.�?7�!?3T;L)"�@�2pi�ٿ� �E�@�AI4��3@.�?7�!?3T;L)"�@��b�ٿo�Xr.�@P��2�3@ ����!?��Τ�ӕ@��b�ٿo�Xr.�@P��2�3@ ����!?��Τ�ӕ@��b�ٿo�Xr.�@P��2�3@ ����!?��Τ�ӕ@��b�ٿo�Xr.�@P��2�3@ ����!?��Τ�ӕ@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@�GFxV�ٿC�8��@�9芕�3@���}�!?eӲ̙b�@��ړd�ٿ$���:�@e�l]��3@�+�a{�!?ӼN�P��@��ړd�ٿ$���:�@e�l]��3@�+�a{�!?ӼN�P��@��ړd�ٿ$���:�@e�l]��3@�+�a{�!?ӼN�P��@��ړd�ٿ$���:�@e�l]��3@�+�a{�!?ӼN�P��@��ړd�ٿ$���:�@e�l]��3@�+�a{�!?ӼN�P��@>�T\��ٿ2%7-�@����L4@�a�{�!?ë�v�˕@>�T\��ٿ2%7-�@����L4@�a�{�!?ë�v�˕@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@�	��!�ٿ�%=�J?�@"����3@i=�d�!?O�Hkl�@bN�w0�ٿł)��+�@mLV���3@��,�H�!?�F�ʕ@bN�w0�ٿł)��+�@mLV���3@��,�H�!?�F�ʕ@p���ٿ�����D�@+����4@d�i�!?�5�n��@p���ٿ�����D�@+����4@d�i�!?�5�n��@p���ٿ�����D�@+����4@d�i�!?�5�n��@�O��N�ٿ���/�D�@8l}�N04@#w����!?��B��@�O��N�ٿ���/�D�@8l}�N04@#w����!?��B��@�O��N�ٿ���/�D�@8l}�N04@#w����!?��B��@�O��N�ٿ���/�D�@8l}�N04@#w����!?��B��@�O��N�ٿ���/�D�@8l}�N04@#w����!?��B��@f|闚ٿ:�����@��}DL4@!����!?�l3lf��@f|闚ٿ:�����@��}DL4@!����!?�l3lf��@f|闚ٿ:�����@��}DL4@!����!?�l3lf��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@`��Y�ٿ%���@&I��.�3@�����!?��Rm��@uuN_�ٿ���D�R�@tIˤ=54@��!�Ӑ!?}��TK�@uuN_�ٿ���D�R�@tIˤ=54@��!�Ӑ!?}��TK�@ 
}�"�ٿ���2�@���3@�"E��!?.Ϊ�ޕ@ 
}�"�ٿ���2�@���3@�"E��!?.Ϊ�ޕ@ 
}�"�ٿ���2�@���3@�"E��!?.Ϊ�ޕ@ 
}�"�ٿ���2�@���3@�"E��!?.Ϊ�ޕ@ 
}�"�ٿ���2�@���3@�"E��!?.Ϊ�ޕ@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@���;�ٿ�LV<�6�@�;�hP�3@��-�W�!?o�����@�R�q��ٿ�v6��6�@?k����3@y�"�]�!?�ψ��@�R�q��ٿ�v6��6�@?k����3@y�"�]�!?�ψ��@�R�q��ٿ�v6��6�@?k����3@y�"�]�!?�ψ��@���J1�ٿOAcymD�@�K�;}�3@�`��!?�1%��@io�
�ٿ<���q=�@*����E4@��K���!?`ͽ� �@io�
�ٿ<���q=�@*����E4@��K���!?`ͽ� �@io�
�ٿ<���q=�@*����E4@��K���!?`ͽ� �@io�
�ٿ<���q=�@*����E4@��K���!?`ͽ� �@io�
�ٿ<���q=�@*����E4@��K���!?`ͽ� �@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@L�X>��ٿ&���2+�@�9��Y�3@)}?�:�!?cn�]Ǖ@P�����ٿ��'A�@G�?��3@��P�!?�\uG��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@54~7Ӟٿ��Hn�5�@�p�{� 4@�{Ɛ!?�b\��@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��]&|�ٿL���F�@H3R	��3@_�W預!?b�P$�@��r6�ٿ }"G8�@�����3@�nY�z�!?� d!l��@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@���6��ٿ��x��,�@A`?�m�3@�G��W�!?M��_ ͕@��ا�ٿ�� +A�@D���3@�ң�v�!?���E��@��ا�ٿ�� +A�@D���3@�ң�v�!?���E��@��g)�ٿ�Ɨ�S=�@�l����3@$���;�!?��Ye��@��g)�ٿ�Ɨ�S=�@�l����3@$���;�!?��Ye��@��g)�ٿ�Ɨ�S=�@�l����3@$���;�!?��Ye��@�2��ٿQ6���;�@�>?>��3@��6z�!?��
���@�2��ٿQ6���;�@�>?>��3@��6z�!?��
���@�2��ٿQ6���;�@�>?>��3@��6z�!?��
���@�2��ٿQ6���;�@�>?>��3@��6z�!?��
���@ȇ�.��ٿ-����@��/��3@|��YO�!?����x�@b@Yl�ٿY�-��2�@��˃��3@3��!?�
�x��@b@Yl�ٿY�-��2�@��˃��3@3��!?�
�x��@b@Yl�ٿY�-��2�@��˃��3@3��!?�
�x��@b@Yl�ٿY�-��2�@��˃��3@3��!?�
�x��@�jR�ٿ�c�_�:�@�└/4@�㲂S�!?��i�d��@��{q��ٿft�H�J�@p����3@�9l�!?ќ�2�@��)��ٿ5{��4�@
�^��3@�p��!?�N��Y�@O����ٿOu���:�@��Vf64@��~!�!?�6����@O����ٿOu���:�@��Vf64@��~!�!?�6����@O����ٿOu���:�@��Vf64@��~!�!?�6����@?� `n�ٿ��D���@{/*��4@xJ���!?���g��@?� `n�ٿ��D���@{/*��4@xJ���!?���g��@���:�ٿ�;i�/�@�"j�`4@���2�!?�^$MzЕ@�V8�v�ٿ䑈%#9�@0h}|G4@�|�U&�!?�D�@�V8�v�ٿ䑈%#9�@0h}|G4@�|�U&�!?�D�@�V8�v�ٿ䑈%#9�@0h}|G4@�|�U&�!?�D�@�V8�v�ٿ䑈%#9�@0h}|G4@�|�U&�!?�D�@�D�!�ٿy%,V+�@u&~�=U4@�i��8�!?����^@�D�!�ٿy%,V+�@u&~�=U4@�i��8�!?����^@#�0ؖ�ٿ�re��@,� ��24@`s=���!?��ºk�@;�3��ٿ�C2��@��s��3@27}KԐ!?��O䚕@;�3��ٿ�C2��@��s��3@27}KԐ!?��O䚕@ʷ��ٿy)��C�@�W@�3@!6D�!?���A��@ʷ��ٿy)��C�@�W@�3@!6D�!?���A��@ʷ��ٿy)��C�@�W@�3@!6D�!?���A��@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@���?�ٿ�I1��>�@�9[���3@���yI�!?���f%�@��'��ٿu���O�@8p����3@�I*k�!?R ���C�@n_�d�ٿ��`�D�@2!����3@�_�˦�!?5Z��e!�@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@�3�5�ٿ:���t�@)�2sH4@$%��!?�N�*���@x�r���ٿ6�O*9�@��M[�3@_�����!?Џ�ӑ��@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@�q4��ٿ�bS�"�@@/�)b�3@����i�!?wv��ʨ�@6*�:A�ٿ��hQ,3�@\��Z$.4@A�+/�!?�
ޖ��@6*�:A�ٿ��hQ,3�@\��Z$.4@A�+/�!?�
ޖ��@6*�:A�ٿ��hQ,3�@\��Z$.4@A�+/�!?�
ޖ��@Ϛ�Q�ٿ#R��LC�@�P ^�F4@��+�!?��}��@Ϛ�Q�ٿ#R��LC�@�P ^�F4@��+�!?��}��@Ϛ�Q�ٿ#R��LC�@�P ^�F4@��+�!?��}��@Ϛ�Q�ٿ#R��LC�@�P ^�F4@��+�!?��}��@����٣ٿ���p\�@�fm��"4@��$�!?}OA�m�@����٣ٿ���p\�@�fm��"4@��$�!?}OA�m�@����٣ٿ���p\�@�fm��"4@��$�!?}OA�m�@�Z/�ٿ���kP�@��͸3K4@����!?y���{B�@�Z/�ٿ���kP�@��͸3K4@����!?y���{B�@�Z/�ٿ���kP�@��͸3K4@����!?y���{B�@�Z/�ٿ���kP�@��͸3K4@����!?y���{B�@�Z/�ٿ���kP�@��͸3K4@����!?y���{B�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@�#����ٿHd�UN�@0[�4@Hg�'�!?.2o?�@_.����ٿ��siHC�@�7���3@�v�AN�!?��$@�@_.����ٿ��siHC�@�7���3@�v�AN�!?��$@�@!g��u�ٿJ����&�@q}>��3@�$j`�!?.�W1}��@!g��u�ٿJ����&�@q}>��3@�$j`�!?.�W1}��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@����ٿyX� %�@}N���3@p�kb�!?18��@v�%�ٿ�5G�[8�@��ؓB4@��ת��!?f��K��@v�%�ٿ�5G�[8�@��ؓB4@��ת��!?f��K��@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@�}���ٿ��|=�@|l�}4@�EyM��!?jo���@HT�ٿ�M�b�9�@ S��44@�s����!?N�����@HT�ٿ�M�b�9�@ S��44@�s����!?N�����@���Z3�ٿ�Bۨ�,�@����G4@���ԙ�!?.L�7�Ǖ@���Z3�ٿ�Bۨ�,�@����G4@���ԙ�!?.L�7�Ǖ@�G�8	�ٿh퓲�1�@b�P&4@��$Kn�!?��E�ܕ@�G�8	�ٿh퓲�1�@b�P&4@��$Kn�!?��E�ܕ@%�ӡٿö��W�@��#�)4@�Y%X1�!?C<L�za�@I�'{A�ٿ�B��V�@^���4@�.�!?�_1��^�@I�'{A�ٿ�B��V�@^���4@�.�!?�_1��^�@�6��ٿ����F�@[.��J4@�o��:�!?3λat$�@�6��ٿ����F�@[.��J4@�o��:�!?3λat$�@:�C��ٿ�Sk��*�@;�K��4@�,�(a�!?��{7Ǖ@:�C��ٿ�Sk��*�@;�K��4@�,�(a�!?��{7Ǖ@(8�H(�ٿʸ7-�^�@M���;4@�5k,�!?}�70~�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@*ĵ�t�ٿ��قpO�@�=�-4@DeL,��!?]���J�@�<�nʚٿb<�P	�@�$���4@�N����!?���胕@�<�nʚٿb<�P	�@�$���4@�N����!?���胕@壘ٿw��1�@$v(�3@Pn��t�!?�p�$���@壘ٿw��1�@$v(�3@Pn��t�!?�p�$���@壘ٿw��1�@$v(�3@Pn��t�!?�p�$���@壘ٿw��1�@$v(�3@Pn��t�!?�p�$���@壘ٿw��1�@$v(�3@Pn��t�!?�p�$���@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@7����ٿd!�԰3�@�5��3@�²�!?�����@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@x�.�e�ٿ��*�=�@��
��4@d�����!?|gl��@�?`ҙ�ٿ��S��;�@����;4@�.5�!?V�����@�?`ҙ�ٿ��S��;�@����;4@�.5�!?V�����@�?`ҙ�ٿ��S��;�@����;4@�.5�!?V�����@�?`ҙ�ٿ��S��;�@����;4@�.5�!?V�����@��8[ܚٿ-�:�D<�@��G9%4@r#\m*�!?�e-\b�@0���ٿ�Z��@�@�P�Q}64@�!�?��!?}����@0���ٿ�Z��@�@�P�Q}64@�!�?��!?}����@0���ٿ�Z��@�@�P�Q}64@�!�?��!?}����@0���ٿ�Z��@�@�P�Q}64@�!�?��!?}����@�
�ٿ|#t�z*�@��}G&4@��xx�!?�w�q��@�
�ٿ|#t�z*�@��}G&4@��xx�!?�w�q��@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@s���ٿ]m���7�@D����3@6;�PO�!?n�Pp�@;V�7�ٿ����F4�@�O��
$4@ǰ���!?s�;��@;V�7�ٿ����F4�@�O��
$4@ǰ���!?s�;��@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@��+�c�ٿn�d��@�9w�4@���@*�!?���#���@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@Iy�,
�ٿ���1�@ܞ�/�4@�~M�!?�R�E��@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@prޚٿ�4L�
'�@Ɠ"*D.4@I�9&�!?����ɪ�@6�+s�ٿYU��"�@�����3@��j��!?�D�pI��@6�+s�ٿYU��"�@�����3@��j��!?�D�pI��@Y�o�z�ٿ�C�+.Z�@�yR��3@��q�c�!?�a�n j�@Y�o�z�ٿ�C�+.Z�@�yR��3@��q�c�!?�a�n j�@Y�o�z�ٿ�C�+.Z�@�yR��3@��q�c�!?�a�n j�@.;Y�ٿG��\+�@�Pɣ24@v�~lS�!?����@.;Y�ٿG��\+�@�Pɣ24@v�~lS�!?����@: `ri�ٿ?�b.�@���4@��!���!?~=Dh�ە@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�L2�\�ٿe��O�@n����3@n
�p�!?sd�W�U�@�LDWR�ٿ��b��)�@^�8��4@�e>��!?P�7�r��@�LDWR�ٿ��b��)�@^�8��4@�e>��!?P�7�r��@�LDWR�ٿ��b��)�@^�8��4@�e>��!?P�7�r��@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@�%$Q�ٿ���(�"�@��D���3@ Đ�!?W�=&���@1�$��ٿ�141=8�@�t]��3@�զ4'�!?�O"�t�@a���ٿ����^C�@A#���3@���E�!?<����@a���ٿ����^C�@A#���3@���E�!?<����@a���ٿ����^C�@A#���3@���E�!?<����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@U%;w�ٿ��<J1�@�3s�a*4@��u%a�!?�o����@@*ۘٿ��:K�-�@�])�n	4@F�qK�!?0�5��ҕ@@*ۘٿ��:K�-�@�])�n	4@F�qK�!?0�5��ҕ@@*ۘٿ��:K�-�@�])�n	4@F�qK�!?0�5��ҕ@����s�ٿ�g��&�@c�c��"4@�O`��!?�|�;��@����s�ٿ�g��&�@c�c��"4@�O`��!?�|�;��@����s�ٿ�g��&�@c�c��"4@�O`��!?�|�;��@,��lءٿPs'X.�@{̼W&4@J�-C�!?�@ۇ�ϕ@,��lءٿPs'X.�@{̼W&4@J�-C�!?�@ۇ�ϕ@,��lءٿPs'X.�@{̼W&4@J�-C�!?�@ۇ�ϕ@,��lءٿPs'X.�@{̼W&4@J�-C�!?�@ۇ�ϕ@b<����ٿ���/�@P���	4@E��0o�!?I���ܕ@b<����ٿ���/�@P���	4@E��0o�!?I���ܕ@�P#�ʞٿ�AL�P�@U2P��4@O��P�!?��P(P�@��E��ٿ���O6�@\@z1� 4@�ms�>�!?>������@��E��ٿ���O6�@\@z1� 4@�ms�>�!?>������@��E��ٿ���O6�@\@z1� 4@�ms�>�!?>������@Æ��T�ٿ18ݖ2�@����3@�~��S�!?�����@Æ��T�ٿ18ݖ2�@����3@�~��S�!?�����@Æ��T�ٿ18ݖ2�@����3@�~��S�!?�����@Æ��T�ٿ18ݖ2�@����3@�~��S�!?�����@�}��N�ٿJd L�D�@o;��8�3@M��▐!?�X=��!�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@W���[�ٿ��2?�@1�֟4@%w����!?���b�@ES��ٿ�8<��j�@���N4@�Q�r�!?�H{ԡ��@ԕ�/2�ٿ=)��gn�@>#[,@4@"�Ð!?�Q�O�Ė@ԕ�/2�ٿ=)��gn�@>#[,@4@"�Ð!?�Q�O�Ė@�sB�ٿTC��V�@� yx�E4@��뷌�!?�U��d�@�sB�ٿTC��V�@� yx�E4@��뷌�!?�U��d�@�sB�ٿTC��V�@� yx�E4@��뷌�!?�U��d�@�sB�ٿTC��V�@� yx�E4@��뷌�!?�U��d�@�sB�ٿTC��V�@� yx�E4@��뷌�!?�U��d�@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@d����ٿ2�f�rI�@F˷�~S4@]�i�z�!?�A` �@�h� ��ٿ��Ii]�@�s��44@׷	Q�!?3�,m�o�@�h� ��ٿ��Ii]�@�s��44@׷	Q�!?3�,m�o�@n�����ٿ��G FN�@��I�4@��tU��!?�Ld@A�@upG��ٿ�d65m#�@^D����3@ą�ɋ�!?U1���@upG��ٿ�d65m#�@^D����3@ą�ɋ�!?U1���@� �ٿ2J��r��@#�'g�3@h���M�!?,�S;�@� �ٿ2J��r��@#�'g�3@h���M�!?,�S;�@� �ٿ2J��r��@#�'g�3@h���M�!?,�S;�@M�WeG�ٿ����@V!q���3@��q�ڏ!?����fh�@M�WeG�ٿ����@V!q���3@��q�ڏ!?����fh�@*�Y�ŦٿVqP�za�@�*���3@|����!?}�����@�Z�6}�ٿ$R '��@|�7X��3@�{�VG�!?O�#r��@�Z�6}�ٿ$R '��@|�7X��3@�{�VG�!?O�#r��@�Z�6}�ٿ$R '��@|�7X��3@�{�VG�!?O�#r��@#m,6/�ٿ,�eu�^�@�U^�`4@ �>�~�!?�tЭ�[�@#m,6/�ٿ,�eu�^�@�U^�`4@ �>�~�!?�tЭ�[�@#m,6/�ٿ,�eu�^�@�U^�`4@ �>�~�!?�tЭ�[�@#m,6/�ٿ,�eu�^�@�U^�`4@ �>�~�!?�tЭ�[�@���#�ٿ-��pH`�@�
Xl�+4@#`B0�!?��3uZu�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@��x��ٿ{E�k�K�@P����:4@��M��!?���"9:�@���ٿ80��A�@fGpf�3@�B��!?��'�$�@���ٿ80��A�@fGpf�3@�B��!?��'�$�@���ٿ80��A�@fGpf�3@�B��!?��'�$�@���ٿ80��A�@fGpf�3@�B��!?��'�$�@�Mվ��ٿ^G�85�@��L�3@�Է��!?�j�w$�@�Mվ��ٿ^G�85�@��L�3@�Է��!?�j�w$�@�qH4�ٿX��B`�@��ߊ7�3@T�Wȥ�!?�jUҜ��@�qH4�ٿX��B`�@��ߊ7�3@T�Wȥ�!?�jUҜ��@�qH4�ٿX��B`�@��ߊ7�3@T�Wȥ�!?�jUҜ��@�qH4�ٿX��B`�@��ߊ7�3@T�Wȥ�!?�jUҜ��@�qH4�ٿX��B`�@��ߊ7�3@T�Wȥ�!?�jUҜ��@F�$��ٿqۜAq@�@^x6UU�3@(IJ���!?@t^�1/�@F�$��ٿqۜAq@�@^x6UU�3@(IJ���!?@t^�1/�@F�$��ٿqۜAq@�@^x6UU�3@(IJ���!?@t^�1/�@F�$��ٿqۜAq@�@^x6UU�3@(IJ���!?@t^�1/�@@�7�ٿ ���@'�@�h�3@�g�T�!?z���.��@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@fu¥ٿ|���]>�@.�]r4@�d�䍐!?Ҳ�K+�@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@�9v댢ٿ$}P�8�@�2�H4@oJ����!?�f,ͯڕ@p���s�ٿ�H�F�=�@'J�Lv64@���wg�!?kk��=�@p���s�ٿ�H�F�=�@'J�Lv64@���wg�!?kk��=�@p���s�ٿ�H�F�=�@'J�Lv64@���wg�!?kk��=�@���8�ٿz4*׵N�@@m��uQ4@3��f"�!?�'�CB�@���8�ٿz4*׵N�@@m��uQ4@3��f"�!?�'�CB�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@>�N]��ٿ���`%T�@W��@��3@y��{�!?:�DFh`�@�Ϯ ��ٿP�/SO�@j3$�3@�#�K<�!?h���V]�@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@Ʒj-�ٿ2��5ZX�@7��D�3@�Jl<J�!?�p����@����H�ٿ�-�`�9�@K.��74@I��̸�!?,ɕo��@����H�ٿ�-�`�9�@K.��74@I��̸�!?,ɕo��@����H�ٿ�-�`�9�@K.��74@I��̸�!?,ɕo��@Y�͸Кٿ�|]�2�@�:�14@V�5p�!?���Oϕ@Y�͸Кٿ�|]�2�@�:�14@V�5p�!?���Oϕ@Y�͸Кٿ�|]�2�@�:�14@V�5p�!?���Oϕ@Y�͸Кٿ�|]�2�@�:�14@V�5p�!?���Oϕ@Q�! �ٿ�K-ڎY�@+!�F�-4@�Ptc=�!?�e�$zH�@Q�! �ٿ�K-ڎY�@+!�F�-4@�Ptc=�!?�e�$zH�@Q�! �ٿ�K-ڎY�@+!�F�-4@�Ptc=�!?�e�$zH�@Q�! �ٿ�K-ڎY�@+!�F�-4@�Ptc=�!?�e�$zH�@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@�쵱�ٿS��b�@�(���3@f\ޛ@�!?f��@����J�ٿ�[�O�@p#�m�4@��f���!?ö8�A�@����J�ٿ�[�O�@p#�m�4@��f���!?ö8�A�@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@=&3bʠٿ��bkA�@<SFr+�3@��{MM�!?��y��@{�؛ٿ/d��K>�@���V�3@oeN^�!?�➭�@{�؛ٿ/d��K>�@���V�3@oeN^�!?�➭�@W;�Ӵ�ٿֆ�%M/�@�����	4@(j���!?�`����@W;�Ӵ�ٿֆ�%M/�@�����	4@(j���!?�`����@W;�Ӵ�ٿֆ�%M/�@�����	4@(j���!?�`����@W;�Ӵ�ٿֆ�%M/�@�����	4@(j���!?�`����@W;�Ӵ�ٿֆ�%M/�@�����	4@(j���!?�`����@p���8�ٿy��Ǉ<�@�_JS4@�;E,�!?S��̼�@p���8�ٿy��Ǉ<�@�_JS4@�;E,�!?S��̼�@p���8�ٿy��Ǉ<�@�_JS4@�;E,�!?S��̼�@p���8�ٿy��Ǉ<�@�_JS4@�;E,�!?S��̼�@p���8�ٿy��Ǉ<�@�_JS4@�;E,�!?S��̼�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@ r���ٿ�'�m!�@��T%s4@JA����!?�4��ɖ�@EcQEO�ٿ���21$�@��V84@���A��!?�D�O�@��g$�ٿ��v��@Ȯ��A4@7��%c�!?�<�Icr�@@�EE?�ٿ:��g82�@��,�X4@ڄ����!?�bLtؕ@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@R���:�ٿ��r5�@��� 6�3@��y���!?��t���@X%뇙�ٿ8�V��\�@=��}4�3@z�:�!?����^�@X%뇙�ٿ8�V��\�@=��}4�3@z�:�!?����^�@��gߞٿ�w[G�@fCB�(D4@��Y�!?A�&p�@��gߞٿ�w[G�@fCB�(D4@��Y�!?A�&p�@�Y�bޡٿ�1ڬC�@�;�4@�s���!?
�U�&�@�Y�bޡٿ�1ڬC�@�;�4@�s���!?
�U�&�@�Y�bޡٿ�1ڬC�@�;�4@�s���!?
�U�&�@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@�M��ٿ�y���<�@}h��@�3@���V�!?S���@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@��I�ٿ�ٽ�-�@�G�&%�3@�$�#�!?o
=�r��@�{İ;�ٿ����OF�@��*�h4@��UO�!?I�~�a�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@��gc1�ٿ;�-�b[�@(O�fh	4@z�2�\�!?�m�Tqg�@����̗ٿ�h�GK�@u�p�3@��b�!?�]�kw)�@m>%Œ�ٿ��N�E�@���EC4@�a~CG�!?�d^e���@m>%Œ�ٿ��N�E�@���EC4@�a~CG�!?�d^e���@m>%Œ�ٿ��N�E�@���EC4@�a~CG�!?�d^e���@m>%Œ�ٿ��N�E�@���EC4@�a~CG�!?�d^e���@����.�ٿ�s�"�@?�NQ�4@�>5�_�!?27C�P��@�3�V3�ٿ'BR �C�@��N��3@�G�)�!?FLt��@�3�V3�ٿ'BR �C�@��N��3@�G�)�!?FLt��@��T	�ٿ�[#4�@�B���3@7],�y�!?��mxS�@��T	�ٿ�[#4�@�B���3@7],�y�!?��mxS�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@�$���ٿ%X��>U�@�V?&�4@\�ӗ:�!?�4�^�@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@��ê*�ٿ?�Y��4�@�`�xe�3@�f�A�!?�j!�ޕ@Ũ�b/�ٿ��D�E�@Y���4@cV�'X�!?3;���'�@Ũ�b/�ٿ��D�E�@Y���4@cV�'X�!?3;���'�@Ũ�b/�ٿ��D�E�@Y���4@cV�'X�!?3;���'�@T�݆]�ٿ���V_�@.'���4@�b��;�!?țH�r�@T�݆]�ٿ���V_�@.'���4@�b��;�!?țH�r�@T�݆]�ٿ���V_�@.'���4@�b��;�!?țH�r�@����ٿ6��/�B�@�#v4@�}��!?��^*�@����ٿ6��/�B�@�#v4@�}��!?��^*�@�g��ٿת��4>�@
-�[~�3@�}
K�!?M|K_]��@�~��T�ٿQ����B�@��4@��O���!?�@`ڕ@�~��T�ٿQ����B�@��4@��O���!?�@`ڕ@�~��T�ٿQ����B�@��4@��O���!?�@`ڕ@�~��T�ٿQ����B�@��4@��O���!?�@`ڕ@�~��T�ٿQ����B�@��4@��O���!?�@`ڕ@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@Yw�R�ٿ����@��C8;�3@S��X#�!?ѹ/�?H�@������ٿq5�tNC�@��3��3@6�癆�!?x�{��'�@������ٿq5�tNC�@��3��3@6�癆�!?x�{��'�@9o��T�ٿ�x?C�<�@3��3@��]���!?3���M�@9o��T�ٿ�x?C�<�@3��3@��]���!?3���M�@9o��T�ٿ�x?C�<�@3��3@��]���!?3���M�@���.4�ٿ�vA5�C�@кi�54@�)�*ܐ!?�a]lM�@Nr,�ٿ���m;�@xxf�!4@�V
�s�!?U1�:�&�@Nr,�ٿ���m;�@xxf�!4@�V
�s�!?U1�:�&�@Nr,�ٿ���m;�@xxf�!4@�V
�s�!?U1�:�&�@h[�d��ٿp�'sL�@v�G 4@��Gz�!?Z�[мT�@h[�d��ٿp�'sL�@v�G 4@��Gz�!?Z�[мT�@݇�ؠٿA{�BK�@!h#4@�!`�r�!?����Mb�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@N��ɢٿh�� ]=�@��ѐ�#4@�ጉ�!?xB�!o=�@�xjW�ٿ�^�{�:�@���}K%4@�;���!?���d��@�xjW�ٿ�^�{�:�@���}K%4@�;���!?���d��@�xjW�ٿ�^�{�:�@���}K%4@�;���!?���d��@�	���ٿ;�q�h�@X{B�4@��d��!?��e4&��@�	���ٿ;�q�h�@X{B�4@��d��!?��e4&��@�	���ٿ;�q�h�@X{B�4@��d��!?��e4&��@�	���ٿ;�q�h�@X{B�4@��d��!?��e4&��@�	���ٿ;�q�h�@X{B�4@��d��!?��e4&��@\o'YҚٿ��� A[�@:$��
4@�k9�!?�J�j��@\o'YҚٿ��� A[�@:$��
4@�k9�!?�J�j��@��*s�ٿ�@�!B�@ِ��4@zG��G�!?R��L�@��*s�ٿ�@�!B�@ِ��4@zG��G�!?R��L�@��*s�ٿ�@�!B�@ِ��4@zG��G�!?R��L�@��*s�ٿ�@�!B�@ِ��4@zG��G�!?R��L�@;����ٿQ�S�^A�@�ӑ�4@����!?���D�M�@;����ٿQ�S�^A�@�ӑ�4@����!?���D�M�@;����ٿQ�S�^A�@�ӑ�4@����!?���D�M�@eA�7�ٿmKc@�/�@`�L���3@��v�!?b�S��@eA�7�ٿmKc@�/�@`�L���3@��v�!?b�S��@�!����ٿg��\�8�@��� 24@�p(L\�!?%)j�sM�@�!����ٿg��\�8�@��� 24@�p(L\�!?%)j�sM�@�!����ٿg��\�8�@��� 24@�p(L\�!?%)j�sM�@�!����ٿg��\�8�@��� 24@�p(L\�!?%)j�sM�@�!����ٿg��\�8�@��� 24@�p(L\�!?%)j�sM�@FAF�l�ٿ�����@���>�4@o]�#��!?:������@FAF�l�ٿ�����@���>�4@o]�#��!?:������@FAF�l�ٿ�����@���>�4@o]�#��!?:������@FAF�l�ٿ�����@���>�4@o]�#��!?:������@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@Zv�9!�ٿ��!�q��@�TQ���3@�G�Zn�!?؞�4�0�@W��ٿw�?J��@5��ǣ�3@�r�"1�!?=g�[ڕ@��@��ٿ7W˘��@"�,�e4@᪞[��!?��؈��@؂��,�ٿiKF��
�@�}�%4@��37�!?�e�[フ@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@և����ٿf^Ov�e�@�%du=4@fca&��!?,I��F�@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@Nz���ٿ��d&�@�ȳ�u�3@���+$�!?%cV˕@p �i�ٿ��"�bJ�@8���<�3@�j�Q�!?ĖXq@��@p �i�ٿ��"�bJ�@8���<�3@�j�Q�!?ĖXq@��@p �i�ٿ��"�bJ�@8���<�3@�j�Q�!?ĖXq@��@p �i�ٿ��"�bJ�@8���<�3@�j�Q�!?ĖXq@��@p �i�ٿ��"�bJ�@8���<�3@�j�Q�!?ĖXq@��@��Y!�ٿ�%��5�@��鬹�3@������!?�0;+_R�@��Y!�ٿ�%��5�@��鬹�3@������!?�0;+_R�@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@�9V�ٿ���l�@�~�'�3@2Ȋ[�!?�M��攕@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@8G�՞ٿ��D#u�@�oJ:��3@�*G�!?#���O�@n�0 *�ٿ�K	�h�@.5�Q��3@u{�>t�!?z���+�@n�0 *�ٿ�K	�h�@.5�Q��3@u{�>t�!?z���+�@n�0 *�ٿ�K	�h�@.5�Q��3@u{�>t�!?z���+�@zO1�ݛٿ'�;N8�@Y��3@lOߏ!?rӵ.&ѕ@��z)�ٿu�zB�@B5��,�3@7��!�!?5�`���@at���ٿ��>�@�=���4@�Z�!?r5�NWz�@��*�]�ٿ����2�@�V�4@�K6��!?A�Uw%�@��*�]�ٿ����2�@�V�4@�K6��!?A�Uw%�@��*�]�ٿ����2�@�V�4@�K6��!?A�Uw%�@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�7$�ٿ����R�@��S3H4@�RW��!?�b��֕@�{�>��ٿ*Pe2�B�@� +���3@��µw�!?�_s���@�{�>��ٿ*Pe2�B�@� +���3@��µw�!?�_s���@�{�>��ٿ*Pe2�B�@� +���3@��µw�!?�_s���@�{�>��ٿ*Pe2�B�@� +���3@��µw�!?�_s���@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@����ٿ�>��Vi�@��I��3@�z�}�!?mǉՕ@�=ݝ�ٿ/��2���@k��3@U1��!?���N��@�=ݝ�ٿ/��2���@k��3@U1��!?���N��@�=ݝ�ٿ/��2���@k��3@U1��!?���N��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@�,���ٿ�1�e��@9*�r[4@&��g�!?/�d��@����ٿ�P���r�@|�i��+4@Y�oS�!?�:;2��@����ٿ�P���r�@|�i��+4@Y�oS�!?�:;2��@����ٿ�P���r�@|�i��+4@Y�oS�!?�:;2��@����ٿ�P���r�@|�i��+4@Y�oS�!?�:;2��@��g �ٿg�ٿ��@��;Y@24@��Y��!?{|��S�@��g �ٿg�ٿ��@��;Y@24@��Y��!?{|��S�@��g �ٿg�ٿ��@��;Y@24@��Y��!?{|��S�@��g �ٿg�ٿ��@��;Y@24@��Y��!?{|��S�@��g �ٿg�ٿ��@��;Y@24@��Y��!?{|��S�@��`I��ٿ�oa���@��.�c 4@�M�*�!?F�uQY�@���"7�ٿ���
��@���4@�<�4ܐ!??]>q`r�@���"7�ٿ���
��@���4@�<�4ܐ!??]>q`r�@���"7�ٿ���
��@���4@�<�4ܐ!??]>q`r�@���"7�ٿ���
��@���4@�<�4ܐ!??]>q`r�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@�Hw�J�ٿ��a���@y�LF�>4@�B�L�!?2T��x�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@h�۠ٿq���Q��@٢W��54@L,�Sb�!?����_D�@N'�ٿ �蘖�@�D��!�3@�vdŜ�!?E�?�MT�@�����ٿ�v�x���@�JR���3@�p���!?�ԫ����@�����ٿ�v�x���@�JR���3@�p���!?�ԫ����@)7F:��ٿ�;OZ%~�@��5�(4@m�y���!?��1jؕ@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@<0(�ٿ�Zp�W�@�ѫ"4@�;�ܕ�!?
t�r��@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@��Xn�ٿ<�����@q*bUY04@��i��!?���q���@s���y�ٿ�=ZMu�@4q)�64@W���z�!?��-�Õ@s���y�ٿ�=ZMu�@4q)�64@W���z�!?��-�Õ@s���y�ٿ�=ZMu�@4q)�64@W���z�!?��-�Õ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@o
l�ٿ�4"��@����$4@F9vS,�!?���ꖕ@C}? �ٿ�'9Or��@a{F+B�3@@��L@�!?S{���g�@C}? �ٿ�'9Or��@a{F+B�3@@��L@�!?S{���g�@綶v�ٿ.]�p�#�@z)T�'�3@��Xh�!?5D�C�d�@綶v�ٿ.]�p�#�@z)T�'�3@��Xh�!?5D�C�d�@綶v�ٿ.]�p�#�@z)T�'�3@��Xh�!?5D�C�d�@綶v�ٿ.]�p�#�@z)T�'�3@��Xh�!?5D�C�d�@��
�N�ٿGR$��@��54@;�9Q�!?��Ⱦ��@��
�N�ٿGR$��@��54@;�9Q�!?��Ⱦ��@��
�N�ٿGR$��@��54@;�9Q�!?��Ⱦ��@��
�N�ٿGR$��@��54@;�9Q�!?��Ⱦ��@h�5��ٿ��E�v�@�u� 4@5�-��!?������@h�5��ٿ��E�v�@�u� 4@5�-��!?������@h�5��ٿ��E�v�@�u� 4@5�-��!?������@h�5��ٿ��E�v�@�u� 4@5�-��!?������@h�5��ٿ��E�v�@�u� 4@5�-��!?������@J�h[��ٿh��fxU�@J�ܛ4@�@U��!?F�?�ev�@J�h[��ٿh��fxU�@J�ܛ4@�@U��!?F�?�ev�@�Nތ��ٿ� o�D�@K�|.ju4@��B�!?/��ߑ�@�Nތ��ٿ� o�D�@K�|.ju4@��B�!?/��ߑ�@�Nތ��ٿ� o�D�@K�|.ju4@��B�!?/��ߑ�@�Nތ��ٿ� o�D�@K�|.ju4@��B�!?/��ߑ�@�Nތ��ٿ� o�D�@K�|.ju4@��B�!?/��ߑ�@�ʉդٿh㈾���@^ս��;4@�S}#��!?N}����@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�����ٿ ���@���4@@�s�J�!?�������@�g3�ٿ)َ�]��@d���3@(�/bG�!?~<�Э!�@�g3�ٿ)َ�]��@d���3@(�/bG�!?~<�Э!�@�g3�ٿ)َ�]��@d���3@(�/bG�!?~<�Э!�@�g3�ٿ)َ�]��@d���3@(�/bG�!?~<�Э!�@S���ٿ&�x%G�@��%Z4@~��Rr�!?�{����@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@"��2�ٿ�?7�@e�-Xg�3@�g���!?M�V�#R�@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@��O�ٿڡilu��@�)Mb��3@kC,���!?8�����@~2l�؟ٿdF�w���@��{���3@��U�!?1�����@��MqZ�ٿ�4����@�����3@x�/�!?_+Z����@��MqZ�ٿ�4����@�����3@x�/�!?_+Z����@��MqZ�ٿ�4����@�����3@x�/�!?_+Z����@��MqZ�ٿ�4����@�����3@x�/�!?_+Z����@|U�-��ٿ��oA���@n�=� 94@�f���!?��M1N�@|U�-��ٿ��oA���@n�=� 94@�f���!?��M1N�@|U�-��ٿ��oA���@n�=� 94@�f���!?��M1N�@|U�-��ٿ��oA���@n�=� 94@�f���!?��M1N�@|U�-��ٿ��oA���@n�=� 94@�f���!?��M1N�@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@�ҕ��ٿ�6	��X�@��N��H4@ҫ@�v�!?*�����@���7�ٿ �.�;��@C�}�4@8Ts�M�!?V�I�̞�@���7�ٿ �.�;��@C�}�4@8Ts�M�!?V�I�̞�@���7�ٿ �.�;��@C�}�4@8Ts�M�!?V�I�̞�@Ǵʌ%�ٿQa*E�@���:�3@-lF���!?+͆s���@Ǵʌ%�ٿQa*E�@���:�3@-lF���!?+͆s���@Ǵʌ%�ٿQa*E�@���:�3@-lF���!?+͆s���@Ǵʌ%�ٿQa*E�@���:�3@-lF���!?+͆s���@ v8��ٿm��]���@��F���3@.�],�!?
�S��@ v8��ٿm��]���@��F���3@.�],�!?
�S��@ v8��ٿm��]���@��F���3@.�],�!?
�S��@Й�n��ٿ!��m���@Ar��G4@����!?���v��@Й�n��ٿ!��m���@Ar��G4@����!?���v��@Й�n��ٿ!��m���@Ar��G4@����!?���v��@��n���ٿ�9�^��@�A;284@<8J�!?���f�@��n���ٿ�9�^��@�A;284@<8J�!?���f�@��n���ٿ�9�^��@�A;284@<8J�!?���f�@��n���ٿ�9�^��@�A;284@<8J�!?���f�@��y��ٿ�������@�!��3@z��\m�!?���4��@vZ��ٿG��C���@��[�p�3@�'�_C�!?�w�Yx�@vZ��ٿG��C���@��[�p�3@�'�_C�!?�w�Yx�@H~��/�ٿ�K�6|��@�
��4@-%�_�!?^3��@�@O�΃l�ٿ��ȴ���@��ԓ��3@1P�E+�!?�s6�@O�΃l�ٿ��ȴ���@��ԓ��3@1P�E+�!?�s6�@O�΃l�ٿ��ȴ���@��ԓ��3@1P�E+�!?�s6�@lU���ٿ����$E�@\��n�3@-��Z�!?�Է�H�@�>ˮ��ٿ�Q�p�@=OipAE4@�5%�!?D��{�@�>ˮ��ٿ�Q�p�@=OipAE4@�5%�!?D��{�@�>ˮ��ٿ�Q�p�@=OipAE4@�5%�!?D��{�@a�j���ٿd�vS/�@�ѼE4@��Yw�!?D$`@b�@a�j���ٿd�vS/�@�ѼE4@��Yw�!?D$`@b�@a�j���ٿd�vS/�@�ѼE4@��Yw�!?D$`@b�@�&.���ٿQ��a��@MI͓E4@��$}�!?��\�F��@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@�w��e�ٿ��'\���@��4Ȧ;4@�k�-��!?�0����@|:�<��ٿ����~��@���4@�O-c�!?v�U��A�@|:�<��ٿ����~��@���4@�O-c�!?v�U��A�@|:�<��ٿ����~��@���4@�O-c�!?v�U��A�@^'��ٿE��r\$�@�H�/4@��b?�!?�o�mf�@^'��ٿE��r\$�@�H�/4@��b?�!?�o�mf�@t#��ٿ�\�LI�@�.��B�3@o��!?JG�};�@t#��ٿ�\�LI�@�.��B�3@o��!?JG�};�@O�"i��ٿю��X��@|�>&��3@�}/��!?�T0R���@O�"i��ٿю��X��@|�>&��3@�}/��!?�T0R���@'x(�ٿ��U���@ּ尌�3@A�kW�!?R�#��@���v�ٿ��c��@��+�+�3@���^�!?�#'*�@�F����ٿ�<_�@���^��3@�1�[�!?W�S��5�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@��Q+��ٿZ�4>��@�^}y�3@xDR�!?W�Q�x�@�\�#�ٿ�k�z��@·|��4@�w�Ib�!?1K�FT�@�\�#�ٿ�k�z��@·|��4@�w�Ib�!?1K�FT�@�o�Id�ٿ��@���@�mt� 4@:/�̐�!?��T�R��@�o�Id�ٿ��@���@�mt� 4@:/�̐�!?��T�R��@�o�Id�ٿ��@���@�mt� 4@:/�̐�!?��T�R��@�o�Id�ٿ��@���@�mt� 4@:/�̐�!?��T�R��@�o�Id�ٿ��@���@�mt� 4@:/�̐�!?��T�R��@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@m��D�ٿd����@����G4@�Ա���!?\	(��ߕ@I˯Vf�ٿfHSm�@8(���14@��hǐ!?+>�&�@I˯Vf�ٿfHSm�@8(���14@��hǐ!?+>�&�@I˯Vf�ٿfHSm�@8(���14@��hǐ!?+>�&�@I˯Vf�ٿfHSm�@8(���14@��hǐ!?+>�&�@������ٿ��w@�"�@�*�m�M4@TTǙ�!?A�m��Օ@q�����ٿ㑷(c=�@���H(4@8O�S��!?�`�?+ϕ@q�����ٿ㑷(c=�@���H(4@8O�S��!?�`�?+ϕ@q�����ٿ㑷(c=�@���H(4@8O�S��!?�`�?+ϕ@q�����ٿ㑷(c=�@���H(4@8O�S��!?�`�?+ϕ@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@�����ٿ�y�u��@o*�K#4@e?���!?<}WZ��@i��Ӫ�ٿ��ȵ��@E�t3�3@p�QԐ!?��b�[�@i��Ӫ�ٿ��ȵ��@E�t3�3@p�QԐ!?��b�[�@i��Ӫ�ٿ��ȵ��@E�t3�3@p�QԐ!?��b�[�@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@r�"�ٿc��_���@�t�e�3@�#����!?���|��@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@����G�ٿ	T�\��@l����3@�4��]�!?۩����@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��Q�ٿ�#�Gi�@ZNT��4@3o��8�!?ULW`N�@��%��ٿ
�V�'�@�mU��%4@D5VB�!?E䭦��@��VJm�ٿv�f(���@���n4@��<�!?Y(��ԕ@��VJm�ٿv�f(���@���n4@��<�!?Y(��ԕ@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@�TO�F�ٿf;���@3]�u�3@񎴞0�!?�-�h��@s	�e۝ٿ����@��?��3@���!?IXQݕ@s	�e۝ٿ����@��?��3@���!?IXQݕ@s	�e۝ٿ����@��?��3@���!?IXQݕ@s	�e۝ٿ����@��?��3@���!?IXQݕ@s	�e۝ٿ����@��?��3@���!?IXQݕ@��Bv��ٿ^l���*�@��@�"4@4(�n2�!?hÏ@��Bv��ٿ^l���*�@��@�"4@4(�n2�!?hÏ@��Bv��ٿ^l���*�@��@�"4@4(�n2�!?hÏ@CM.l�ٿ·P�i�@[;R`4@�1 �!?��@���@CM.l�ٿ·P�i�@[;R`4@�1 �!?��@���@CM.l�ٿ·P�i�@[;R`4@�1 �!?��@���@CM.l�ٿ·P�i�@[;R`4@�1 �!?��@���@CM.l�ٿ·P�i�@[;R`4@�1 �!?��@���@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@'�Mv�ٿ(�V��B�@8���S4@�`rA�!?��y�@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@S��?�ٿ:f=e��@,FJr44@P�ji�!?���'��@�2�:\�ٿƣx"�3�@tC\t�3@&xIu�!?�w�I?��@�2�:\�ٿƣx"�3�@tC\t�3@&xIu�!?�w�I?��@�2�:\�ٿƣx"�3�@tC\t�3@&xIu�!?�w�I?��@�2�:\�ٿƣx"�3�@tC\t�3@&xIu�!?�w�I?��@�2�:\�ٿƣx"�3�@tC\t�3@&xIu�!?�w�I?��@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@���m�ٿï#�#�@�(y��4@0��J�!?W�)j�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@V-)�D�ٿ
�M~��@���c,34@6�#z�!?&�%�@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@߷�p��ٿ$���@�@�+L=C4@�/4#�!?�����@&��̝ٿ��p��)�@�(W��24@��T���!?7�_��@&��̝ٿ��p��)�@�(W��24@��T���!?7�_��@&��̝ٿ��p��)�@�(W��24@��T���!?7�_��@���J4�ٿ�^�YC�@6ŋ&\x4@)�1���!?��7E"�@���J4�ٿ�^�YC�@6ŋ&\x4@)�1���!?��7E"�@���J4�ٿ�^�YC�@6ŋ&\x4@)�1���!?��7E"�@���J4�ٿ�^�YC�@6ŋ&\x4@)�1���!?��7E"�@���J4�ٿ�^�YC�@6ŋ&\x4@)�1���!?��7E"�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@[��Z��ٿ#����M�@]b�d4@io�I�!?,�)Y�@����[�ٿͦ�((��@�w��4@J�^�!?1.����@����[�ٿͦ�((��@�w��4@J�^�!?1.����@����[�ٿͦ�((��@�w��4@J�^�!?1.����@��@�0�ٿ�@�`B6�@�P�L��3@�2��!?1��s�"�@��@�0�ٿ�@�`B6�@�P�L��3@�2��!?1��s�"�@��@�0�ٿ�@�`B6�@�P�L��3@�2��!?1��s�"�@��:���ٿ��]\�@�<m#K�3@�ʱ�!�!?���x[,�@��:���ٿ��]\�@�<m#K�3@�ʱ�!�!?���x[,�@��:���ٿ��]\�@�<m#K�3@�ʱ�!�!?���x[,�@��:���ٿ��]\�@�<m#K�3@�ʱ�!�!?���x[,�@��:���ٿ��]\�@�<m#K�3@�ʱ�!�!?���x[,�@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@`.�{�ٿin5�l�@J�� 4@�o{��!?
K��ѕ@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@d�\О�ٿ�����@R�J44@���!?]�JQ@�@q}��%�ٿ�ׯ&��@9�A4@ϟ���!?!��Ѷ��@��'�E�ٿ����`��@����QD4@�}!ڻ�!?� 9�ß�@��'�E�ٿ����`��@����QD4@�}!ڻ�!?� 9�ß�@Чq�B�ٿ�1-��@��i�S4@62G�!?���_a�@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@"롳q�ٿ�L#B��@J�\q.4@�s�5Z�!?#��9Օ@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@d�_��ٿ�';V���@"�F	�"4@�T%�!?"/�JA͕@b� �ٿ~��U�@����3@JyAԽ�!?����@b� �ٿ~��U�@����3@JyAԽ�!?����@b� �ٿ~��U�@����3@JyAԽ�!?����@b� �ٿ~��U�@����3@JyAԽ�!?����@b� �ٿ~��U�@����3@JyAԽ�!?����@��ez�ٿ���0��@ ��4@�-	�j�!?d�n�J7�@��ez�ٿ���0��@ ��4@�-	�j�!?d�n�J7�@��ez�ٿ���0��@ ��4@�-	�j�!?d�n�J7�@��ez�ٿ���0��@ ��4@�-	�j�!?d�n�J7�@�iΗٿ��Q�Z��@9�.TJK4@��Vc�!?;0��{�@�iΗٿ��Q�Z��@9�.TJK4@��Vc�!?;0��{�@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@R:ρ��ٿ-I�L�@Q(�Ɨ'4@�Qݐ!?����@��5�ٿ�6a�W��@TH�2�X4@)�J�f�!?ɚ䍙ϕ@��5�ٿ�6a�W��@TH�2�X4@)�J�f�!?ɚ䍙ϕ@��5�ٿ�6a�W��@TH�2�X4@)�J�f�!?ɚ䍙ϕ@��5�ٿ�6a�W��@TH�2�X4@)�J�f�!?ɚ䍙ϕ@���<�ٿD��ok�@G����14@�}R�o�!?D��Ѐ�@���<�ٿD��ok�@G����14@�}R�o�!?D��Ѐ�@���<�ٿD��ok�@G����14@�}R�o�!?D��Ѐ�@���<�ٿD��ok�@G����14@�}R�o�!?D��Ѐ�@���<�ٿD��ok�@G����14@�}R�o�!?D��Ѐ�@-�(���ٿڼg��@Η���I4@q���u�!?J�#T↕@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@���2��ٿ�Ix��)�@�]š'�3@��䶐!?.���b��@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@L���,�ٿ���$F�@y�&"4@��'�!?�	�ʕ@�*�t�ٿ�_Mzֿ�@�m��3@��^!?F����@�*�t�ٿ�_Mzֿ�@�m��3@��^!?F����@���.��ٿ�z��7�@����[�3@ʐ"��!?!v�JM�@���.��ٿ�z��7�@����[�3@ʐ"��!?!v�JM�@���.��ٿ�z��7�@����[�3@ʐ"��!?!v�JM�@���.��ٿ�z��7�@����[�3@ʐ"��!?!v�JM�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@K�a�ٿ��0� �@�+�4@��?�U�!?�,3��Q�@�o���ٿw�����@�rےX*4@�r.X�!?���&��@�o���ٿw�����@�rےX*4@�r.X�!?���&��@���r�ٿ������@�y�4@��h>�!?�/�#�@���r�ٿ������@�y�4@��h>�!?�/�#�@�W���ٿD�r���@m�d��=4@�Q�9w�!?m��,o�@�W���ٿD�r���@m�d��=4@�Q�9w�!?m��,o�@�W���ٿD�r���@m�d��=4@�Q�9w�!?m��,o�@1����ٿ���s��@!N����3@�[
=t�!?��q�H�@1����ٿ���s��@!N����3@�[
=t�!?��q�H�@1����ٿ���s��@!N����3@�[
=t�!?��q�H�@1����ٿ���s��@!N����3@�[
=t�!?��q�H�@1����ٿ���s��@!N����3@�[
=t�!?��q�H�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@�y�.��ٿ��2�%@�@��%O�4@.8�k��!?�R��q�@/�ᠶ�ٿt)����@^�DUp4@~�~�$�!?�{��H�@�����ٿN&��<��@c:9Y�*4@D�ɓ�!?��99: �@�����ٿN&��<��@c:9Y�*4@D�ɓ�!?��99: �@�����ٿN&��<��@c:9Y�*4@D�ɓ�!?��99: �@�����ٿN&��<��@c:9Y�*4@D�ɓ�!?��99: �@�.1���ٿ�z�l��@M�l=4@u`%�ߐ!?�X��؃�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@?:���ٿ6*	���@�2���04@��A�!?��[�-u�@ƇeD��ٿ)��s��@�-Z3*4@���!?O}�L�@����ٿ�G��F��@��B�;4@�bL��!?}Q,��ڕ@����ٿ�G��F��@��B�;4@�bL��!?}Q,��ڕ@����ٿ�G��F��@��B�;4@�bL��!?}Q,��ڕ@����ٿ�G��F��@��B�;4@�bL��!?}Q,��ڕ@z�m��ٿFtP`���@�(�+�g4@hA�'�!?��[���@z�m��ٿFtP`���@�(�+�g4@hA�'�!?��[���@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@��/���ٿH�V0$�@���04@�N�V�!?�[jg�:�@�_��ٿ3J�k~��@��
4@1�'Z�!?��: �W�@�_��ٿ3J�k~��@��
4@1�'Z�!?��: �W�@�_��ٿ3J�k~��@��
4@1�'Z�!?��: �W�@�_��ٿ3J�k~��@��
4@1�'Z�!?��: �W�@�_��ٿ3J�k~��@��
4@1�'Z�!?��: �W�@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@\-�n��ٿU�D̼�@�`�-��3@�����!?�� B
 �@i�L��ٿ��8����@���3@�r�ߔ�!?N�6�n5�@i�L��ٿ��8����@���3@�r�ߔ�!?N�6�n5�@i�L��ٿ��8����@���3@�r�ߔ�!?N�6�n5�@i�L��ٿ��8����@���3@�r�ߔ�!?N�6�n5�@i�L��ٿ��8����@���3@�r�ߔ�!?N�6�n5�@�L���ٿa��H�6�@z�֎�3@�4�Ċ�!?2HPT�@�L���ٿa��H�6�@z�֎�3@�4�Ċ�!?2HPT�@�L���ٿa��H�6�@z�֎�3@�4�Ċ�!?2HPT�@�L���ٿa��H�6�@z�֎�3@�4�Ċ�!?2HPT�@�L���ٿa��H�6�@z�֎�3@�4�Ċ�!?2HPT�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@�BU-̠ٿ�ڛ�%�@-�@*4@��=�!?r�7x2�@��T}��ٿ����2�@�S+���3@�h-�^�!?D����b�@��T}��ٿ����2�@�S+���3@�h-�^�!?D����b�@��T}��ٿ����2�@�S+���3@�h-�^�!?D����b�@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@��:���ٿw�'���@(-�+�4@2�PR�!?�u�g��@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@H1���ٿ�`���@V>4@��$�J�!?��4-p�@���I�ٿ�����@B־���3@�i2n�!?�D�� �@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��Hc^�ٿ@ �!�@��c3��3@e�|Q��!?�dߢЕ@��mʞٿ����s��@wV
�;4@Y��-�!?�8Z܎ԕ@��mʞٿ����s��@wV
�;4@Y��-�!?�8Z܎ԕ@�o��ٿ	k&!��@�;�!4@��'"��!?l��Y�@�o��ٿ	k&!��@�;�!4@��'"��!?l��Y�@�o��ٿ	k&!��@�;�!4@��'"��!?l��Y�@�!���ٿ �*Nk�@`�A��"4@Cc%c�!?�̑��@�!���ٿ �*Nk�@`�A��"4@Cc%c�!?�̑��@�!���ٿ �*Nk�@`�A��"4@Cc%c�!?�̑��@d��|�ٿ�1����@?g`a,�3@Lj[v�!?8�Mͬ�@d��|�ٿ�1����@?g`a,�3@Lj[v�!?8�Mͬ�@d��|�ٿ�1����@?g`a,�3@Lj[v�!?8�Mͬ�@x�PUy�ٿL�k�c!�@��w*�4@K[�Gq�!?���3��@x�PUy�ٿL�k�c!�@��w*�4@K[�Gq�!?���3��@�v�� �ٿ�	�9���@��C^4@&V�Β�!?!KL�|��@�v�� �ٿ�	�9���@��C^4@&V�Β�!?!KL�|��@�v�� �ٿ�	�9���@��C^4@&V�Β�!?!KL�|��@e���ٿ������@=O�4@ӹ�T��!?��5D��@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@���ٿ\�J(��@���@�3@ �����!?~3�[Ĉ�@u1�נٿC� ��$�@���?�3@�d1�ǐ!??	LR�@` ��ʞٿSM��@��e�|�3@�/sͷ�!?
��D�1�@�R�s�ٿ{������@J}�3@�	�(��!?5V-%�@�R�s�ٿ{������@J}�3@�	�(��!?5V-%�@�R�s�ٿ{������@J}�3@�	�(��!?5V-%�@?j�sm�ٿ��z'�@� �A��3@y��g��!?8'd����@��zK�ٿ][]�K�@q��{�3@�5�d��!?��<�W�@^d��_�ٿl��q�@�R�b�4@���l �!?=8g@	��@^d��_�ٿl��q�@�R�b�4@���l �!?=8g@	��@{Z|�r�ٿ��Ghʯ�@�L�!.4@TB�!?��qb�p�@�|��ٿ��}�6��@t��ޤ54@Q�ð�!?�+�ʋ��@�|��ٿ��}�6��@t��ޤ54@Q�ð�!?�+�ʋ��@�|��ٿ��}�6��@t��ޤ54@Q�ð�!?�+�ʋ��@]$ż�ٿ��w(��@��1Z��3@�T�6m�!?���83�@��pzϟٿ,����@XsT�5 4@:�Ь��!?��W��@��pzϟٿ,����@XsT�5 4@:�Ь��!?��W��@��pzϟٿ,����@XsT�5 4@:�Ь��!?��W��@��pzϟٿ,����@XsT�5 4@:�Ь��!?��W��@.����ٿ�{?g��@[�o��4@_�qjl�!?7��=�@.����ٿ�{?g��@[�o��4@_�qjl�!?7��=�@��.���ٿ�o�*!��@�y�">4@�pC��!?�kF����@��.���ٿ�o�*!��@�y�">4@�pC��!?�kF����@��.���ٿ�o�*!��@�y�">4@�pC��!?�kF����@��.���ٿ�o�*!��@�y�">4@�pC��!?�kF����@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�i���ٿτ��;X�@T����3@���Ƀ�!?�~�(��@�{�W0�ٿ��.[��@�`z�?4@��r��!?`\�]��@�{�W0�ٿ��.[��@�`z�?4@��r��!?`\�]��@�{�W0�ٿ��.[��@�`z�?4@��r��!?`\�]��@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@9*P=��ٿ��-B��@�{���4@)���a�!?@��cĕ@�R���ٿ6#Iџ��@u���q,4@�/g�!?���o��@�R���ٿ6#Iџ��@u���q,4@�/g�!?���o��@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@:-Ebܞٿox�5���@)���#4@�XUg��!?(i0mŕ@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@ ����ٿ�Ħ��@c��:�3@B���!?�*MH/N�@6���ٿ��F����@8��"��3@�d�x�!?�� ���@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@���ٿ����@��@�,��3@���^�!?�N��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@�d-&�ٿ������@^�Q��3@��=`�!?�eq�U��@}�ýњٿ��tY׸�@�RW�!4@z��3 �!?x��k]ʕ@}�ýњٿ��tY׸�@�RW�!4@z��3 �!?x��k]ʕ@�"�Tp�ٿ�B�-�@jE�\<4@��(3�!?2h����@�"�Tp�ٿ�B�-�@jE�\<4@��(3�!?2h����@�"�Tp�ٿ�B�-�@jE�\<4@��(3�!?2h����@�"�Tp�ٿ�B�-�@jE�\<4@��(3�!?2h����@k�b!��ٿ�9�n+�@�� &4@e�C#�!?-T2��@��#��ٿ�?X���@���j�%4@]�~;�!?��m��,�@��#��ٿ�?X���@���j�%4@]�~;�!?��m��,�@Ǜ"���ٿ�~,���@(M�d��3@�	�y�!?���=�@Q��Y��ٿ��Gۅ��@60��Q4@�L����!?�j��g�@Q��Y��ٿ��Gۅ��@60��Q4@�L����!?�j��g�@Q��Y��ٿ��Gۅ��@60��Q4@�L����!?�j��g�@<1�d��ٿ�d�k<-�@A)���4@���^�!?���D3�@<1�d��ٿ�d�k<-�@A)���4@���^�!?���D3�@<1�d��ٿ�d�k<-�@A)���4@���^�!?���D3�@c�Z�ѝٿ O�IE\�@6�"��	4@���<|�!?x�#���@c�Z�ѝٿ O�IE\�@6�"��	4@���<|�!?x�#���@c�Z�ѝٿ O�IE\�@6�"��	4@���<|�!?x�#���@��r2V�ٿ�3>���@6�}���3@T���!?��?!h%�@��r2V�ٿ�3>���@6�}���3@T���!?��?!h%�@&�}{�ٿ��L��@w�{�74@�ǐ!?��#���@Jħ'�ٿ��6�0��@dy��4@��;d��!?I�.�t:�@Jħ'�ٿ��6�0��@dy��4@��;d��!?I�.�t:�@Jħ'�ٿ��6�0��@dy��4@��;d��!?I�.�t:�@Jħ'�ٿ��6�0��@dy��4@��;d��!?I�.�t:�@���j�ٿ�	A���@��
iL4@XxD��!?��dw�@���j�ٿ�	A���@��
iL4@XxD��!?��dw�@����ٿ�v$y���@3���Q$4@-�Ѐې!?f�a!us�@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@~XӲZ�ٿB=�b��@w��w74@��F�ߐ!?+��䜕@P�V- �ٿ�������@����j14@� ʓ��!?��L�7�@P�V- �ٿ�������@����j14@� ʓ��!?��L�7�@P�V- �ٿ�������@����j14@� ʓ��!?��L�7�@*�^O��ٿ.��5;��@�l�A4@��'{��!?��8�9�@*�^O��ٿ.��5;��@�l�A4@��'{��!?��8�9�@*�^O��ٿ.��5;��@�l�A4@��'{��!?��8�9�@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@�sM�g�ٿH�I���@�l��"4@a��[z�!?Ğ��l��@!��Q�ٿ b���Z�@��wx]�3@��8IJ�!?��0��@!��Q�ٿ b���Z�@��wx]�3@��8IJ�!?��0��@!��Q�ٿ b���Z�@��wx]�3@��8IJ�!?��0��@!��Q�ٿ b���Z�@��wx]�3@��8IJ�!?��0��@�7�4̛ٿ]�
�i�@��?4@�t�_�!?���*ӹ�@�7�4̛ٿ]�
�i�@��?4@�t�_�!?���*ӹ�@�7�4̛ٿ]�
�i�@��?4@�t�_�!?���*ӹ�@N6H���ٿ�H�y��@�>��24@�K,I�!?V��c]�@N6H���ٿ�H�y��@�>��24@�K,I�!?V��c]�@N6H���ٿ�H�y��@�>��24@�K,I�!?V��c]�@N6H���ٿ�H�y��@�>��24@�K,I�!?V��c]�@N6H���ٿ�H�y��@�>��24@�K,I�!?V��c]�@�t�z�ٿ�����@(�?{*14@뉆2l�!?����*�@�t�z�ٿ�����@(�?{*14@뉆2l�!?����*�@�t�z�ٿ�����@(�?{*14@뉆2l�!?����*�@�t�z�ٿ�����@(�?{*14@뉆2l�!?����*�@Z4zW�ٿ�w��@a'�T�84@��jh�!?3�F^��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�n�a��ٿx�zO���@�!u���3@��Eh��!?�<�!��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@�Ձ�b�ٿ{�k�r��@�T2�4@zdD^�!?C̨�V��@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@A��"-�ٿ(l����@ �N Z(4@gp
w�!?P@����@s����ٿN��fn��@����4@�}b�_�!?|Ǖ��7�@��0|�ٿ6�4���@	7��~�3@!����!?)��L��@E2Md��ٿͥ��1��@� �"�3@w��~��!?:j}t�Õ@���9�ٿ�Fs^��@��B��3@j0� �!?y��U�{�@���9�ٿ�Fs^��@��B��3@j0� �!?y��U�{�@UH�ڛٿm��-���@
��T,4@��
�!?�b�%~`�@�.���ٿ���{3�@����N4@Ѳ�V�!?���ۗ�@�.���ٿ���{3�@����N4@Ѳ�V�!?���ۗ�@�.���ٿ���{3�@����N4@Ѳ�V�!?���ۗ�@�.���ٿ���{3�@����N4@Ѳ�V�!?���ۗ�@�v��ٿ��yh�%�@��8}':4@�\�;n�!?��!��8�@�>Zc�ٿ�t��A��@B؋�3@�*����!?����q!�@�>Zc�ٿ�t��A��@B؋�3@�*����!?����q!�@�>Zc�ٿ�t��A��@B؋�3@�*����!?����q!�@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@��Da�ٿ�_�T_u�@�h5��3@;�t��!?��5u���@�&_��ٿ�1�� ��@��S��3@�#�!?���H�n�@)���|�ٿ
Ц�5��@B;g�4@`��\�!?
s��ؖ@)���|�ٿ
Ц�5��@B;g�4@`��\�!?
s��ؖ@;]�m��ٿz,���@�@�0V�84@T�Vjp�!?7-�	J��@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@4ω�!�ٿ 6>Y���@�����'4@"�+�P�!?�O�R���@q��S��ٿ�����@�~Ǆ(4@Ow_0�!?�9�P�@���Ԭ�ٿ����^�@�����4@M-��r�!?
�\V��@���Ԭ�ٿ����^�@�����4@M-��r�!?
�\V��@���Ԭ�ٿ����^�@�����4@M-��r�!?
�\V��@���Ԭ�ٿ����^�@�����4@M-��r�!?
�\V��@���Ԭ�ٿ����^�@�����4@M-��r�!?
�\V��@6�k֚ٿޚ<(���@��V�n+4@�oJ.��!?�{&���@���LY�ٿ~  ��S�@K�S��4@���!?�W�D�q�@d}�a�ٿ�{R0�@�ڰ��3@b��S�!?�sЁgS�@d}�a�ٿ�{R0�@�ڰ��3@b��S�!?�sЁgS�@d}�a�ٿ�{R0�@�ڰ��3@b��S�!?�sЁgS�@ў;�x�ٿ��-�@XB45�3@���!�!?n�ꞇ͕@ў;�x�ٿ��-�@XB45�3@���!�!?n�ꞇ͕@��¸��ٿ�;{�@�;�!��3@+:�y�!?��x����@���Ҝٿ�mʹ�@�Y�Y��3@v�(
;�!?=ʓ�}Е@���Ҝٿ�mʹ�@�Y�Y��3@v�(
;�!?=ʓ�}Е@���Ҝٿ�mʹ�@�Y�Y��3@v�(
;�!?=ʓ�}Е@���Ҝٿ�mʹ�@�Y�Y��3@v�(
;�!?=ʓ�}Е@��^��ٿ���A�@ț^�+4@l.Y�m�!?d���x"�@��^��ٿ���A�@ț^�+4@l.Y�m�!?d���x"�@��^��ٿ���A�@ț^�+4@l.Y�m�!?d���x"�@��^��ٿ���A�@ț^�+4@l.Y�m�!?d���x"�@_��fI�ٿ�<&`�H�@��/@4@yJ-�M�!?�����@_��fI�ٿ�<&`�H�@��/@4@yJ-�M�!?�����@_��fI�ٿ�<&`�H�@��/@4@yJ-�M�!?�����@_��fI�ٿ�<&`�H�@��/@4@yJ-�M�!?�����@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@C[󑶚ٿ�!7�W%�@
T�#4@{FD�!?\�z�_�@��b}�ٿr�����@����3@���s�!?툤���@��b}�ٿr�����@����3@���s�!?툤���@��b}�ٿr�����@����3@���s�!?툤���@��b}�ٿr�����@����3@���s�!?툤���@��b}�ٿr�����@����3@���s�!?툤���@��b}�ٿr�����@����3@���s�!?툤���@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@����ٿ��<f��@+�^�K&4@�[�R�!?S�	��@�.�Q�ٿ���q�@�ӸJ94@���!�!?xOH���@�.�Q�ٿ���q�@�ӸJ94@���!�!?xOH���@�.�Q�ٿ���q�@�ӸJ94@���!�!?xOH���@5�>�f�ٿg�X�c|�@H�R*4@�n�m�!?�)WP�ӕ@5�>�f�ٿg�X�c|�@H�R*4@�n�m�!?�)WP�ӕ@L�2�ٿL�%��@���)4@ٔaQ�!?�F�`�@<ig���ٿ ��o�@İ�g4E4@���'�!?]�g���@<ig���ٿ ��o�@İ�g4E4@���'�!?]�g���@<ig���ٿ ��o�@İ�g4E4@���'�!?]�g���@�U'�ٿ��.Uw�@��84@"�`~�!? ������@����E�ٿ�2u���@�_[K<4@_o�F�!?�,kq�@����E�ٿ�2u���@�_[K<4@_o�F�!?�,kq�@����E�ٿ�2u���@�_[K<4@_o�F�!?�,kq�@����E�ٿ�2u���@�_[K<4@_o�F�!?�,kq�@����E�ٿ�2u���@�_[K<4@_o�F�!?�,kq�@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@�"�G��ٿ�ڡ��@��)C	%4@�-��t�!?�v
���@8�!.]�ٿ�U�*�Z�@�-@�4@ Hx�|�!?�^ �᜕@8�!.]�ٿ�U�*�Z�@�-@�4@ Hx�|�!?�^ �᜕@8�!.]�ٿ�U�*�Z�@�-@�4@ Hx�|�!?�^ �᜕@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@2"�R�ٿR��8�@�J%(�3@J�ZuL�!?�����@�8��Ҟٿ�D�%���@�v2��3@�}�~�!?��w����@�8��Ҟٿ�D�%���@�v2��3@�}�~�!?��w����@�8��Ҟٿ�D�%���@�v2��3@�}�~�!?��w����@�8��Ҟٿ�D�%���@�v2��3@�}�~�!?��w����@�_��Ρٿ���"�@�)-�"�3@*hNꔐ!?�
�a��@�_��Ρٿ���"�@�)-�"�3@*hNꔐ!?�
�a��@�_��Ρٿ���"�@�)-�"�3@*hNꔐ!?�
�a��@=~���ٿ1��X��@�F%Z��3@��m2��!?D��ѕ@=~���ٿ1��X��@�F%Z��3@��m2��!?D��ѕ@�R,뷞ٿ�v.�i�@(�tWn�3@SC��!?�EA/f@�@�R,뷞ٿ�v.�i�@(�tWn�3@SC��!?�EA/f@�@�R,뷞ٿ�v.�i�@(�tWn�3@SC��!?�EA/f@�@�R,뷞ٿ�v.�i�@(�tWn�3@SC��!?�EA/f@�@Sȷ�,�ٿְ=��%�@��b��+4@V��U�!?P�H��8�@Sȷ�,�ٿְ=��%�@��b��+4@V��U�!?P�H��8�@�|�O�ٿ�2��o!�@4ZO:�>4@S��*�!?;�N���@��g���ٿ��HI��@kE�O�F4@bv|^�!?� �����@��g���ٿ��HI��@kE�O�F4@bv|^�!?� �����@��g���ٿ��HI��@kE�O�F4@bv|^�!?� �����@��g���ٿ��HI��@kE�O�F4@bv|^�!?� �����@C�I~f�ٿWg�W���@��rn�-4@k��}T�!?�b����@C�I~f�ٿWg�W���@��rn�-4@k��}T�!?�b����@C�I~f�ٿWg�W���@��rn�-4@k��}T�!?�b����@C�I~f�ٿWg�W���@��rn�-4@k��}T�!?�b����@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@yK9��ٿ"�2M��@`���4@��j�\�!?N&���@}�z�ʘٿ~i�A���@Z����I4@�7𣐐!?�����@}�z�ʘٿ~i�A���@Z����I4@�7𣐐!?�����@ݞ8$�ٿ��dv���@h���84@L�Kk�!?v�fו@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@M��T�ٿ@�i8D�@��֟G)4@~Z��!?��?H<�@/m�Δٿm	�ye��@��	�24@�%����!?X@��@�aX�E�ٿǓ�'��@3��]@4@>�#t�!?N,����@�aX�E�ٿǓ�'��@3��]@4@>�#t�!?N,����@���L�ٿ����(�@�o��D4@��&I9�!?&q�?C�@���L�ٿ����(�@�o��D4@��&I9�!?&q�?C�@���L�ٿ����(�@�o��D4@��&I9�!?&q�?C�@���L�ٿ����(�@�o��D4@��&I9�!?&q�?C�@���L�ٿ����(�@�o��D4@��&I9�!?&q�?C�@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@>��S�ٿD���@nS��� 4@+�QUD�!?��N���@�p�O�ٿ�L'��@�`[��L4@��� �!?U6��Ǖ@�p�O�ٿ�L'��@�`[��L4@��� �!?U6��Ǖ@�p�O�ٿ�L'��@�`[��L4@��� �!?U6��Ǖ@�p�%��ٿH�.z��@���U�4@���K�!?����S2�@�p�%��ٿH�.z��@���U�4@���K�!?����S2�@�p�%��ٿH�.z��@���U�4@���K�!?����S2�@�p�%��ٿH�.z��@���U�4@���K�!?����S2�@�p�%��ٿH�.z��@���U�4@���K�!?����S2�@^ڣ�ܠٿ�:I���@��'�4@�ĝd�!?���Qc\�@^ڣ�ܠٿ�:I���@��'�4@�ĝd�!?���Qc\�@M�Lg��ٿv;u�Y�@����24@ӂz�i�!?@�2�?f�@M�Lg��ٿv;u�Y�@����24@ӂz�i�!?@�2�?f�@M�Lg��ٿv;u�Y�@����24@ӂz�i�!?@�2�?f�@M�Lg��ٿv;u�Y�@����24@ӂz�i�!?@�2�?f�@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@������ٿ��',h�@�O@X4@�s�;��!?��� ��@���>f�ٿ���M��@�f��C4@'�$?��!?�ա�6�@�1��Ƙٿ�ه�dW�@��oK�4@� ���!?;%�D���@{��L
�ٿU�@��@�+U��3@����!?1#9@8ە@HV���ٿHGu���@�	���3@dѣB��!?�D|m˕@HV���ٿHGu���@�	���3@dѣB��!?�D|m˕@HV���ٿHGu���@�	���3@dѣB��!?�D|m˕@HV���ٿHGu���@�	���3@dѣB��!?�D|m˕@HV���ٿHGu���@�	���3@dѣB��!?�D|m˕@����ٿW�i���@�j6$4@z����!?8E�c<��@����ٿW�i���@�j6$4@z����!?8E�c<��@�����ٿ��l1Y�@�W�X�4@N�F��!?�4ї�ʕ@�t	P�ٿ���4��@޺�S4@�4��Ӑ!?w5�#�@�t	P�ٿ���4��@޺�S4@�4��Ӑ!?w5�#�@�t	P�ٿ���4��@޺�S4@�4��Ӑ!?w5�#�@�/4M˚ٿQ�����@��"_�F4@9x���!?����-<�@�/4M˚ٿQ�����@��"_�F4@9x���!?����-<�@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@O���ٿ���}t��@L��e\T4@D�	ק�!?��x@oߕ@�M�i�ٿp�P��v�@#��<4@��	���!?��}����@�M�i�ٿp�P��v�@#��<4@��	���!?��}����@�M�i�ٿp�P��v�@#��<4@��	���!?��}����@�M�i�ٿp�P��v�@#��<4@��	���!?��}����@�M�i�ٿp�P��v�@#��<4@��	���!?��}����@��A�ٿeP�"�@%�+��?4@��.���!?�ju��|�@��A�ٿeP�"�@%�+��?4@��.���!?�ju��|�@��A�ٿeP�"�@%�+��?4@��.���!?�ju��|�@��A�ٿeP�"�@%�+��?4@��.���!?�ju��|�@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@a%��1�ٿ�9=~g�@�t��p(4@Pڷ�W�!?�֙����@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@q�	a��ٿw����@�&��64@��V�x�!?q�O*L��@Fx�o͘ٿu*�f�@���4@�x�3�!?%�:+�@�GV��ٿ���e��@����3@+��X�!?�wJ{C�@�GV��ٿ���e��@����3@+��X�!?�wJ{C�@v���ٿ�?�-�@�x�k�3@���Q�!?טI��9�@v���ٿ�?�-�@�x�k�3@���Q�!?טI��9�@v���ٿ�?�-�@�x�k�3@���Q�!?טI��9�@v���ٿ�?�-�@�x�k�3@���Q�!?טI��9�@�v����ٿȗ����@��n���3@,�Y�}�!?o��y��@���u�ٿ�|���@ ���p�3@V��W
�!?�HJ)���@���u�ٿ�|���@ ���p�3@V��W
�!?�HJ)���@2r�~�ٿ{�b.�t�@�EtAu4@&�H�s�!?����@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@�e���ٿ�N��x�@@ܳ��3@-�㉀�!?&�2�ӕ@B~�!�ٿ0�ܳ0�@��!�,4@��Y�!?�=�Gb��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@+֜B��ٿ*i����@�{޳�\4@?�~�f�!?ÊX��@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@������ٿa\7�w�@��\�I4@�-W�c�!?+j����@�4%�ٿ�X@�2�@ruoó4@�{{>�!?!��@�@�4%�ٿ�X@�2�@ruoó4@�{{>�!?!��@�@�4%�ٿ�X@�2�@ruoó4@�{{>�!?!��@�@�ݩ`�ٿ���N���@}��{*4@�\p0�!?n���&�@�ݩ`�ٿ���N���@}��{*4@�\p0�!?n���&�@�ݩ`�ٿ���N���@}��{*4@�\p0�!?n���&�@ٱ5b�ٿ3���<l�@��4���3@����#�!?�cn��@9�V�ٿ$<��J�@��A��3@49��C�!?��ǭ�3�@9�ڞٿ�m�Z]��@���\g4@VS�!?���0�@9�ڞٿ�m�Z]��@���\g4@VS�!?���0�@9�ڞٿ�m�Z]��@���\g4@VS�!?���0�@9�ڞٿ�m�Z]��@���\g4@VS�!?���0�@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@��<�ٿ�6dJ��@�5�;4@��#/�!?T!��@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@�7�	˞ٿ��K�@��@�ë�D4@��@�!?��zil�@n/�n�ٿ�aE��@>��L�C4@�� |V�!?f��w7�@n/�n�ٿ�aE��@>��L�C4@�� |V�!?f��w7�@n/�n�ٿ�aE��@>��L�C4@�� |V�!?f��w7�@n/�n�ٿ�aE��@>��L�C4@�� |V�!?f��w7�@�F�LT�ٿ2��y= �@�&�R�U4@H.�[�!?��0>�&�@�F�LT�ٿ2��y= �@�&�R�U4@H.�[�!?��0>�&�@�F�LT�ٿ2��y= �@�&�R�U4@H.�[�!?��0>�&�@�F�LT�ٿ2��y= �@�&�R�U4@H.�[�!?��0>�&�@�F�LT�ٿ2��y= �@�&�R�U4@H.�[�!?��0>�&�@�!V��ٿ��)��e�@��%r8\4@�_�ɕ�!?s�p��@<δ�<�ٿ��LgRk�@,=��z4@�7���!?�O�9��@<δ�<�ٿ��LgRk�@,=��z4@�7���!?�O�9��@<δ�<�ٿ��LgRk�@,=��z4@�7���!?�O�9��@��7qԤٿ�u´{�@��@��-4@bA��'�!?�bw�o��@��7qԤٿ�u´{�@��@��-4@bA��'�!?�bw�o��@�O�.&�ٿeL��/C�@_�i@4@z)c-�!?�ԙ��@�O�.&�ٿeL��/C�@_�i@4@z)c-�!?�ԙ��@���v�ٿ�Ǆe���@w�@�4@P��'�!?N���fd�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@�"�y��ٿ$�9�e�@47�/\4@�e92�!?�tYQM�@��Vv�ٿ�Y[�V�@�mD��4@��08D�!?�/�w�!�@+�ٿ�Ԙ���@�'�34@ۺ��!?PT����@+�ٿ�Ԙ���@�'�34@ۺ��!?PT����@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@�D�@�ٿ+�����@@޶tW4@:MBO�!?,��P�$�@����6�ٿC��wa�@sA:gNV4@����!?ز�w�@����6�ٿC��wa�@sA:gNV4@����!?ز�w�@����6�ٿC��wa�@sA:gNV4@����!?ز�w�@����6�ٿC��wa�@sA:gNV4@����!?ز�w�@,���B�ٿu1���2�@W,M<eL4@R[k]�!?�)N��@,���B�ٿu1���2�@W,M<eL4@R[k]�!?�)N��@,���B�ٿu1���2�@W,M<eL4@R[k]�!?�)N��@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@?��!-�ٿ��}�@�3�U4@9��ϒ�!?P�f���@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@�GJ�3�ٿ!��8N�@��z�}34@7VAU�!?�K8�)�@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@��@_y�ٿ]�:�z��@	�»P 4@��aIO�!?��ӻ���@�����ٿ6�΄���@�_V�?L4@�o���!?�IO�Õ@�����ٿ6�΄���@�_V�?L4@�o���!?�IO�Õ@�����ٿ6�΄���@�_V�?L4@�o���!?�IO�Õ@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@唌���ٿ�������@���W4@\3�tw�!?�����@�<	�ٿ�Q���y�@Ǎ��I4@�/�a�!?��6��@�@�К�=�ٿ��[���@�<Չ2F4@�l��z�!?L+�Lו@s�^{��ٿ�)9���@U2�#+4@擕l�!?p)�]���@��/���ٿI{X
C�@����4@j^0�C�!?�W��{��@�	��ڜٿr�V~w��@�Kc�%;4@��<�!?��È���@�	��ڜٿr�V~w��@�Kc�%;4@��<�!?��È���@�	��ڜٿr�V~w��@�Kc�%;4@��<�!?��È���@�	��ڜٿr�V~w��@�Kc�%;4@��<�!?��È���@�	��ڜٿr�V~w��@�Kc�%;4@��<�!?��È���@��h�"�ٿ�����@t�Rj4@�|��0�!?m�b	:�@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@9x�� �ٿ?�Ƈ\�@�M� M4@�,� P�!?��(b�ȕ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@�����ٿ�D���s�@��\ 4@�)	`j�!?˸���Õ@i�X{��ٿ�l���@f��%4@���ce�!?3�v9�~�@�f)���ٿߜF�?#�@�i�OeC4@��"���!?��ӂ�@�f)���ٿߜF�?#�@�i�OeC4@��"���!?��ӂ�@���]]�ٿh�!F0��@8��
,84@�b$��!?�i��@���]]�ٿh�!F0��@8��
,84@�b$��!?�i��@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@��dD�ٿ��ik��@��-��4@6���F�!?��D�V�@~��7��ٿ?�v6�@M2�nM 4@?��.�!?/5��Е@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�#���ٿ2%4RjR�@e���3@�j�^4�!?Ta��ӕ@�I1,�ٿ�����y�@�c$*�3@�lP�\�!?�9�v�@���9ɛٿ����p�@y(Ivn4@��ѥ��!?Z�o��@Gص���ٿ��Σ��@�DP� 4@'�ݘ��!?!�Z���@Gص���ٿ��Σ��@�DP� 4@'�ݘ��!?!�Z���@Gص���ٿ��Σ��@�DP� 4@'�ݘ��!?!�Z���@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�
R(�ٿɡrF�@�J|�I4@��xP��!?V�����@�W��ٿ2%����@���4�
4@�]��!?0����@�W��ٿ2%����@���4�
4@�]��!?0����@Cv lA�ٿ�%��CV�@A�%i�4@z��I�!?h�6�*��@Cv lA�ٿ�%��CV�@A�%i�4@z��I�!?h�6�*��@Cv lA�ٿ�%��CV�@A�%i�4@z��I�!?h�6�*��@Cv lA�ٿ�%��CV�@A�%i�4@z��I�!?h�6�*��@�C�j��ٿ F���a�@D�%!4@#�@�[�!?�Q��8�@�C�j��ٿ F���a�@D�%!4@#�@�[�!?�Q��8�@�̩x��ٿ{s{ �%�@����64@�/?�H�!?��6�@�̩x��ٿ{s{ �%�@����64@�/?�H�!?��6�@.�<g�ٿ鸑\K!�@D���|)4@Nǈ� �!?%�ޏ�Е@.�<g�ٿ鸑\K!�@D���|)4@Nǈ� �!?%�ޏ�Е@.�<g�ٿ鸑\K!�@D���|)4@Nǈ� �!?%�ޏ�Е@.�<g�ٿ鸑\K!�@D���|)4@Nǈ� �!?%�ޏ�Е@�Q�e�ٿ̩э���@SJy��4@gL�r!�!?���c��@�Q�e�ٿ̩э���@SJy��4@gL�r!�!?���c��@�Q�e�ٿ̩э���@SJy��4@gL�r!�!?���c��@ލ&�C�ٿ�i��@��ΰ�4@{Oh8/�!?Y����@ލ&�C�ٿ�i��@��ΰ�4@{Oh8/�!?Y����@ލ&�C�ٿ�i��@��ΰ�4@{Oh8/�!?Y����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@�&�XS�ٿT%HW8��@�Ђ�:4@@�-ڋ�!?P8����@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@���bw�ٿ�$"�?��@AK럘)4@���U�!?G�f��*�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@�9���ٿ�&ɇv_�@v��*�3@�J�P�!?�i�ټP�@���Yg�ٿX�� 	�@*y#�3@ۭ$�w�!?�ޞ�5u�@ob$;l�ٿ8�5���@�]��3@Q��1Ӑ!?Q6���A�@ob$;l�ٿ8�5���@�]��3@Q��1Ӑ!?Q6���A�@ob$;l�ٿ8�5���@�]��3@Q��1Ӑ!?Q6���A�@���k*�ٿW�ױ|�@H�k��3@��L��!?Br���@���k*�ٿW�ױ|�@H�k��3@��L��!?Br���@���k*�ٿW�ױ|�@H�k��3@��L��!?Br���@���k*�ٿW�ױ|�@H�k��3@��L��!?Br���@���k*�ٿW�ױ|�@H�k��3@��L��!?Br���@B�հ��ٿ����7�@i�Eς'4@�<���!?���;�@A�q�ٿ6������@�X��~�3@zj�!?d'�H�$�@A�q�ٿ6������@�X��~�3@zj�!?d'�H�$�@A�q�ٿ6������@�X��~�3@zj�!?d'�H�$�@��O>[�ٿz����7�@�G!�O�3@f]�o�!?~P�:�@����~�ٿ������@1�{�3@[&f��!?,��f؟�@����~�ٿ������@1�{�3@[&f��!?,��f؟�@����~�ٿ������@1�{�3@[&f��!?,��f؟�@������ٿ��~���@>��M�4@����ɐ!?�0�Z �@������ٿ��~���@>��M�4@����ɐ!?�0�Z �@������ٿ��~���@>��M�4@����ɐ!?�0�Z �@�&���ٿC�B�:�@e4�~�R4@���^�!?QK@��@�&���ٿC�B�:�@e4�~�R4@���^�!?QK@��@�&���ٿC�B�:�@e4�~�R4@���^�!?QK@��@�-!��ٿ�˺�.1�@�R�'�3@̤Xw�!?^wi��Ε@���ٿfش��@n��F�3@������!?~)�8��@���ٿfش��@n��F�3@������!?~)�8��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@?N$�"�ٿ�ϕn��@A�v��4@o�]��!?�,��|��@���>�ٿA�[]��@}믳�&4@;;�+�!?�őՕ@���>�ٿA�[]��@}믳�&4@;;�+�!?�őՕ@���>�ٿA�[]��@}믳�&4@;;�+�!?�őՕ@���>�ٿA�[]��@}믳�&4@;;�+�!?�őՕ@�L��ٿ�ר�$�@����'4@%#̶X�!?d����@�L��ٿ�ר�$�@����'4@%#̶X�!?d����@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@����n�ٿ��X�Y��@��L@�34@��jn�!?~mCV9ԕ@f	e�ٿ�85�@Q�2��3@dB}�!?��rڇ��@f	e�ٿ�85�@Q�2��3@dB}�!?��rڇ��@f	e�ٿ�85�@Q�2��3@dB}�!?��rڇ��@f	e�ٿ�85�@Q�2��3@dB}�!?��rڇ��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@8��kE�ٿ|�yXu	�@�q���3@P^�S�!?��Z�5��@�;T~Y�ٿ��!����@y�i��3@$P��k�!?������@��ổٿ'�b���@Vv��-	4@��'5z�!?��B�Bb�@��ổٿ'�b���@Vv��-	4@��'5z�!?��B�Bb�@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@���c�ٿ=l^�>L�@(�|�54@ڼ�`��!?��d>� �@F��M�ٿ<!%�@_[�+�3@��9��!?�7�ߖ�@F��M�ٿ<!%�@_[�+�3@��9��!?�7�ߖ�@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@���Ƽ�ٿ�w���A�@��6��4@H_`��!?�rPNbΕ@Z���ٿ	6����@=�g*��3@��!�!?��{I9��@Z���ٿ	6����@=�g*��3@��!�!?��{I9��@�EQ&i�ٿ������@�����3@'v�J�!?لV�n��@�t<~�ٿ�_ɚ��@�����3@�>��8�!?C����@�t<~�ٿ�_ɚ��@�����3@�>��8�!?C����@�t<~�ٿ�_ɚ��@�����3@�>��8�!?C����@��k՛ٿ�ݻ���@��E�3@-��8�!?�듟nӕ@��k՛ٿ�ݻ���@��E�3@-��8�!?�듟nӕ@��k՛ٿ�ݻ���@��E�3@-��8�!?�듟nӕ@��k՛ٿ�ݻ���@��E�3@-��8�!?�듟nӕ@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@��Xq�ٿ
"�.=��@R
q��3@/���!?ȋl��t�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@2�Y��ٿ�2Ef��@	�2|4@�d4�!?��ʩ�,�@BT����ٿ`���d2�@x���s"4@(O���!?����~�@@��-��ٿ�y���@��	��84@FP�]��!?�%��`��@@��-��ٿ�y���@��	��84@FP�]��!?�%��`��@5�ީ�ٿ�p�(��@��)1R4@d`��ϐ!?߁n��@�w�Q�ٿ?#6�M��@���v�G4@7��/i�!?P��(�@�w�Q�ٿ?#6�M��@���v�G4@7��/i�!?P��(�@�w�Q�ٿ?#6�M��@���v�G4@7��/i�!?P��(�@�w�Q�ٿ?#6�M��@���v�G4@7��/i�!?P��(�@�w�Q�ٿ?#6�M��@���v�G4@7��/i�!?P��(�@�	`g2�ٿ����*�@���E4@�W�<@�!?N�	���@�	`g2�ٿ����*�@���E4@�W�<@�!?N�	���@�	`g2�ٿ����*�@���E4@�W�<@�!?N�	���@�	`g2�ٿ����*�@���E4@�W�<@�!?N�	���@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@���,��ٿ;ǹbx��@�=�X�\4@E|V��!?�/��Е@�̗禖ٿ��ɦ�}�@t3�,M4@�<Ho%�!?1x*�Y��@�̗禖ٿ��ɦ�}�@t3�,M4@�<Ho%�!?1x*�Y��@��e>�ٿU�Z�}��@�f�q4@��ٷ��!?�5�b�z�@�يm�ٿ������@~/�C4@����!?<nxgs�@�يm�ٿ������@~/�C4@����!?<nxgs�@�يm�ٿ������@~/�C4@����!?<nxgs�@�يm�ٿ������@~/�C4@����!?<nxgs�@Wʭ�	�ٿ���y��@j�a��4@4b�2�!?Q��ZV�@Wʭ�	�ٿ���y��@j�a��4@4b�2�!?Q��ZV�@ܷe!4�ٿ@��h�\�@��"^p4@Qg-�!?��f�#ȕ@ܷe!4�ٿ@��h�\�@��"^p4@Qg-�!?��f�#ȕ@^�Q��ٿoKv��S�@�.��r%4@�5(v�!?�Oe.��@�����ٿ�����@7���� 4@�h� �!?��}%V�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@�	�w��ٿU^�<ž�@0�/�4@I����!?�A��2�@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@rW�i�ٿ���k���@o�j���3@Z{���!?��uU���@�C��j�ٿ��T�@o��3~4@_	b�!?Q{>kJ��@08��r�ٿ��ؑ���@BԊcc4@�ӋQM�!?�4J��@08��r�ٿ��ؑ���@BԊcc4@�ӋQM�!?�4J��@08��r�ٿ��ؑ���@BԊcc4@�ӋQM�!?�4J��@08��r�ٿ��ؑ���@BԊcc4@�ӋQM�!?�4J��@i�GG��ٿ�Ĭ6���@DNK��4@�� �<�!?� �4��@�7�Y��ٿ@V򁑁�@�!+U/4@R�Ż}�!?'���@
��}|�ٿ��>���@z@�}4@"p�td�!?2���+�@
��}|�ٿ��>���@z@�}4@"p�td�!?2���+�@
��}|�ٿ��>���@z@�}4@"p�td�!?2���+�@
��}|�ٿ��>���@z@�}4@"p�td�!?2���+�@
��}|�ٿ��>���@z@�}4@"p�td�!?2���+�@��,X)�ٿ������@3|�v�4@���홐!?�e�)F�@g|`Җٿ��(��t�@Λ��04@��x��!?y z|��@g|`Җٿ��(��t�@Λ��04@��x��!?y z|��@g|`Җٿ��(��t�@Λ��04@��x��!?y z|��@gw�X��ٿ287�� �@��|�@4@wt�,�!?�r��@gw�X��ٿ287�� �@��|�@4@wt�,�!?�r��@gw�X��ٿ287�� �@��|�@4@wt�,�!?�r��@wʲ�$�ٿ�twH�@�^n�B4@��!i�!?����>�@wʲ�$�ٿ�twH�@�^n�B4@��!i�!?����>�@wʲ�$�ٿ�twH�@�^n�B4@��!i�!?����>�@m��ٿph%��p�@:dQ��<4@��܋�!?簙&S�@m��ٿph%��p�@:dQ��<4@��܋�!?簙&S�@m��ٿph%��p�@:dQ��<4@��܋�!?簙&S�@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@ve�ٿ�Q��1�@'���X4@Xj2q�!?^0���@B�	�ݚٿ���1�@���54@�����!?����.1�@B�	�ݚٿ���1�@���54@�����!?����.1�@B�	�ݚٿ���1�@���54@�����!?����.1�@B�	�ݚٿ���1�@���54@�����!?����.1�@B�	�ݚٿ���1�@���54@�����!?����.1�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@m&𖟚ٿae;�@o;�T�#4@���	��!?F��H�@�rE�ɡٿ�lo�R�@��n}�3@
Xͯ�!?��XZ���@�rE�ɡٿ�lo�R�@��n}�3@
Xͯ�!?��XZ���@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@��G�W�ٿI�����@;Vo1��3@���C��!?[�����@�yJ)<�ٿ�W�	S�@{@u�14@�8��3�!?o�����@lş}�ٿS�.D��@�ȱ�h�3@(���M�!?#Ha�u�@lş}�ٿS�.D��@�ȱ�h�3@(���M�!?#Ha�u�@lş}�ٿS�.D��@�ȱ�h�3@(���M�!?#Ha�u�@lş}�ٿS�.D��@�ȱ�h�3@(���M�!?#Ha�u�@��Ɂ2�ٿnP��7��@�?ڇ14@ M�]d�!?	�, LÕ@��Ɂ2�ٿnP��7��@�?ڇ14@ M�]d�!?	�, LÕ@��Ɂ2�ٿnP��7��@�?ڇ14@ M�]d�!?	�, LÕ@��Ɂ2�ٿnP��7��@�?ڇ14@ M�]d�!?	�, LÕ@��Ɂ2�ٿnP��7��@�?ڇ14@ M�]d�!?	�, LÕ@o]۠ٿ�ի�_�@ui1��3@�{��r�!?��6�Õ@o]۠ٿ�ի�_�@ui1��3@�{��r�!?��6�Õ@�q�A�ٿ�|SQ�W�@���'"4@GK:Uc�!?��s�@�I~���ٿК����@�k�'4@� �tk�!?��WO<�@�I~���ٿК����@�k�'4@� �tk�!?��WO<�@�I~���ٿК����@�k�'4@� �tk�!?��WO<�@�I~���ٿК����@�k�'4@� �tk�!?��WO<�@it��=�ٿ�'ڼ=��@�����3@C�7�!?X�%�愕@it��=�ٿ�'ڼ=��@�����3@C�7�!?X�%�愕@h�d�d�ٿw豀���@�l����3@�~�.�!?�ʭ����@���d�ٿ�2�����@%����3@(��!?��gWԕ@�b��ٿ|����@}��qq4@��ؚ_�!?�s�c��@�b��ٿ|����@}��qq4@��ؚ_�!?�s�c��@8�*f�ٿC�EN��@��u�S,4@�~j�n�!?��hXE�@8�*f�ٿC�EN��@��u�S,4@�~j�n�!?��hXE�@8�*f�ٿC�EN��@��u�S,4@�~j�n�!?��hXE�@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@�.˖�ٿ�N��@��?#4@� �
5�!?�4����@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@A�{-�ٿ�uy8��@<�5$4@��\�!?�C9���@�z�H�ٿI|����@J:��*4@� ~qW�!?	O%(�@�z�H�ٿI|����@J:��*4@� ~qW�!?	O%(�@�z�H�ٿI|����@J:��*4@� ~qW�!?	O%(�@�z�H�ٿI|����@J:��*4@� ~qW�!?	O%(�@�z�H�ٿI|����@J:��*4@� ~qW�!?	O%(�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@P휏�ٿ�k6{�@;�T;4@)��iP�!?3 #�@��ٿE�̪�@]Z?�34@Ȑ0vO�!?�ҙor�@b�R�ٞٿ`����b�@n<�&4@�W�	�!?�EtW��@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@7�@�ٿ���&N�@6�	4@�d�0[�!?HV�}_�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@�3�w�ٿs&����@r2���4@����u�!?���s�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@Lu��ٿ��©n�@��f3�*4@��Cא�!?����S�@tI�2�ٿC�_����@��Op�=4@2ן�*�!?z Jڕ@tI�2�ٿC�_����@��Op�=4@2ן�*�!?z Jڕ@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@���ȷ�ٿFBG簞�@�]�::4@�k��H�!?���o���@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@�r�k�ٿI}�?+�@�����(4@$���h�!?&�}R�
�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@����ٿV�x�ܨ�@�^14@r×�+�!?�"j��*�@0ނP�ٿ�)�O.�@��ELD+4@~�2��!?;�]��K�@0ނP�ٿ�)�O.�@��ELD+4@~�2��!?;�]��K�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@��w	�ٿ���O��@G����4@
�Q�!?vje�@�\4�T�ٿ�v8��=�@i
?D4@�M2�'�!?>�V����@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@&Z�#�ٿ�e�N�@C��R[4@�2HK�!?[�Ӝ�>�@h3�s��ٿ��5���@�y,.�3@9�Ƙ/�!?�f��Å�@h3�s��ٿ��5���@�y,.�3@9�Ƙ/�!?�f��Å�@h3�s��ٿ��5���@�y,.�3@9�Ƙ/�!?�f��Å�@h3�s��ٿ��5���@�y,.�3@9�Ƙ/�!?�f��Å�@h3�s��ٿ��5���@�y,.�3@9�Ƙ/�!?�f��Å�@�%��ٿ�T*����@0�V��3@�@��z�!?g��g�@�%��ٿ�T*����@0�V��3@�@��z�!?g��g�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@݈��(�ٿ�6�kb��@܋(Q�3@�%���!?�0�1C�@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@0�V\�ٿ��p��Z�@)(3HB�3@��AҚ�!?�,��@>�e��ٿTX�����@��gP� 4@�^��!?s�d�"��@>�e��ٿTX�����@��gP� 4@�^��!?s�d�"��@���r	�ٿ��Y��@"�;L��3@��MӐ!?[	��飕@���r	�ٿ��Y��@"�;L��3@��MӐ!?[	��飕@z�*:]�ٿ�lZ�	�@)���3@j]�Z��!?���e��@z�*:]�ٿ�lZ�	�@)���3@j]�Z��!?���e��@�̀��ٿ�T�MS��@��oy44@��Ǹ��!?e{�)Io�@�̀��ٿ�T�MS��@��oy44@��Ǹ��!?e{�)Io�@N�`�ٿ`�8��@=mm��3@�x���!?��0>��@�ݴ�1�ٿ#�s��@)R����3@sۼ�~�!?#��*�@�ݴ�1�ٿ#�s��@)R����3@sۼ�~�!?#��*�@�ݴ�1�ٿ#�s��@)R����3@sۼ�~�!?#��*�@�ݴ�1�ٿ#�s��@)R����3@sۼ�~�!?#��*�@�ݴ�1�ٿ#�s��@)R����3@sۼ�~�!?#��*�@H���ٿ۟����@����4@w���[�!?��zy4��@��L���ٿ���p��@���B4@̡��5�!?Y^�hЕ@��L���ٿ���p��@���B4@̡��5�!?Y^�hЕ@?^�Z�ٿ������@���'4@h�����!?QCø֕@��)Ad�ٿ~ю	f�@5A�T�"4@b���!?�-D���@��)Ad�ٿ~ю	f�@5A�T�"4@b���!?�-D���@��)Ad�ٿ~ю	f�@5A�T�"4@b���!?�-D���@��)Ad�ٿ~ю	f�@5A�T�"4@b���!?�-D���@���ʘٿ�ԑ�@G�&W04@�j�x0�!?�*�.��@���ʘٿ�ԑ�@G�&W04@�j�x0�!?�*�.��@���ʘٿ�ԑ�@G�&W04@�j�x0�!?�*�.��@���ʘٿ�ԑ�@G�&W04@�j�x0�!?�*�.��@���ʘٿ�ԑ�@G�&W04@�j�x0�!?�*�.��@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@7ݝޠ�ٿ�#Ǚ,��@�����"4@�z���!?S��9�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@L��c�ٿQU�p�e�@���6F4@O)�ki�!?p���5q�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@�x�a��ٿ*B��x�@��d7�+4@� �F�!?�����3�@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@!�E�ٿj!T=���@:��n)4@����/�!?p`�j͕@��l��ٿi���6��@{�祥-4@A�r���!?�?��͕@��l��ٿi���6��@{�祥-4@A�r���!?�?��͕@��l��ٿi���6��@{�祥-4@A�r���!?�?��͕@��l��ٿi���6��@{�祥-4@A�r���!?�?��͕@��l��ٿi���6��@{�祥-4@A�r���!?�?��͕@Ҧ���ٿ�	�|V��@�A�64@g9H6g�!?FQѕ@|�P��ٿ���>��@Zq��-4@7T�� �!?�Ґcm�@|�P��ٿ���>��@Zq��-4@7T�� �!?�Ґcm�@|�P��ٿ���>��@Zq��-4@7T�� �!?�Ґcm�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@5d�H�ٿ	؋���@�]��D%4@heo>�!?:QN��c�@�-}�T�ٿ���k�@-Dk��4@�t�-�!?�x`;�@�-}�T�ٿ���k�@-Dk��4@�t�-�!?�x`;�@�-}�T�ٿ���k�@-Dk��4@�t�-�!?�x`;�@�-}�T�ٿ���k�@-Dk��4@�t�-�!?�x`;�@�-}�T�ٿ���k�@-Dk��4@�t�-�!?�x`;�@�8M|�ٿ��T'��@�����14@t�M�!?���bh�@�8M|�ٿ��T'��@�����14@t�M�!?���bh�@�8M|�ٿ��T'��@�����14@t�M�!?���bh�@�8M|�ٿ��T'��@�����14@t�M�!?���bh�@�[���ٿ8d�Xz�@��;P�84@|�1�8�!?���zy�@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@��5��ٿJ�y/:�@-Z2)�N4@=N��+�!?޻P#i��@v���$�ٿf`�(��@�vw_�64@�̝Pe�!?����R��@v���$�ٿf`�(��@�vw_�64@�̝Pe�!?����R��@v���$�ٿf`�(��@�vw_�64@�̝Pe�!?����R��@v���$�ٿf`�(��@�vw_�64@�̝Pe�!?����R��@v���$�ٿf`�(��@�vw_�64@�̝Pe�!?����R��@�CEs��ٿ��!����@�0���4@؟ZWS�!?���!�@�CEs��ٿ��!����@�0���4@؟ZWS�!?���!�@�CEs��ٿ��!����@�0���4@؟ZWS�!?���!�@�CEs��ٿ��!����@�0���4@؟ZWS�!?���!�@ýxw�ٿ���2��@Ȉ�x�:4@��E)�!?��s"�%�@ýxw�ٿ���2��@Ȉ�x�:4@��E)�!?��s"�%�@ýxw�ٿ���2��@Ȉ�x�:4@��E)�!?��s"�%�@ýxw�ٿ���2��@Ȉ�x�:4@��E)�!?��s"�%�@ ��淨ٿ����@c�!R04@��vX�!?�
�u��@ ��淨ٿ����@c�!R04@��vX�!?�
�u��@ ��淨ٿ����@c�!R04@��vX�!?�
�u��@��(E��ٿ`]�!Օ�@ppEe^4@�Ⱥ�W�!?;��꾜�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@.R�Ӛٿ�t�K�@ra�4@��C�O�!?�L�,A{�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�H$ �ٿ��)E*��@��Y4@}zk�?�!?wۂ��v�@�
�=i�ٿO"'%��@砌��4@;0����!?�m�G�@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�0Y��ٿ�9tΒ+�@kj�4@0���ُ!?�Z�ƕ@�d�F��ٿ���@�I�@�~���
4@��s�!?n0�AU�@�d�F��ٿ���@�I�@�~���
4@��s�!?n0�AU�@��/S�ٿ��� ͠�@@�H�g4@���6�!?�$+ےݕ@��/S�ٿ��� ͠�@@�H�g4@���6�!?�$+ےݕ@��/S�ٿ��� ͠�@@�H�g4@���6�!?�$+ےݕ@��/S�ٿ��� ͠�@@�H�g4@���6�!?�$+ےݕ@��/S�ٿ��� ͠�@@�H�g4@���6�!?�$+ےݕ@n�l���ٿq��:�@��%s4@��p�!?�����@n�l���ٿq��:�@��%s4@��p�!?�����@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@�U>�c�ٿAH_d�E�@���"4@�`2�!?���>F �@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@���ٿ�����@mdL��4@���["�!?���m�ϕ@N^�ũ�ٿ0{�d�@�@��ڢ1�3@4x�\�!?MB
<�Е@N^�ũ�ٿ0{�d�@�@��ڢ1�3@4x�\�!?MB
<�Е@N^�ũ�ٿ0{�d�@�@��ڢ1�3@4x�\�!?MB
<�Е@N^�ũ�ٿ0{�d�@�@��ڢ1�3@4x�\�!?MB
<�Е@�c����ٿ���5��@�wq4@�X�R�!?���{Kt�@�c����ٿ���5��@�wq4@�X�R�!?���{Kt�@Ƃ�V&�ٿ��Q`�@΀g��%4@��`��!?��:���@Ƃ�V&�ٿ��Q`�@΀g��%4@��`��!?��:���@Ƃ�V&�ٿ��Q`�@΀g��%4@��`��!?��:���@o��ߗٿ���b���@��g�.$4@F�!`��!?z$Л.��@Բf�A�ٿ|�����@y$"D�/4@f�R�)�!?-Ie�ƕ@Բf�A�ٿ|�����@y$"D�/4@f�R�)�!?-Ie�ƕ@Բf�A�ٿ|�����@y$"D�/4@f�R�)�!?-Ie�ƕ@� r~x�ٿDqe�@���#4@G��	%�!?_��7:��@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@Y���O�ٿDIqĸ��@D�r�""4@��!?f��s �@��l��ٿ�T�g�@T�^ �3@{��!?��J�I�@��l��ٿ�T�g�@T�^ �3@{��!?��J�I�@vl#�J�ٿP�'��@D���W�3@[����!?�Z0u�r�@vl#�J�ٿP�'��@D���W�3@[����!?�Z0u�r�@vl#�J�ٿP�'��@D���W�3@[����!?�Z0u�r�@ܭ]T�ٿU��;��@��4@�2j�!?oaM�(�@�"HU��ٿN,%�A�@���u4@������!?�n��ⴖ@�"HU��ٿN,%�A�@���u4@������!?�n��ⴖ@i�6��ٿ�l-��B�@��-�;4@'3��!?�Q�4@i�6��ٿ�l-��B�@��-�;4@'3��!?�Q�4@i�6��ٿ�l-��B�@��-�;4@'3��!?�Q�4@�v$�,�ٿ�gR�,�@�L_o�4@�t	���!?��^��Z�@�v$�,�ٿ�gR�,�@�L_o�4@�t	���!?��^��Z�@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@�Mٛٿ���Q��@�j{-�4@F��O�!?�?��ȕ@Tc����ٿ�Q:RG��@�/\4@�`Nd�!?�8�Ȣ��@Tc����ٿ�Q:RG��@�/\4@�`Nd�!?�8�Ȣ��@Tc����ٿ�Q:RG��@�/\4@�`Nd�!?�8�Ȣ��@N�AK�ٿ�_�ڃ=�@�ɹ�S,4@����!?�ǻ�D��@N�AK�ٿ�_�ڃ=�@�ɹ�S,4@����!?�ǻ�D��@N�AK�ٿ�_�ڃ=�@�ɹ�S,4@����!?�ǻ�D��@C��q֠ٿq�?��#�@�o��(04@�נ�L�!?�v�E���@C��q֠ٿq�?��#�@�o��(04@�נ�L�!?�v�E���@����ٿ������@���4@K(voe�!?O!�̕@����ٿ������@���4@K(voe�!?O!�̕@����ٿ������@���4@K(voe�!?O!�̕@����ٿ������@���4@K(voe�!?O!�̕@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@MH̆ٝٿ��1���@W��"4@�=^�c�!?��ɺ�@M��!8�ٿ6\����@�{Z~�>4@6D�/��!?b�P��@4tt���ٿ��8K�@)w���N4@���W��!?|�:A�@4tt���ٿ��8K�@)w���N4@���W��!?|�:A�@4tt���ٿ��8K�@)w���N4@���W��!?|�:A�@8�b{ӝٿ$[�t��@�"�e4@��5_�!?������@���2l�ٿ�XYo	��@���J4@/04;�!?��{Zl�@���2l�ٿ�XYo	��@���J4@/04;�!?��{Zl�@�Z��-�ٿ���e#��@Eρx�.4@��?�!?Fq�D�@�Z��-�ٿ���e#��@Eρx�.4@��?�!?Fq�D�@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@�@CJ�ٿ�bs��@�i��A'4@O�3/_�!?5�.���@-K��[�ٿQ����@悇��4@�cn@?�!?2���@-K��[�ٿQ����@悇��4@�cn@?�!?2���@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@cQ���ٿ5~2���@3t��`4@�mG�:�!?��&&w��@xϖT؜ٿ�.����@��m�!+4@#��Mf�!?0Yh��@�΄��ٿ�c���C�@�g��>"4@!�<���!?m_Ѫ��@�΄��ٿ�c���C�@�g��>"4@!�<���!?m_Ѫ��@�΄��ٿ�c���C�@�g��>"4@!�<���!?m_Ѫ��@�΄��ٿ�c���C�@�g��>"4@!�<���!?m_Ѫ��@|KTzp�ٿY�$��@�F�K�'4@V��)M�!?r9�kR��@�(��F�ٿ8�J�@���2(4@D���A�!?�I�ccv�@�(��F�ٿ8�J�@���2(4@D���A�!?�I�ccv�@N���ٿ���*��@�<I?M4@�8u��!?��G�:�@N���ٿ���*��@�<I?M4@�8u��!?��G�:�@N���ٿ���*��@�<I?M4@�8u��!?��G�:�@N���ٿ���*��@�<I?M4@�8u��!?��G�:�@N���ٿ���*��@�<I?M4@�8u��!?��G�:�@��d�ٿ�.�3Zr�@_:��;P4@+cx�!?i����@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@w�P-T�ٿ�/��i��@s��
-4@��D�j�!?v���ו@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@��0��ٿ�?�Vi�@�O<�K4@Y挅s�!?_+�����@6o�ٿ�>G[�@��B4@�Jk�@�!?J�(�G�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@X�
�ڝٿ�hj4c�@^tf��84@����a�!?*��&#E�@���ٿޅ���@΄^�44@լ�}�!?�B��ە@���ٿޅ���@΄^�44@լ�}�!?�B��ە@ԧMF�ٿF�z��J�@��~��E4@��Hk�!?�"�+�@ԧMF�ٿF�z��J�@��~��E4@��Hk�!?�"�+�@ԧMF�ٿF�z��J�@��~��E4@��Hk�!?�"�+�@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@}eGǜٿX��@�wf�D4@�NH�d�!?꟤���@�+��)�ٿ�{�)bi�@v%��4@t���!?ڌ��J˕@�+��)�ٿ�{�)bi�@v%��4@t���!?ڌ��J˕@�+��)�ٿ�{�)bi�@v%��4@t���!?ڌ��J˕@�2vO�ٿN��Y��@�SQWq!4@�P�ԕ�!?��u�P�@�2vO�ٿN��Y��@�SQWq!4@�P�ԕ�!?��u�P�@�2vO�ٿN��Y��@�SQWq!4@�P�ԕ�!?��u�P�@��8�ٿs<p���@��r�4@Lq	��!?�r��F�@��8�ٿs<p���@��r�4@Lq	��!?�r��F�@��8�ٿs<p���@��r�4@Lq	��!?�r��F�@��8�ٿs<p���@��r�4@Lq	��!?�r��F�@a���ٿp2�^S�@�Ƃ��3@�s�c��!?WNQ��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@	S�G��ٿ@�j�8�@�Ҫj)�3@e�G͐!?M�	�R��@��� ��ٿ'���5�@	c���3@��^S��!?P��6��@��� ��ٿ'���5�@	c���3@��^S��!?P��6��@��� ��ٿ'���5�@	c���3@��^S��!?P��6��@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@Gc�/�ٿ(|�o�@1x��4@�-�析!?���.�@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@ju!H�ٿſ;���@�t��- 4@�2��!?�xp�֕@�zc2�ٿ��2�a�@�W/7�=4@��&?�!?%y�F2��@�zc2�ٿ��2�a�@�W/7�=4@��&?�!?%y�F2��@��hx��ٿ������@�#;�(]4@��Ke�!?0����@�ğLͤٿ_��!}��@yY�c�D4@��Fkߐ!?f�|XK
�@�ğLͤٿ_��!}��@yY�c�D4@��Fkߐ!?f�|XK
�@�w~ k�ٿ�&�tm��@Ɠ�7	4@��!?����@�w~ k�ٿ�&�tm��@Ɠ�7	4@��!?����@�w~ k�ٿ�&�tm��@Ɠ�7	4@��!?����@�w~ k�ٿ�&�tm��@Ɠ�7	4@��!?����@�1�)�ٿ�5�Ox��@�$MP�3@5@.�ܐ!?*T�����@(�q��ٿu��\݀�@�~7�3@2�t�ڐ!?@�Σ��@(�q��ٿu��\݀�@�~7�3@2�t�ڐ!?@�Σ��@(�q��ٿu��\݀�@�~7�3@2�t�ڐ!?@�Σ��@(�q��ٿu��\݀�@�~7�3@2�t�ڐ!?@�Σ��@��9�
�ٿ��yV��@(J��3@0�ݡ��!?g�!g�ŕ@�1$���ٿ�r�;���@>}n�g�3@�����!?f�j��@�P��Ֆٿ�,v�NF�@$�����3@hZ����!?"E.}�ߕ@�P��Ֆٿ�,v�NF�@$�����3@hZ����!?"E.}�ߕ@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@#�Nλ�ٿ?�6V+��@���}�3@a"�+��!?k�v��N�@'��Y��ٿBd�d�@8[w��3@��ђ_�!?#O�}�,�@'��Y��ٿBd�d�@8[w��3@��ђ_�!?#O�}�,�@R�8���ٿƷ�d��@�d����3@��%w�!?����^d�@H-o+r�ٿn�+Ɉ�@�����3@��63�!?���V�@H-o+r�ٿn�+Ɉ�@�����3@��63�!?���V�@H-o+r�ٿn�+Ɉ�@�����3@��63�!?���V�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@3<܀ �ٿmz�,�@�֍��3@$��:�!?��#�Я�@	��'��ٿ� �XB�@����M4@ҕQ �!?*�
�Y�@	��'��ٿ� �XB�@����M4@ҕQ �!?*�
�Y�@X��8КٿN��r�@��PfZd4@P��#�!?�X���@X��8КٿN��r�@��PfZd4@P��#�!?�X���@�G ��ٿ�o�>��@�|;��<4@�����!?����Fe�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@'�Aŷ�ٿzɹE�Z�@f���4@��q��!?�0p�@~SwJ�ٿ�"l��@ë��h4@�
G�א!?�-�5�@~SwJ�ٿ�"l��@ë��h4@�
G�א!?�-�5�@~SwJ�ٿ�"l��@ë��h4@�
G�א!?�-�5�@~SwJ�ٿ�"l��@ë��h4@�
G�א!?�-�5�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@14'T��ٿܴ�ܧ�@��R�4@ZR���!?��|�@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@y�졜ٿ@��a�@��Y|4@v��c&�!?[3�Z]��@�Ұ?Ŗٿ��@�:�@�d��&4@�ڙ�`�!?�AC�dE�@�Ұ?Ŗٿ��@�:�@�d��&4@�ڙ�`�!?�AC�dE�@��>��ٿ�d�!$��@���3b�3@��74�!?f	nK#�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@d@kژٿ��~��5�@Վ���4@����G�!?c��B�@o��F�ٿB�O�&��@.$BH
4@_����!?�df�!�@o��F�ٿB�O�&��@.$BH
4@_����!?�df�!�@o��F�ٿB�O�&��@.$BH
4@_����!?�df�!�@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@7Lvs�ٿ�IR]���@Ȝ/
�:4@3���l�!?E���@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@��](�ٿ��[���@�晣.�3@��Cw�!?��ǚq�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@v�˒]�ٿ@d��U�@2�����3@�u{F�!?�͙'8�@V�k�ٿ��0��V�@0v@*�3@Q�����!?���t(�@ߡ;	?�ٿЎ��n��@ֿ>S�3@��o�J�!?������@ߡ;	?�ٿЎ��n��@ֿ>S�3@��o�J�!?������@�M��ٿ	���(�@gC����3@�[a5�!?��D���@�M��ٿ	���(�@gC����3@�[a5�!?��D���@�M��ٿ	���(�@gC����3@�[a5�!?��D���@�n��{�ٿ�'���@��\%j�3@���P�!??�כ]�@�n��{�ٿ�'���@��\%j�3@���P�!??�כ]�@�n��{�ٿ�'���@��\%j�3@���P�!??�כ]�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�V�ES�ٿ}nD�e�@~�X�4@��rKU�!?�ǥ��=�@�b���ٿ�H[Kq��@��?��4@������!?����@M@�C�ٿҢ���@�f��W4@jԥ�z�!?R}�k��@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@�2,ƙٿ5�4�@�{�'4@[�)@}�!?�)���Е@C���ٿ-����@K�ي4@���"��!?y�H��@C���ٿ-����@K�ي4@���"��!?y�H��@C���ٿ-����@K�ي4@���"��!?y�H��@C���ٿ-����@K�ي4@���"��!?y�H��@C���ٿ-����@K�ي4@���"��!?y�H��@w�|h��ٿ=B.҆��@�4C�=44@.���{�!?���pbٕ@w�|h��ٿ=B.҆��@�4C�=44@.���{�!?���pbٕ@w�|h��ٿ=B.҆��@�4C�=44@.���{�!?���pbٕ@w�|h��ٿ=B.҆��@�4C�=44@.���{�!?���pbٕ@�&�Üٿ�	��Ҳ�@��m�O4@���hg�!?�޽x��@�&�Üٿ�	��Ҳ�@��m�O4@���hg�!?�޽x��@h�m�ٿ�'���@&�$�84@����$�!?��'~� �@h�m�ٿ�'���@&�$�84@����$�!?��'~� �@{�2�֢ٿW��Qy��@{�t4�44@wø�|�!?������@{�2�֢ٿW��Qy��@{�t4�44@wø�|�!?������@{�2�֢ٿW��Qy��@{�t4�44@wø�|�!?������@�_-�ٿy��n��@5�����3@��V�!?	��89�@�_-�ٿy��n��@5�����3@��V�!?	��89�@�_-�ٿy��n��@5�����3@��V�!?	��89�@�_-�ٿy��n��@5�����3@��V�!?	��89�@�_-�ٿy��n��@5�����3@��V�!?	��89�@�_-�ٿy��n��@5�����3@��V�!?	��89�@��#T�ٿ/z3t�@���0W�3@z�h.�!?.�&뺓�@��#T�ٿ/z3t�@���0W�3@z�h.�!?.�&뺓�@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@^��ٿ��<]�x�@9�[���3@)�*�!?H�y8p��@*CӠ��ٿ��=�0�@@�{�V�3@��6le�!?[��@*CӠ��ٿ��=�0�@@�{�V�3@��6le�!?[��@*CӠ��ٿ��=�0�@@�{�V�3@��6le�!?[��@*CӠ��ٿ��=�0�@@�{�V�3@��6le�!?[��@�Rn�ٿ�/�z�@��߆�3@{얼�!?�[.�7ݕ@�Rn�ٿ�/�z�@��߆�3@{얼�!?�[.�7ݕ@�Rn�ٿ�/�z�@��߆�3@{얼�!?�[.�7ݕ@�Rn�ٿ�/�z�@��߆�3@{얼�!?�[.�7ݕ@�N���ٿ�	$�R��@
�lC>4@8����!?h�	"@�N���ٿ�	$�R��@
�lC>4@8����!?h�	"@O�Q�K�ٿ+�-:a�@�&w{�O4@e�#�Y�!?����y�@O�Q�K�ٿ+�-:a�@�&w{�O4@e�#�Y�!?����y�@O�Q�K�ٿ+�-:a�@�&w{�O4@e�#�Y�!?����y�@:�vy��ٿ���YA��@����e4@F�����!?�l%A���@:�vy��ٿ���YA��@����e4@F�����!?�l%A���@:�vy��ٿ���YA��@����e4@F�����!?�l%A���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@�>,_r�ٿ�$n%�r�@��[t4@bS�ٛ�!?��l���@E&� T�ٿ�o��|z�@S֙�R4@Y�9<��!?�*���@�c�qќٿa�K8<�@�|��&4@,cɐ!?��y�p�@�c�qќٿa�K8<�@�|��&4@,cɐ!?��y�p�@�c�qќٿa�K8<�@�|��&4@,cɐ!?��y�p�@���Oטٿ�b7p�@k����3@QN����!?�Β)~e�@���Oטٿ�b7p�@k����3@QN����!?�Β)~e�@���Oטٿ�b7p�@k����3@QN����!?�Β)~e�@���Oטٿ�b7p�@k����3@QN����!?�Β)~e�@\,���ٿ"��(���@�J��3@6=��|�!?5"���=�@\,���ٿ"��(���@�J��3@6=��|�!?5"���=�@\,���ٿ"��(���@�J��3@6=��|�!?5"���=�@�o7rA�ٿ2������@F=����3@0�+��!?W��	��@U��	��ٿ/L��3�@�5 V�3@~'��y�!?��e��@U��	��ٿ/L��3�@�5 V�3@~'��y�!?��e��@�b�b��ٿ�f���@�f�_�3@~�j�̐!?T�� �ɕ@�b�b��ٿ�f���@�f�_�3@~�j�̐!?T�� �ɕ@�b�b��ٿ�f���@�f�_�3@~�j�̐!?T�� �ɕ@�b�b��ٿ�f���@�f�_�3@~�j�̐!?T�� �ɕ@�b�b��ٿ�f���@�f�_�3@~�j�̐!?T�� �ɕ@eWp�ٿ@�����@D�EDA4@
~ �H�!?���Һƕ@eWp�ٿ@�����@D�EDA4@
~ �H�!?���Һƕ@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@�Ȋ�ٿ��e�1Q�@Y6a+�.4@���(m�!?S����@j�$I�ٿʟR�	�@�-���"4@T�	p�!?D\-Xﳕ@j�$I�ٿʟR�	�@�-���"4@T�	p�!?D\-Xﳕ@���.�ٿq��j� �@ےa��3@G�X:�!?���N��@���.�ٿq��j� �@ےa��3@G�X:�!?���N��@���.�ٿq��j� �@ےa��3@G�X:�!?���N��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@Ţ<��ٿh��ʗ@�@�Ԛ�9�3@�yKM �!?�$�%��@�1
�/�ٿc0����@���5�3@�V��F�!?^�0f���@�1
�/�ٿc0����@���5�3@�V��F�!?^�0f���@�1
�/�ٿc0����@���5�3@�V��F�!?^�0f���@�0�j�ٿ2�n��@�����3@
P=�m�!?�����̕@�0�j�ٿ2�n��@�����3@
P=�m�!?�����̕@�0�j�ٿ2�n��@�����3@
P=�m�!?�����̕@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@B���ٿc�{�A�@�X��V4@��0G�!?D%nW,��@AU��ٿ*"�]�@}dz�N4@�'P�*�!?xY��[�@AU��ٿ*"�]�@}dz�N4@�'P�*�!?xY��[�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@�=�	�ٿ��7��^�@���g�b4@$�-��!?��h�b�@v˙:�ٿT��=
��@��]C4@|k�|y�!?+�v#	�@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@d�g��ٿ�(!'}b�@On�E$4@�i��e�!?�du�r��@VDU	G�ٿ����@���`yB4@�n�<�!?շ�NYܕ@b�E��ٿ	��??�@�G���P4@J�>e�!?�@\2]��@���z�ٿ^u�ϧ��@�2��:4@�(��!?�fԄ��@���z�ٿ^u�ϧ��@�2��:4@�(��!?�fԄ��@���z�ٿ^u�ϧ��@�2��:4@�(��!?�fԄ��@Ɇ��ܚٿɭE���@��0�:=4@��CD��!?�Ξ��@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@���ٿ��ٓ���@n]���F4@J����!?������@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@lQF�ؖٿ1��4�@x�rO4@9iWH��!?R8?�杕@IǸv�ٿ��-�G��@�C?t�14@jC�I��!?���cÕ@IǸv�ٿ��-�G��@�C?t�14@jC�I��!?���cÕ@IǸv�ٿ��-�G��@�C?t�14@jC�I��!?���cÕ@IǸv�ٿ��-�G��@�C?t�14@jC�I��!?���cÕ@IǸv�ٿ��-�G��@�C?t�14@jC�I��!?���cÕ@.���ٿvpPz�@x�3�4@�ː2o�!?,�?���@.���ٿvpPz�@x�3�4@�ː2o�!?,�?���@.���ٿvpPz�@x�3�4@�ː2o�!?,�?���@.���ٿvpPz�@x�3�4@�ː2o�!?,�?���@=Q��r�ٿoۓ`���@3��4@�=vE��!?fG�����@=Q��r�ٿoۓ`���@3��4@�=vE��!?fG�����@=Q��r�ٿoۓ`���@3��4@�=vE��!?fG�����@�f��q�ٿ��8�z�@�W�"94@Q���s�!?:-�q�@�f��q�ٿ��8�z�@�W�"94@Q���s�!?:-�q�@(�s>�ٿ=��o�@��5��64@R+�ډ�!?F^�Ow�@(�s>�ٿ=��o�@��5��64@R+�ډ�!?F^�Ow�@(�s>�ٿ=��o�@��5��64@R+�ډ�!?F^�Ow�@<��M��ٿ:!=��@�q�7	4@����j�!?�nH7d�@<��M��ٿ:!=��@�q�7	4@����j�!?�nH7d�@<��M��ٿ:!=��@�q�7	4@����j�!?�nH7d�@<��M��ٿ:!=��@�q�7	4@����j�!?�nH7d�@+}3��ٿ�N;���@�
��3@�q�Ap�!?���NaD�@*1|��ٿx�S�8�@"3���4@��7Z�!?�j9c�F�@*1|��ٿx�S�8�@"3���4@��7Z�!?�j9c�F�@*1|��ٿx�S�8�@"3���4@��7Z�!?�j9c�F�@�Q���ٿ߂]S<"�@c��w
#4@��,�!?��B�L�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@ы���ٿ�%x��S�@C���m4@S��+�!?g��dcF�@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@7x�^��ٿV���=��@uc4h;4@�?K�!?Dd����@.=���ٿB�?�2��@S���GK4@eJ"�,�!?�� ՂJ�@.=���ٿB�?�2��@S���GK4@eJ"�,�!?�� ՂJ�@��Z��ٿ�?ڗ��@�j��4@|
��/�!?u7���\�@��Z��ٿ�?ڗ��@�j��4@|
��/�!?u7���\�@��Z��ٿ�?ڗ��@�j��4@|
��/�!?u7���\�@��Z��ٿ�?ڗ��@�j��4@|
��/�!?u7���\�@��Z��ٿ�?ڗ��@�j��4@|
��/�!?u7���\�@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@ ��w��ٿ��i�)�@1mYJ4@�vEX�!?�������@(�����ٿ�����(�@��!��	4@a� �&�!?S�j�ޕ@,�����ٿ��ځ&��@�e�c�	4@�ra��!?��� ͕@,�����ٿ��ځ&��@�e�c�	4@�ra��!?��� ͕@,�����ٿ��ځ&��@�e�c�	4@�ra��!?��� ͕@,�����ٿ��ځ&��@�e�c�	4@�ra��!?��� ͕@��'�ۤٿ�U�����@�3�74@��I�!?�D0~m�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�:�>N�ٿ\ed� ��@���3@�2��@�!?�4��8D�@�v��Ӝٿ����?�@�Ř^n34@��a`>�!?����)�@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@K1N95�ٿ1��>5��@�"�:�3@�l�D��!?%9f�- �@�c�p7�ٿ�$#���@�LnRn�3@a8;mV�!?<��~ƕ@�c�p7�ٿ�$#���@�LnRn�3@a8;mV�!?<��~ƕ@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@K����ٿpV]d���@��C1�3@�G}9�!?��$9���@C���ٿ�n9�7�@�"�Z+4@&�[cE�!?x�����@C���ٿ�n9�7�@�"�Z+4@&�[cE�!?x�����@C���ٿ�n9�7�@�"�Z+4@&�[cE�!?x�����@C���ٿ�n9�7�@�"�Z+4@&�[cE�!?x�����@C���ٿ�n9�7�@�"�Z+4@&�[cE�!?x�����@LU�9�ٿą��s��@�8�p�4@�9gѐ!?,�̲�ŕ@LU�9�ٿą��s��@�8�p�4@�9gѐ!?,�̲�ŕ@LU�9�ٿą��s��@�8�p�4@�9gѐ!?,�̲�ŕ@LU�9�ٿą��s��@�8�p�4@�9gѐ!?,�̲�ŕ@T\驚ٿC���,��@��.>�04@��靐!?,�/M< �@U���ٿj@�~(�@�'94@f&�w��!?���-�Ε@U���ٿj@�~(�@�'94@f&�w��!?���-�Ε@U���ٿj@�~(�@�'94@f&�w��!?���-�Ε@U���ٿj@�~(�@�'94@f&�w��!?���-�Ε@P�%�ٿ���=��@�TP�94@Q%�ŵ�!?&a��&%�@S�6�ٿR�~��@�*�S 4@r�l���!?% ֩M8�@S�6�ٿR�~��@�*�S 4@r�l���!?% ֩M8�@S�6�ٿR�~��@�*�S 4@r�l���!?% ֩M8�@�N�2'�ٿ�Gf1�@�_���3@*�1��!?L�Ġ1 �@i���ٿ��Jo���@C��.p�3@W,�V�!?�w���)�@���ٿ4.��^��@��q764@�q]fZ�!?
����S�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�Nx�J�ٿ���+���@��z��(4@��T���!?��{2'�@�c7S�ٿċ��R��@ı,��4@Vl�Qv�!?=��˛ȕ@X�����ٿ�C��%-�@Rn�
�3@Ϳ�uX�!?1�[p��@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@��(q�ٿY��]��@������3@�-�u�!?�g1u�y�@W���ٿ���D��@k�n�4@�S���!?�}1��@W���ٿ���D��@k�n�4@�S���!?�}1��@W���ٿ���D��@k�n�4@�S���!?�}1��@31�v�ٿ���Z��@;0�'fQ4@�k��}�!?�!`NU֕@31�v�ٿ���Z��@;0�'fQ4@�k��}�!?�!`NU֕@�C����ٿ��F�@,`�0.u4@��=��!?u6L(���@�C����ٿ��F�@,`�0.u4@��=��!?u6L(���@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@�\''�ٿ>o	���@�қ�Yl4@�(𰢐!?���C|��@��Upe�ٿD����@�Nè"�3@HKV��!?.[]`�@��Upe�ٿD����@�Nè"�3@HKV��!?.[]`�@��Upe�ٿD����@�Nè"�3@HKV��!?.[]`�@��Upe�ٿD����@�Nè"�3@HKV��!?.[]`�@��Upe�ٿD����@�Nè"�3@HKV��!?.[]`�@}�Y���ٿK�<��@1Ԕw�	4@�n�34�!?T�Ǳ��@��=�ŚٿWw��?�@\h��o 4@���!?�0�r�@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@]��塛ٿ&�JF��@� _�84@���`�!?��b�Nޕ@ז��N�ٿp�&2/�@�K-�L4@���x�!?I�~�N�@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@�Lۛ��ٿ�Ϻ?Z/�@��?�54@��!.�!?n�`����@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@Z�K3��ٿ�����=�@p����44@CJ}�)�!?��A#���@]n��ٿ/<���k�@�˶��C4@Q��kb�!?j��"c�@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@u�����ٿj�wX�@/P��4@Z[���!?�j�A}��@C��\�ٿ��\ڔ�@���\�F4@�8�:�!?d���tؕ@C��\�ٿ��\ڔ�@���\�F4@�8�:�!?d���tؕ@C��\�ٿ��\ڔ�@���\�F4@�8�:�!?d���tؕ@B�k� �ٿ(���-�@����4@��=�N�!?9�*�:Ε@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@D����ٿ�`�xI&�@$��;��3@�A�A�!?؝̧�=�@/���Ԛٿ�}��m��@��=�3�3@ĵ���!?�)(P�@/���Ԛٿ�}��m��@��=�3�3@ĵ���!?�)(P�@.�ٿb�Wo��@���u�3@��>7�!?׫/�d�@.�ٿb�Wo��@���u�3@��>7�!?׫/�d�@�G���ٿ�=�m�@N�Q4@'l	B1�!?�W��R�@�G���ٿ�=�m�@N�Q4@'l	B1�!?�W��R�@�G���ٿ�=�m�@N�Q4@'l	B1�!?�W��R�@�G���ٿ�=�m�@N�Q4@'l	B1�!?�W��R�@��m�ٿ.zӢI&�@��5��4@H9>�G�!?2�*0ҕ@��m�ٿ.zӢI&�@��5��4@H9>�G�!?2�*0ҕ@ƣ�c�ٿ`A�&���@�{�]��3@��M*q�!?��Ս��@ƣ�c�ٿ`A�&���@�{�]��3@��M*q�!?��Ս��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@�9]ޛٿ�&�-�@s<��3@�Wxi_�!?|z]\��@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@��� �ٿ��u#��@�Y�
"4@}0��#�!?6?�H5N�@�����ٿ�}Tm��@���>4@��i�!?IG�pGٕ@�����ٿ�}Tm��@���>4@��i�!?IG�pGٕ@�����ٿ�}Tm��@���>4@��i�!?IG�pGٕ@�����ٿ�}Tm��@���>4@��i�!?IG�pGٕ@����V�ٿb�(�@��,�x�3@FŐ�!?m�{�]ӕ@����V�ٿb�(�@��,�x�3@FŐ�!?m�{�]ӕ@��{�>�ٿ8:>M���@�ݹ�3@�֡j�!?�m!�H�@9�ޛ&�ٿ�bkjo�@#9�@4�3@�
�mj�!?��H(p�@9�ޛ&�ٿ�bkjo�@#9�@4�3@�
�mj�!?��H(p�@9�ޛ&�ٿ�bkjo�@#9�@4�3@�
�mj�!?��H(p�@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@�(Ş�ٿO��7��@���34@;�q���!?�������@[&5K�ٿ�ve ֋�@ �[�4@��Y]�!?%B'秕@[&5K�ٿ�ve ֋�@ �[�4@��Y]�!?%B'秕@[&5K�ٿ�ve ֋�@ �[�4@��Y]�!?%B'秕@�O1��ٿ��o5k�@x�l2�4@L� �n�!??�Z�P��@�O1��ٿ��o5k�@x�l2�4@L� �n�!??�Z�P��@�O1��ٿ��o5k�@x�l2�4@L� �n�!??�Z�P��@E�[�n�ٿ�����m�@h�;�/4@��H���!?�g�ą��@E�[�n�ٿ�����m�@h�;�/4@��H���!?�g�ą��@�[���ٿBzCZ��@�*S��D4@i2� ��!?2�����@w��Ht�ٿf�n�;�@�ݒ04@'����!?�y�z��@w��Ht�ٿf�n�;�@�ݒ04@'����!?�y�z��@�2
���ٿӳU�@�Ǯ�@4@h�a�u�!?���`!�@�2
���ٿӳU�@�Ǯ�@4@h�a�u�!?���`!�@�2
���ٿӳU�@�Ǯ�@4@h�a�u�!?���`!�@��v˙ٿ��3�@Q5�E4@�Z?�i�!?U�����@��W⸛ٿ�@y�'��@��?<44@Tn�y&�!?T��fc�@��W⸛ٿ�@y�'��@��?<44@Tn�y&�!?T��fc�@���9�ٿ���O���@���:4@���խ�!?3c��@	��P�ٿL`�H�@���m�24@q&�Ƃ�!?�c��
�@	��P�ٿL`�H�@���m�24@q&�Ƃ�!?�c��
�@	��P�ٿL`�H�@���m�24@q&�Ƃ�!?�c��
�@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@��/ڡٿO���V��@:KѾ�K4@#h��M�!?J��0ʕ@�'�_ƥٿI2�5���@��ʾ�4@F��YF�!?�Q�]�!�@�'�_ƥٿI2�5���@��ʾ�4@F��YF�!?�Q�]�!�@�'�_ƥٿI2�5���@��ʾ�4@F��YF�!?�Q�]�!�@z�nd�ٿH�N����@x ��4@�Ǭ~��!?_J��l�@L�&�k�ٿ3?�V�@G�H�d:4@�GF�2�!?/�u���@L�&�k�ٿ3?�V�@G�H�d:4@�GF�2�!?/�u���@L�&�k�ٿ3?�V�@G�H�d:4@�GF�2�!?/�u���@����)�ٿ �z{l[�@a��9O+4@W7��!?�f�x�@����)�ٿ �z{l[�@a��9O+4@W7��!?�f�x�@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@a����ٿb�k��@����'4@�����!?�$����@�X�ٿ4�.�@Q�@�L2�3@`�mz�!?����̕@�X�ٿ4�.�@Q�@�L2�3@`�mz�!?����̕@�X�ٿ4�.�@Q�@�L2�3@`�mz�!?����̕@�X�ٿ4�.�@Q�@�L2�3@`�mz�!?����̕@N�ꓡٿ=9��q��@���Uf�3@߭1g�!?���� �@��)�ٿ��+��@)�����3@4�E��!?��VD	�@��)�ٿ��+��@)�����3@4�E��!?��VD	�@��)�ٿ��+��@)�����3@4�E��!?��VD	�@��)�ٿ��+��@)�����3@4�E��!?��VD	�@��)�ٿ��+��@)�����3@4�E��!?��VD	�@�e��[�ٿ���%$�@<G��54@dӍ�!?�Csx��@�e��[�ٿ���%$�@<G��54@dӍ�!?�Csx��@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@_��?�ٿ�*�uD$�@�<54@�%��d�!?B�����@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@I�>��ٿ� �3��@���
4@Se{�~�!?�%�漕@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@��f:�ٿ)�b���@�Z$4@���扐!?HAY��@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@ȃ� U�ٿ�'~a�!�@��*K%4@�>�bT�!?N�{~Е@+�I��ٿ|h�k��@n�n�"4@:r)�!?��2U�@+�I��ٿ|h�k��@n�n�"4@:r)�!?��2U�@+�I��ٿ|h�k��@n�n�"4@:r)�!?��2U�@C%b��ٿ`���5��@Z���@�3@�쵕G�!?hCMf�J�@���l%�ٿ��+ێn�@�?�Z~$4@�>/8�!?�݌)@G�@O����ٿ��"���@}1e�n�3@�� 9�!?���Ze��@O����ٿ��"���@}1e�n�3@�� 9�!?���Ze��@O����ٿ��"���@}1e�n�3@�� 9�!?���Ze��@C?�F�ٿG#KP�@�(�g�3@l*�&t�!?��0��@C?�F�ٿG#KP�@�(�g�3@l*�&t�!?��0��@��I���ٿ|i��`�@�U����3@w�L�!?���wU�@�ꑻ��ٿ����[��@�u���3@�!�e7�!?>P��)a�@�ꑻ��ٿ����[��@�u���3@�!�e7�!?>P��)a�@�ꑻ��ٿ����[��@�u���3@�!�e7�!?>P��)a�@�G�ٿw����@V�jF�3@\?��!?"�����@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@������ٿfﶇ.�@���q?�3@��/�X�!?��ܔ�@���?��ٿoq�@���@��c	�4@Ʈ��)�!?�U��^��@���?��ٿoq�@���@��c	�4@Ʈ��)�!?�U��^��@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@:�8�|�ٿ��L�}^�@G��TA$4@�&?9�!?*�:�[�@z #���ٿs��gB��@�E��4@�8Bw�!?���@z #���ٿs��gB��@�E��4@�8Bw�!?���@z #���ٿs��gB��@�E��4@�8Bw�!?���@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�O�-��ٿ�c��d�@��G4@R{:_�!?��~�H�@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@�{�3�ٿF��g7�@��q�4@C����!?P2;~H��@O��q�ٿ���X���@�T�l4@(�o��!?C^�J��@y8�?�ٿ�U0+���@ �vy4@�"�`��!?}�WW��@y8�?�ٿ�U0+���@ �vy4@�"�`��!?}�WW��@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@L�@|�ٿ��ru�@Op��F4@��[�!?�'�b�ԕ@�S��ٿ��!~�@2c�G4@I��拐!?��!F���@�S��ٿ��!~�@2c�G4@I��拐!?��!F���@�S��ٿ��!~�@2c�G4@I��拐!?��!F���@�ls'_�ٿ�Q�c��@�gշ�74@�v��Ɛ!?��x���@�ls'_�ٿ�Q�c��@�gշ�74@�v��Ɛ!?��x���@�ls'_�ٿ�Q�c��@�gշ�74@�v��Ɛ!?��x���@�ls'_�ٿ�Q�c��@�gշ�74@�v��Ɛ!?��x���@G�����ٿA��%���@��p܅^4@�"W��!?c~` k�@v�A��ٿ{>�K�@ b�24@Pw�y
�!?�M߮�9�@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@kqj�טٿ6p,�%�@R�|=�%4@��fs�!?P��#��@`a\��ٿ09��jI�@iMh*C4@�~�m��!?��Qdb>�@`a\��ٿ09��jI�@iMh*C4@�~�m��!?��Qdb>�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@���*�ٿϝv�:�@�]j<�4@)`!��!?�>	J�@�U�|�ٿ��\E��@��o���3@���8��!?�q���O�@�U�|�ٿ��\E��@��o���3@���8��!?�q���O�@�U�|�ٿ��\E��@��o���3@���8��!?�q���O�@�U�|�ٿ��\E��@��o���3@���8��!?�q���O�@�U�|�ٿ��\E��@��o���3@���8��!?�q���O�@������ٿM�,1��@t@w���3@��փ�!?�1I��W�@������ٿM�,1��@t@w���3@��փ�!?�1I��W�@������ٿM�,1��@t@w���3@��փ�!?�1I��W�@�>o�	�ٿ�ڲMz�@m���4@�;r�O�!?��r�s�@�>o�	�ٿ�ڲMz�@m���4@�;r�O�!?��r�s�@�>o�	�ٿ�ڲMz�@m���4@�;r�O�!?��r�s�@�>o�	�ٿ�ڲMz�@m���4@�;r�O�!?��r�s�@��_��ٿx���I-�@�v ��4@D��5��!?�%~���@�?��ٿ2�
���@���T�3@L_�܂�!?	�ɭו@��y�ٿ�J@���@�Q���4@~-���!?(�@Pѕ@��y�ٿ�J@���@�Q���4@~-���!?(�@Pѕ@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@�	Ue�ٿ�X�URD�@�r�&&4@�S�v�!?�E(�<c�@��C$c�ٿq�]#e�@��G�4@� _s��!?Y���N��@��C$c�ٿq�]#e�@��G�4@� _s��!?Y���N��@�����ٿ��M�%�@�r64@x�+(��!?�z��H�@�����ٿ��M�%�@�r64@x�+(��!?�z��H�@�����ٿ��M�%�@�r64@x�+(��!?�z��H�@Z<;��ٿ�Q/Z��@]_\�64@�>O�h�!?����q�@Z<;��ٿ�Q/Z��@]_\�64@�>O�h�!?����q�@���x�ٿ6�R��@���3@�(��!?�d�ϕ@;6T�[�ٿ��f���@ ����3@Z�,��!?� c�Vѕ@M���t�ٿN�1��2�@���#��3@�Xx���!?��;���@M���t�ٿN�1��2�@���#��3@�Xx���!?��;���@M���t�ٿN�1��2�@���#��3@�Xx���!?��;���@M���t�ٿN�1��2�@���#��3@�Xx���!?��;���@N�|,�ٿ��5Opr�@��C)4@���B�!?��A����@N�|,�ٿ��5Opr�@��C)4@���B�!?��A����@N�|,�ٿ��5Opr�@��C)4@���B�!?��A����@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@�gbݜٿz��+��@�d{F�4@�im�m�!?{��f[�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@䐼�Κٿk�/|�@�q6��_4@P?�Ah�!?�B'�,�@��񎺗ٿ��M��@����4@�ZdT�!?�����@��񎺗ٿ��M��@����4@�ZdT�!?�����@��񎺗ٿ��M��@����4@�ZdT�!?�����@�����ٿ����x��@?@�U�$4@8�(�!?���*:F�@��g�%�ٿ@��j&�@	��M4@�u����!?��5or�@��g�%�ٿ@��j&�@	��M4@�u����!?��5or�@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@:��EZ�ٿ�I����@�[Mq4@6G����!?���._Ε@Aİҩ�ٿ��ʂ)�@��P�<4@O*�-�!?�>�7쫕@�hLB�ٿ�����@6����3@<�@*�!?�Z��h�@�hLB�ٿ�����@6����3@<�@*�!?�Z��h�@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@aS�͜ٿ�&O ��@��3KB4@�+��W�!?� -{ѕ@���4�ٿR��t��@�;�bG^4@1��8�!?��k��s�@���4�ٿR��t��@�;�bG^4@1��8�!?��k��s�@�}W�V�ٿW퉰��@^�ƪbN4@�~q2�!?w�P�H"�@��@zF�ٿT��(�@�}�P�?4@���(��!?r�#���@��@zF�ٿT��(�@�}�P�?4@���(��!?r�#���@��@zF�ٿT��(�@�}�P�?4@���(��!?r�#���@��@zF�ٿT��(�@�}�P�?4@���(��!?r�#���@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@�Ėy>�ٿ*�.��6�@�#eT9>4@��U�U�!?n���Q�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@lul��ٿPG�p��@ F��F4@��R��!?�h�h�c�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@��⏕�ٿxKǋ�@��x�G4@��o)h�!?�s�_�@v��c�ٿY�É.�@��GXic4@�	�=��!?;z��U�@v��c�ٿY�É.�@��GXic4@�	�=��!?;z��U�@7L6ed�ٿ:�t�#��@�?���C4@����ǐ!?��!���@7L6ed�ٿ:�t�#��@�?���C4@����ǐ!?��!���@7L6ed�ٿ:�t�#��@�?���C4@����ǐ!?��!���@7L6ed�ٿ:�t�#��@�?���C4@����ǐ!?��!���@7L6ed�ٿ:�t�#��@�?���C4@����ǐ!?��!���@�e�n�ٿ�!}���@�^DD4@9��C��!?er���@}�@%�ٿ���N� �@4/��3@�k�>N�!?������@}�@%�ٿ���N� �@4/��3@�k�>N�!?������@QAo|��ٿ��B���@ߨ���	4@��-s�!?wKNj�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@!���q�ٿ dzI6�@ۈ�4�,4@�����!?�v���,�@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@FGY�&�ٿ�9�r�@�.m?�3@�,�g�!?R.�ו@d�tǞٿ��XD0X�@v���4@��o�!?�?AT��@8)�՝ٿPGm��h�@�Z�y� 4@X��I�!?Е�!�B�@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@���ٕ�ٿ��=�}��@��S�;4@��6�!?NmD�jƕ@	3
���ٿ��38�@��)�UQ4@S�=�!?wc���@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@�)Թ�ٿ�V��@��Z�3@A܈:c�!?Q�T3��@	�	��ٿ��:C�@�E�4@SЧ-;�!?)��'(�@	�	��ٿ��:C�@�E�4@SЧ-;�!?)��'(�@"��%ۜٿ~���i�@�!@��4@��i1�!?_?s/v$�@��)*Ϛٿz�K����@��	a�4@��ܶR�!?��C�E�@���i�ٿ��l��@���#4@�4[/��!?�i��^�@���i�ٿ��l��@���#4@�4[/��!?�i��^�@���i�ٿ��l��@���#4@�4[/��!?�i��^�@���i�ٿ��l��@���#4@�4[/��!?�i��^�@o�'�ٿz�J�?��@�Cj[4@�,����!?��[�m�@o�'�ٿz�J�?��@�Cj[4@�,����!?��[�m�@o�'�ٿz�J�?��@�Cj[4@�,����!?��[�m�@o�'�ٿz�J�?��@�Cj[4@�,����!?��[�m�@o�'�ٿz�J�?��@�Cj[4@�,����!?��[�m�@�a|x�ٿEGlPV�@�<�5�G4@,3��!?sY��V�@�"�b�ٿ�,�B��@c���44@���Jې!?���^_;�@�"�b�ٿ�,�B��@c���44@���Jې!?���^_;�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@��i�؝ٿ>��  �@��)4@��b���!?9�QjQh�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@~��$�ٿ7Z��!�@C3V��4@�5�֢�!?���O�@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@���f�ٿ��`����@S'���4@� ���!?t�Z�ʕ@��=_�ٿ5.�����@nq�l'4@�7P�3�!?a��:[�@��=_�ٿ5.�����@nq�l'4@�7P�3�!?a��:[�@��v˞ٿM�7��U�@�@���3@*�L�5�!?��Bt*�@��v˞ٿM�7��U�@�@���3@*�L�5�!?��Bt*�@��v˞ٿM�7��U�@�@���3@*�L�5�!?��Bt*�@��v˞ٿM�7��U�@�@���3@*�L�5�!?��Bt*�@U;*���ٿ�J�ȼ��@����[�3@��w�|�!?=0��*�@����ޘٿ,�@���@e�gĵ�3@�FL��!?� ��ĕ@����ޘٿ,�@���@e�gĵ�3@�FL��!?� ��ĕ@����Փٿ�� 5��@����3@�o!�r�!?jK��=�@����Փٿ�� 5��@����3@�o!�r�!?jK��=�@����Փٿ�� 5��@����3@�o!�r�!?jK��=�@���Śٿc��~��@A\e�3@1h �!?K��L�@���Śٿc��~��@A\e�3@1h �!?K��L�@��e�ٿ�����@��\��3@�r�fO�!?~_���@��e�ٿ�����@��\��3@�r�fO�!?~_���@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@��I��ٿX�<���@6x�{��3@SU-���!?�\y-��@�*b�o�ٿ�HB���@�.D"B4@���|�!?e�IF�{�@�*b�o�ٿ�HB���@�.D"B4@���|�!?e�IF�{�@�*b�o�ٿ�HB���@�.D"B4@���|�!?e�IF�{�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@(AS��ٿzWM�8�@���RU4@�N_(�!?s(�a\�@g����ٿ��P6@u�@����#4@�*d���!?�~h�E�@g����ٿ��P6@u�@����#4@�*d���!?�~h�E�@g����ٿ��P6@u�@����#4@�*d���!?�~h�E�@��)o��ٿ�����@��nk��3@�m���!?.Z��ޕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�'��ٿ�4�	&+�@��ԥ?�3@DS�i�!?'
��ϕ@�W ��ٿ8��Z��@a��F�4@�� �:�!?~M����@�W ��ٿ8��Z��@a��F�4@�� �:�!?~M����@�W ��ٿ8��Z��@a��F�4@�� �:�!?~M����@�W ��ٿ8��Z��@a��F�4@�� �:�!?~M����@�X�ԝٿ�_ t�@#��3@���s�!?������@�X�ԝٿ�_ t�@#��3@���s�!?������@�X�ԝٿ�_ t�@#��3@���s�!?������@�X�ԝٿ�_ t�@#��3@���s�!?������@�X�ԝٿ�_ t�@#��3@���s�!?������@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@s=���ٿ�/���s�@h���3@�ƽe��!?=&�oT9�@[+�=w�ٿA
���u�@�*�XH�3@��$��!?����)�@[+�=w�ٿA
���u�@�*�XH�3@��$��!?����)�@[+�=w�ٿA
���u�@�*�XH�3@��$��!?����)�@[+�=w�ٿA
���u�@�*�XH�3@��$��!?����)�@�?�N�ٿQ���@�;��<4@�tg�!?�"Bӽ��@�?�N�ٿQ���@�;��<4@�tg�!?�"Bӽ��@�~�"��ٿ<F�?��@��34@	k��!?��)0b�@�~�"��ٿ<F�?��@��34@	k��!?��)0b�@�~�"��ٿ<F�?��@��34@	k��!?��)0b�@�~�"��ٿ<F�?��@��34@	k��!?��)0b�@�F�Ϫ�ٿov��?�@��X��G4@�2���!?)�BIb�@�F�Ϫ�ٿov��?�@��X��G4@�2���!?)�BIb�@�F�Ϫ�ٿov��?�@��X��G4@�2���!?)�BIb�@�F�Ϫ�ٿov��?�@��X��G4@�2���!?)�BIb�@5q��=�ٿ�/"�@M��h��3@�$}=r�!?�����@5q��=�ٿ�/"�@M��h��3@�$}=r�!?�����@5q��=�ٿ�/"�@M��h��3@�$}=r�!?�����@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@i�tT��ٿ�w�.A�@MLM�3@��o�!?��l��@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@@f��k�ٿa�:[r��@3���
�3@0N�(��!?�=�	?�@���~��ٿ/��d���@���O��3@��m@G�!?mv@���~��ٿ/��d���@���O��3@��m@G�!?mv@�J�;��ٿ�CMos�@����4@w���!?��Ɯ��@� q�@�ٿ�߭k��@�{�GQ4@SK�92�!?���zݣ�@� q�@�ٿ�߭k��@�{�GQ4@SK�92�!?���zݣ�@� q�@�ٿ�߭k��@�{�GQ4@SK�92�!?���zݣ�@���ٿ�S��+�@�H
�3@���k�!?��ܔ�W�@���ٿ�S��+�@�H
�3@���k�!?��ܔ�W�@���ٿ�S��+�@�H
�3@���k�!?��ܔ�W�@���ٿ�S��+�@�H
�3@���k�!?��ܔ�W�@�_��y�ٿ]4Ot��@��Xp)4@"2���!?���;�@��k�&�ٿ�T�k��@i�g�=14@�B+@��!?4���]��@��k�&�ٿ�T�k��@i�g�=14@�B+@��!?4���]��@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@42 .�ٿ/[�:(~�@%G���c4@�5�:k�!?�z�>�@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��uaМٿ�U����@�ʄh�3@�+9N�!?l0(Xԕ@��F�0�ٿHْ��{�@��Η�:4@H��W�!?y�0��@+����ٿS?�(���@��)�=4@P%S2��!?\����@+����ٿS?�(���@��)�=4@P%S2��!?\����@+����ٿS?�(���@��)�=4@P%S2��!?\����@+����ٿS?�(���@��)�=4@P%S2��!?\����@+����ٿS?�(���@��)�=4@P%S2��!?\����@+����ٿS?�(���@��)�=4@P%S2��!?\����@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�~�&�ٿ��*��@]J���&4@˗+���!? �9��Е@�p^�m�ٿ�Y���@�H=�$4@��.-t�!?�4�:;�@�p^�m�ٿ�Y���@�H=�$4@��.-t�!?�4�:;�@�p^�m�ٿ�Y���@�H=�$4@��.-t�!?�4�:;�@�p^�m�ٿ�Y���@�H=�$4@��.-t�!?�4�:;�@�p^�m�ٿ�Y���@�H=�$4@��.-t�!?�4�:;�@TB's�ٿ�)��x�@%���AJ4@��EUY�!?���#Q��@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@J��ii�ٿS�m���@��<]w4@s,�H:�!?S������@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@�G!�1�ٿ���"���@V��24@N$R�Q�!?理ԕ@9<Mu"�ٿ�����@+�t�D4@���f2�!?�ތ3Õ@i�\,�ٿjq�����@�� L@4@���h^�!?�&�`��@i�\,�ٿjq�����@�� L@4@���h^�!?�&�`��@�wV�b�ٿ���L�Y�@���,R4@��X�!?�����@�wV�b�ٿ���L�Y�@���,R4@��X�!?�����@�wV�b�ٿ���L�Y�@���,R4@��X�!?�����@�wV�b�ٿ���L�Y�@���,R4@��X�!?�����@���WՙٿV�w�|7�@�<�h�64@o�)��!?X`�ԯ�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@]���ܟٿ&���N��@R�]sY4@cvH�V�!?n�?=lL�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@-��<�ٿ����F��@���\4@����Ð!?$}��c2�@u�i�H�ٿeTl�C��@�� Oz4@J  �p�!?�6�j���@u�i�H�ٿeTl�C��@�� Oz4@J  �p�!?�6�j���@u�i�H�ٿeTl�C��@�� Oz4@J  �p�!?�6�j���@�E����ٿ�O�VJ�@�->e14@��r�!?$ ��3�@�E����ٿ�O�VJ�@�->e14@��r�!?$ ��3�@�E����ٿ�O�VJ�@�->e14@��r�!?$ ��3�@�E����ٿ�O�VJ�@�->e14@��r�!?$ ��3�@�E����ٿ�O�VJ�@�->e14@��r�!?$ ��3�@1\4'�ٿJ��>�^�@a�J�4@fM�s��!?�6�}���@����ٿu\�x�<�@�3�"�3@�!E�-�!?�+�m��@����ٿu\�x�<�@�3�"�3@�!E�-�!?�+�m��@����ٿu\�x�<�@�3�"�3@�!E�-�!?�+�m��@����ٿu\�x�<�@�3�"�3@�!E�-�!?�+�m��@����ٿu\�x�<�@�3�"�3@�!E�-�!?�+�m��@��-��ٿ��c�	8�@s!�I	�3@�{�`d�!?V)l5_��@��-��ٿ��c�	8�@s!�I	�3@�{�`d�!?V)l5_��@��-��ٿ��c�	8�@s!�I	�3@�{�`d�!?V)l5_��@�T��j�ٿ�d�g�@ۦ�^74@N�N��!?2��}�@�T��j�ٿ�d�g�@ۦ�^74@N�N��!?2��}�@�T��j�ٿ�d�g�@ۦ�^74@N�N��!?2��}�@�T��j�ٿ�d�g�@ۦ�^74@N�N��!?2��}�@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@�4��c�ٿ�^�"���@��Y���3@r�~v�!?�< ��@5���ٿ�p�@���C�4@�����!?s��lt�@5���ٿ�p�@���C�4@�����!?s��lt�@5���ٿ�p�@���C�4@�����!?s��lt�@�ͦ�"�ٿJ܄	��@�KU��3@����a�!?#\�`5�@�ͦ�"�ٿJ܄	��@�KU��3@����a�!?#\�`5�@5�O��ٿ'�j����@;㘧�4@��y,�!?��6iR\�@5�O��ٿ'�j����@;㘧�4@��y,�!?��6iR\�@5�O��ٿ'�j����@;㘧�4@��y,�!?��6iR\�@��@ �ٿ)��/��@U��8�3@�{��>�!?�:�Hv͕@��@ �ٿ)��/��@U��8�3@�{��>�!?�:�Hv͕@��@ �ٿ)��/��@U��8�3@�{��>�!?�:�Hv͕@��@ �ٿ)��/��@U��8�3@�{��>�!?�:�Hv͕@��@ �ٿ)��/��@U��8�3@�{��>�!?�:�Hv͕@�ٿ��/��z�@�L�14@�G� �!?�I��ؕ@�ٿ��/��z�@�L�14@�G� �!?�I��ؕ@�ٿ��/��z�@�L�14@�G� �!?�I��ؕ@�@	�1�ٿ�:q�@o6��4@�3�֏!?�"`�tݕ@�����ٿ82���*�@�P)�(�3@҅����!?��*aϕ@],����ٿ�a��Y�@e���C�3@89+2�!?�H?;��@],����ٿ�a��Y�@e���C�3@89+2�!?�H?;��@],����ٿ�a��Y�@e���C�3@89+2�!?�H?;��@],����ٿ�a��Y�@e���C�3@89+2�!?�H?;��@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@9r론ٿ;(m~9��@qT�Q*4@;�q�*�!?,b��̕@�Oz�t�ٿ�^�Ce��@'J�E84@U���,�!?ԭvq�4�@�Oz�t�ٿ�^�Ce��@'J�E84@U���,�!?ԭvq�4�@�Oz�t�ٿ�^�Ce��@'J�E84@U���,�!?ԭvq�4�@�Oz�t�ٿ�^�Ce��@'J�E84@U���,�!?ԭvq�4�@�Oz�t�ٿ�^�Ce��@'J�E84@U���,�!?ԭvq�4�@�o���ٿ�8��@���&)4@2J�R�!?��BꟋ�@�o���ٿ�8��@���&)4@2J�R�!?��BꟋ�@�o���ٿ�8��@���&)4@2J�R�!?��BꟋ�@s(ٽ�ٿ�y�*%��@��BT4@�kf.�!?���ŏ�@s(ٽ�ٿ�y�*%��@��BT4@�kf.�!?���ŏ�@�����ٿ��p�\��@t'��~4@:�Gt��!?�CQB%�@�Z�n�ٿI��g��@k�:o�X4@[�2o�!?��7����@�Z�n�ٿI��g��@k�:o�X4@[�2o�!?��7����@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@��;�^�ٿ�@����@���d�3@��~f�!?�
�5*��@a�ԕ}�ٿ��	���@��ؖ�3@����!?� Չs�@�Uǧ�ٿ��pu�E�@�����3@��^�!?�t_�p�@�Uǧ�ٿ��pu�E�@�����3@��^�!?�t_�p�@&�V���ٿ�P?*�@�h�\A4@~�d���!?�NL��@&�V���ٿ�P?*�@�h�\A4@~�d���!?�NL��@&�V���ٿ�P?*�@�h�\A4@~�d���!?�NL��@�� �ٿd+�\��@0�V"Vp4@)�|�|�!?o&�'�	�@�� �ٿd+�\��@0�V"Vp4@)�|�|�!?o&�'�	�@�� �ٿd+�\��@0�V"Vp4@)�|�|�!?o&�'�	�@�� �ٿd+�\��@0�V"Vp4@)�|�|�!?o&�'�	�@��h�ٿL�9"�@/f�4p4@�4 ڃ�!?!/��a�@��h�ٿL�9"�@/f�4p4@�4 ڃ�!?!/��a�@��h�ٿL�9"�@/f�4p4@�4 ڃ�!?!/��a�@�f7q�ٿ}k�0��@���\�*4@qi���!? l`��@���v]�ٿ��6d�@1�����3@J/��O�!?��Pb�@�*`OF�ٿ�Q��c�@��l,4@VY�R�!?�C��D0�@�*`OF�ٿ�Q��c�@��l,4@VY�R�!?�C��D0�@�*`OF�ٿ�Q��c�@��l,4@VY�R�!?�C��D0�@�*`OF�ٿ�Q��c�@��l,4@VY�R�!?�C��D0�@'i:���ٿ[�0>���@}�"��3@�ә|;�!?�ʣ���@�oS��ٿQ�]b�@`�*��3@T$�c�!?t ,tɴ�@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@�ϐ$��ٿw_�Ήt�@Z�S�d�3@�Co�[�!?
�t%��@o?|&I�ٿ�C(r���@��i�?4@�;�+�!?�󸫅ە@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�#!Zi�ٿV C��@��or4@H�i"�!?�?t>�@�lƜٿ���
I�@|�ԩ�3@e%��!�!?^/�@�lƜٿ���
I�@|�ԩ�3@e%��!�!?^/�@ɤAȜ�ٿ��C����@.٧�~4@�\T�<�!?�?���@ɤAȜ�ٿ��C����@.٧�~4@�\T�<�!?�?���@ɤAȜ�ٿ��C����@.٧�~4@�\T�<�!?�?���@(��߿�ٿ������@.6���$4@�g� �!?�Xa�iԕ@(��߿�ٿ������@.6���$4@�g� �!?�Xa�iԕ@(��߿�ٿ������@.6���$4@�g� �!?�Xa�iԕ@(��߿�ٿ������@.6���$4@�g� �!?�Xa�iԕ@(��߿�ٿ������@.6���$4@�g� �!?�Xa�iԕ@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@[����ٿ�ݫ���@�+��3@��K(�!?+uhh2��@)�	��ٿ8�WLG�@�@��4@j.p�!?�r�ܓ�@�@<���ٿ�aJ����@j�-��4@:�~��!?�X��\�@�@<���ٿ�aJ����@j�-��4@:�~��!?�X��\�@��T�
�ٿ?<b�s�@L�u?�4@���H�!?�)o����@��T�
�ٿ?<b�s�@L�u?�4@���H�!?�)o����@��T�
�ٿ?<b�s�@L�u?�4@���H�!?�)o����@�`�,��ٿ�G	���@�.5��3@���T�!?Zr+�@�`�,��ٿ�G	���@�.5��3@���T�!?Zr+�@�`�,��ٿ�G	���@�.5��3@���T�!?Zr+�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�!aC��ٿB�(�0�@!b����3@�\�^>�!?5Lv��8�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@�Y�¾�ٿ�N���@<��"4@I�ǂ?�!?U"u$�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@MA�Y��ٿ�? �v�@�?�q�4@�*�:�!?�.�E�K�@���q�ٿ�lL���@�,ݾ4@.w?��!?}��C��@���q�ٿ�lL���@�,ݾ4@.w?��!?}��C��@���q�ٿ�lL���@�,ݾ4@.w?��!?}��C��@���q�ٿ�lL���@�,ݾ4@.w?��!?}��C��@�P��ٿvv�.�@��t?#4@$��:��!?���
�@2��CD�ٿ�@�e�@���[�4@f|����!?���&���@V��g�ٿ��ECh��@
�(C�*4@m�F#y�!?�z�4��@V��g�ٿ��ECh��@
�(C�*4@m�F#y�!?�z�4��@V��g�ٿ��ECh��@
�(C�*4@m�F#y�!?�z�4��@V��g�ٿ��ECh��@
�(C�*4@m�F#y�!?�z�4��@V��g�ٿ��ECh��@
�(C�*4@m�F#y�!?�z�4��@ڣ��٤ٿ��s���@��&h�74@bL�G�!?�٥dϕ@ڣ��٤ٿ��s���@��&h�74@bL�G�!?�٥dϕ@ڣ��٤ٿ��s���@��&h�74@bL�G�!?�٥dϕ@r,���ٿ��)1�@���c�(4@��`���!?��
�/�@ܬ_	�ٿ�8 Cݦ�@�Y8yK#4@�;����!?��f�Ǖ@�;�y�ٿǶ8���@ �ѱ2!4@�a�@y�!?(<����@ۈ+Z�ٿh�!ޕ�@���3@�_���!?���试@ۈ+Z�ٿh�!ޕ�@���3@�_���!?���试@ۈ+Z�ٿh�!ޕ�@���3@�_���!?���试@ۈ+Z�ٿh�!ޕ�@���3@�_���!?���试@rY��L�ٿ�m����@̠��H4@�0���!?A^gu۲�@rY��L�ٿ�m����@̠��H4@�0���!?A^gu۲�@rY��L�ٿ�m����@̠��H4@�0���!?A^gu۲�@rY��L�ٿ�m����@̠��H4@�0���!?A^gu۲�@f�v�ٿ��15j�@;ڤݭ54@�	�cw�!?��+���@f�v�ٿ��15j�@;ڤݭ54@�	�cw�!?��+���@f�v�ٿ��15j�@;ڤݭ54@�	�cw�!?��+���@f�v�ٿ��15j�@;ڤݭ54@�	�cw�!?��+���@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@�Ͻ��ٿU��0�J�@<��h4@�	p+��!?��]Ń��@g�(�ٿ�������@!����3@��WVo�!?��9���@g�(�ٿ�������@!����3@��WVo�!?��9���@g�(�ٿ�������@!����3@��WVo�!?��9���@g�(�ٿ�������@!����3@��WVo�!?��9���@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@���O�ٿ�A��FE�@�kKr�4@�MN蜐!?3�A'�ܕ@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@�>�D�ٿ�(m8gm�@��^94@t��\u�!?����@D�mN�ٿy�0E0�@��ʧ484@6�P�!?�rEP���@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�Ƶf~�ٿ{)��`	�@4���?`4@��@�!?Dk�&�@�a;��ٿ�\�	��@S ���A4@G�ўL�!?Ǿ�9��@���ٿ����1�@omJ��+4@��v!x�!?^Oʍ���@���ٿ����1�@omJ��+4@��v!x�!?^Oʍ���@���ٿ����1�@omJ��+4@��v!x�!?^Oʍ���@���ٿ����1�@omJ��+4@��v!x�!?^Oʍ���@R�<O�ٿ�^�g/�@����4@�15�m�!?8����@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@��*��ٿ�-��@ת^�4@)��J�!?�<"ו@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@Y07��ٿ$óY��@��j��3@�[�$�!?<%m��@�l=�ٿ(Ը�N4�@�����3@���{q�!?ڶ��=�@�l=�ٿ(Ը�N4�@�����3@���{q�!?ڶ��=�@�l=�ٿ(Ը�N4�@�����3@���{q�!?ڶ��=�@�@}1�ٿH}�q;�@z�T 4@ͼߺ��!?��'�1ԕ@�@}1�ٿH}�q;�@z�T 4@ͼߺ��!?��'�1ԕ@�@}1�ٿH}�q;�@z�T 4@ͼߺ��!?��'�1ԕ@�@}1�ٿH}�q;�@z�T 4@ͼߺ��!?��'�1ԕ@�@}1�ٿH}�q;�@z�T 4@ͼߺ��!?��'�1ԕ@�$(��ٿK&�1$�@h���4@]���N�!?LDO���@�$(��ٿK&�1$�@h���4@]���N�!?LDO���@��R��ٿ�m��*�@	�D�4@5r�,��!??��x��@��R��ٿ�m��*�@	�D�4@5r�,��!??��x��@��R��ٿ�m��*�@	�D�4@5r�,��!??��x��@��R��ٿ�m��*�@	�D�4@5r�,��!??��x��@��R��ٿ�m��*�@	�D�4@5r�,��!??��x��@����/�ٿ�r��=�@��(�3@��L�*�!?�Y���@�� j��ٿ��&/�@�\՛�3@[��$�!?X׹�zΕ@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@��Qi9�ٿ��FG^�@���34@���"�!? �s%���@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@8d�k��ٿ�� ����@���3A4@wI @B�!?9w�1��@�(d$֞ٿ3����0�@�X)4@1�6�!?$�'�/�@�g�͜ٿ��V�	�@N�Zla4@wi�3�!?�����@�Q�@�ٿ\�	�@n��2�=4@�!��!?{I(}���@�F��|�ٿ�B.g��@��T��	4@|�8�!?�|a��@�F��|�ٿ�B.g��@��T��	4@|�8�!?�|a��@�F��|�ٿ�B.g��@��T��	4@|�8�!?�|a��@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@���?�ٿ������@�H���3@_�� �!?�Xʯ�Ǖ@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@j�a�B�ٿ�Y�.�@�6T�L�3@���!?�z13���@9�.ʵ�ٿ.H1��@��vu4@}#���!?�RT3��@�V%n�ٿC&.���@p�d��)4@4g23x�!?6�	j�ϕ@�V%n�ٿC&.���@p�d��)4@4g23x�!?6�	j�ϕ@�V%n�ٿC&.���@p�d��)4@4g23x�!?6�	j�ϕ@0�4�ٿq�B�G�@��YL64@/�AL��!?s��R��@0�4�ٿq�B�G�@��YL64@/�AL��!?s��R��@0�4�ٿq�B�G�@��YL64@/�AL��!?s��R��@|��|�ٿ�Ug��@���*4@] +u��!?�5���˕@|��|�ٿ�Ug��@���*4@] +u��!?�5���˕@|��|�ٿ�Ug��@���*4@] +u��!?�5���˕@al9�~�ٿ������@����R!4@)RB��!?'�����@al9�~�ٿ������@����R!4@)RB��!?'�����@al9�~�ٿ������@����R!4@)RB��!?'�����@L$���ٿ)�\�9��@�e&>4@���r�!?�ـ:�@L$���ٿ)�\�9��@�e&>4@���r�!?�ـ:�@L$���ٿ)�\�9��@�e&>4@���r�!?�ـ:�@������ٿD�gq�p�@�Pj}v<4@�S��!?�0�"�@������ٿD�gq�p�@�Pj}v<4@�S��!?�0�"�@�9�+�ٿ�\N�r�@vk�+[4@bk�8�!?m�S���@�9�+�ٿ�\N�r�@vk�+[4@bk�8�!?m�S���@�9�+�ٿ�\N�r�@vk�+[4@bk�8�!?m�S���@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@˝�0�ٿ��0����@s��Q4@�㎝��!?��2"�,�@���^�ٿ1{u����@h� ���3@��+ߏ!?���Ʉ��@�;M�ٿ� oT���@�+9��3@�Ҿp,�!?��M��@�;M�ٿ� oT���@�+9��3@�Ҿp,�!?��M��@�;M�ٿ� oT���@�+9��3@�Ҿp,�!?��M��@�;M�ٿ� oT���@�+9��3@�Ҿp,�!?��M��@�duÝ�ٿ�cA�x��@���a��3@����ې!?A2��䧕@�duÝ�ٿ�cA�x��@���a��3@����ې!?A2��䧕@�duÝ�ٿ�cA�x��@���a��3@����ې!?A2��䧕@�duÝ�ٿ�cA�x��@���a��3@����ې!?A2��䧕@�duÝ�ٿ�cA�x��@���a��3@����ې!?A2��䧕@@p��ҟٿ|�2����@&��!�4@`�b���!?�(�p'�@��Y=0�ٿ���S�@���N4@5q�瞐!?�n� ��@��Y=0�ٿ���S�@���N4@5q�瞐!?�n� ��@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@�}�]šٿ�'����@���]"4@��7{�!?���_�@��Aܰ�ٿD9�<��@'�~��3@}��o��!?Q똼��@��Aܰ�ٿD9�<��@'�~��3@}��o��!?Q똼��@��Aܰ�ٿD9�<��@'�~��3@}��o��!?Q똼��@l����ٿ�v�߲��@��$u�3@E#����!?H���[n�@l����ٿ�v�߲��@��$u�3@E#����!?H���[n�@����ٿ�JS��@�O+�;4@�+��g�!?�PA�8F�@����ٿ�JS��@�O+�;4@�+��g�!?�PA�8F�@����ٿ�JS��@�O+�;4@�+��g�!?�PA�8F�@V�h�ٿ�I�t�@h�o��4@�)B�8�!?(��E"�@}�p4˛ٿy��F��@x��bd 4@�lrc�!?s���,�@}�p4˛ٿy��F��@x��bd 4@�lrc�!?s���,�@�]��ٿh���9�@W�>�4@�rD*K�!??�J2���@�]��ٿh���9�@W�>�4@�rD*K�!??�J2���@�]��ٿh���9�@W�>�4@�rD*K�!??�J2���@� L�v�ٿ��~�(�@|��{:4@��S���!?d@wQ�@� L�v�ٿ��~�(�@|��{:4@��S���!?d@wQ�@� L�v�ٿ��~�(�@|��{:4@��S���!?d@wQ�@� L�v�ٿ��~�(�@|��{:4@��S���!?d@wQ�@� L�v�ٿ��~�(�@|��{:4@��S���!?d@wQ�@c�FƠ�ٿ���=��@N���<�3@�;5DY�!?L�\�ŕ@8��he�ٿ�/��R��@����y�3@��*N�!?�l�^��@8��he�ٿ�/��R��@����y�3@��*N�!?�l�^��@X�p�9�ٿ7c�2��@!�04@��2��!?.��Z=�@X�p�9�ٿ7c�2��@!�04@��2��!?.��Z=�@9�g� �ٿ{��#���@5?��e4@h�@Nڐ!?-�p��@Ἵ���ٿ���Q͐�@�3u?�/4@�d��А!?�|  ܕ@ru�J��ٿ�Ɉ�@��=C��3@�pH)��!?���̏�@ru�J��ٿ�Ɉ�@��=C��3@�pH)��!?���̏�@�{�K}�ٿ/�8�.��@�4+7�4@x
�̐!?z�N|��@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@��X�ٿ+\��5�@�W#>.4@��lC��!? >����@�J=��ٿ���ʵg�@�����4@�g�п�!?m�G�/a�@�J=��ٿ���ʵg�@�����4@�g�п�!?m�G�/a�@n+�脡ٿ��"y��@�����3@wC����!?/.���%�@n+�脡ٿ��"y��@�����3@wC����!?/.���%�@n+�脡ٿ��"y��@�����3@wC����!?/.���%�@n+�脡ٿ��"y��@�����3@wC����!?/.���%�@n+�脡ٿ��"y��@�����3@wC����!?/.���%�@@f��f�ٿ~qv�i�@�>V4@�����!?Ӭ���&�@�M �I�ٿ���e��@ t�[�&4@:f2���!?�B�%P�@�M �I�ٿ���e��@ t�[�&4@:f2���!?�B�%P�@+��	�ٿ�'ޥ�S�@�8|C4@`65��!?��&P�a�@+��	�ٿ�'ޥ�S�@�8|C4@`65��!?��&P�a�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@���j+�ٿj��G]�@:��14@���u[�!?�񆍄�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@i��sD�ٿ��uȞ�@�)�Ȗ4@���!?�9Yu:}�@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@џF���ٿ�T�<�[�@�s!n4@��Ց�!?�-�����@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@�.��r�ٿxB����@T�
�34@υ/�w�!?���̂�@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@��A���ٿ%;�����@�cHu�34@�}��u�!?�O��@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@�ݮ�ٿ�ߓ?��@A�kM@4@N��Z$�!?mtJ룕@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@&�r��ٿ�uh��6�@-�*4@����G�!?:_l�	��@t��Ԡٿ�w�"��@��׾�4@)��&��!?���՘�@�L�ٿM������@ƝU.4@G��E�!?��rZ�@�L�ٿM������@ƝU.4@G��E�!?��rZ�@�L�ٿM������@ƝU.4@G��E�!?��rZ�@�L�ٿM������@ƝU.4@G��E�!?��rZ�@�L�ٿM������@ƝU.4@G��E�!?��rZ�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@�P��H�ٿ>���;��@�ƕ�?4@Q@ �?�!?���T�@���"�ٿ�#�4��@W)��4@j�_�l�!?��/�尕@���"�ٿ�#�4��@W)��4@j�_�l�!?��/�尕@���"�ٿ�#�4��@W)��4@j�_�l�!?��/�尕@_��%�ٿ���0=��@p��gb*4@{ky>��!?�G�3*��@_��%�ٿ���0=��@p��gb*4@{ky>��!?�G�3*��@_��%�ٿ���0=��@p��gb*4@{ky>��!?�G�3*��@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@����x�ٿ��)!x;�@/4R)4@y���!?(/��$�@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@AH�5D�ٿ�A7���@؄BN��3@��V
��!?������@}A��֝ٿʷw+��@PP��74@��Yc�!?�J��w�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��24�ٿ�,;1�@���44@f��r�!?Qk��V�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@��v���ٿ#���A�@lԨ���3@
_��q�!?\��i�@t���%�ٿ�<��g/�@��T�.4@�hh5�!?g�E�@t���%�ٿ�<��g/�@��T�.4@�hh5�!?g�E�@t���%�ٿ�<��g/�@��T�.4@�hh5�!?g�E�@u��ٿ@��� �@�Ev>4@�mhJ�!?��r��@u��ٿ@��� �@�Ev>4@�mhJ�!?��r��@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@��r((�ٿ�}����@?�wP�4@9�׃f�!?c$�.Mԕ@U򪟕�ٿ�qԜ��@L�M/4@�,?�!?iK�AaΕ@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@���ٿ���re�@��$74@-)�L�!?[p��S�@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@ބ<�ٿ0h��M�@�y�H�;4@g�w?i�!?Ľ����@�3C�[�ٿ/W�~'�@��$4@�o�99�!?+�`~�@KW�>k�ٿ��8���@�Y��!4@���!?:v��h�@KW�>k�ٿ��8���@�Y��!4@���!?:v��h�@KW�>k�ٿ��8���@�Y��!4@���!?:v��h�@KW�>k�ٿ��8���@�Y��!4@���!?:v��h�@?0��ٿW�M�@�u�e4@X�!�!?�C7���@?0��ٿW�M�@�u�e4@X�!�!?�C7���@?0��ٿW�M�@�u�e4@X�!�!?�C7���@?0��ٿW�M�@�u�e4@X�!�!?�C7���@?0��ٿW�M�@�u�e4@X�!�!?�C7���@�� �ٿ��&�a�@�p-��
4@�ȡuR�!?8��@�� �ٿ��&�a�@�p-��
4@�ȡuR�!?8��@"�j��ٿ�F��#+�@ˬ)A4@~�� L�!?Y8����@"�j��ٿ�F��#+�@ˬ)A4@~�� L�!?Y8����@��,���ٿ���W��@`<.I4@�y$�!?h�o���@�E�z�ٿșQ����@##S^�F4@c�"�R�!?��Cƣ
�@�E�z�ٿșQ����@##S^�F4@c�"�R�!?��Cƣ
�@�E�z�ٿșQ����@##S^�F4@c�"�R�!?��Cƣ
�@�����ٿ]zPܹ�@�\�Y�64@"���!?Ɩ%E��@�����ٿ]zPܹ�@�\�Y�64@"���!?Ɩ%E��@�����ٿ]zPܹ�@�\�Y�64@"���!?Ɩ%E��@�����ٿ]zPܹ�@�\�Y�64@"���!?Ɩ%E��@�����ٿ]zPܹ�@�\�Y�64@"���!?Ɩ%E��@2�f��ٿ�ߗ�^�@D
�eS4@��$D�!?1[ƕ@2�f��ٿ�ߗ�^�@D
�eS4@��$D�!?1[ƕ@2�f��ٿ�ߗ�^�@D
�eS4@��$D�!?1[ƕ@2�f��ٿ�ߗ�^�@D
�eS4@��$D�!?1[ƕ@}����ٿ:�u����@ho�'�24@���V�!?��c-a�@}����ٿ:�u����@ho�'�24@���V�!?��c-a�@}����ٿ:�u����@ho�'�24@���V�!?��c-a�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@4�Xy��ٿ�]v`�I�@Q�5P4@GЯ��!?���>0U�@�;��#�ٿ�{�����@F&��.4@��y�!?űd�XE�@�;��#�ٿ�{�����@F&��.4@��y�!?űd�XE�@P�Y���ٿ)
!$�@ ��O4@KĆ��!? }H�@�`SW�ٿ|��^��@��?J4@98<��!?��� �@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@��'O�ٿ�&㵜�@��|�]4@�	�U�!?D���G�@���ٿ�&^D�O�@��34@�Ȟ��!?�(?K�@���ٿ�&^D�O�@��34@�Ȟ��!?�(?K�@��?T�ٿ���5p�@��"�/4@`��5�!?�4EZ�@��?T�ٿ���5p�@��"�/4@`��5�!?�4EZ�@��?T�ٿ���5p�@��"�/4@`��5�!?�4EZ�@��?T�ٿ���5p�@��"�/4@`��5�!?�4EZ�@��?T�ٿ���5p�@��"�/4@`��5�!?�4EZ�@��Dp�ٿ�k* 6d�@����3@aCσ�!?��M�8�@���%Ιٿ�PT�	��@eҰ*4@)�V�!?0�>n��@���%Ιٿ�PT�	��@eҰ*4@)�V�!?0�>n��@��]��ٿ��Wb�@E�����3@��3��!?�0R�w4�@��]��ٿ��Wb�@E�����3@��3��!?�0R�w4�@ӫfɕٿ��ܿ�@��2�L4@W
����!?E�\��@ӫfɕٿ��ܿ�@��2�L4@W
����!?E�\��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@rV6.�ٿ��u��@��.4@0T=k��!?8"p�^��@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@֡��˛ٿR�G�%��@yo+{4@p؜���!?!4���@��v�3�ٿ��b�<��@����k4@G����!?;JN���@��v�3�ٿ��b�<��@����k4@G����!?;JN���@��v�3�ٿ��b�<��@����k4@G����!?;JN���@�\�x�ٿX7��,�@�i��3@t����!?�%����@+��ٿ�FZ���@?r���3@?3�yU�!?]��h��@+��ٿ�FZ���@?r���3@?3�yU�!?]��h��@+��ٿ�FZ���@?r���3@?3�yU�!?]��h��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@:��@�ٿ��n��@I1r��4@�����!?`�SC��@x�]j�ٿ{1.h�@P�Gyg?4@�{��:�!?�=�
�H�@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@�6���ٿ��hZG�@U4pӰ4@@t
I�!?�� ܕ@ՕG^+�ٿw�c ��@���w�3@H��r��!?���:a�@���ۚٿ3g��_�@RXoU�4@BK	D��!?R��B�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@c���ٿK���(�@���t5@4@�[��a�!?�uѥ�@�%���ٿ������@���64@��5V�!?��Egٕ@�%���ٿ������@���64@��5V�!?��Egٕ@��-	ٿ6�L5]��@�i�"4@y0�>j�!?Jd�u*�@��-	ٿ6�L5]��@�i�"4@y0�>j�!?Jd�u*�@��-	ٿ6�L5]��@�i�"4@y0�>j�!?Jd�u*�@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@���vx�ٿ��"��@��V�d,4@�>S^G�!?����@z��5��ٿ��z2��@��o]��3@��r�!?�l7V�@z��5��ٿ��z2��@��o]��3@��r�!?�l7V�@z��5��ٿ��z2��@��o]��3@��r�!?�l7V�@g��X<�ٿ��M���@��ꚱ�3@�*�l8�!?*z^r��@g��X<�ٿ��M���@��ꚱ�3@�*�l8�!?*z^r��@g��X<�ٿ��M���@��ꚱ�3@�*�l8�!?*z^r��@��E�$�ٿI���_��@p��+�3@�|.=�!?������@��E�$�ٿI���_��@p��+�3@�|.=�!?������@��E�$�ٿI���_��@p��+�3@�|.=�!?������@���%�ٿ*(����@YA���3@���W�!?�F�C\N�@�ɻN��ٿ*��Nn��@k�+g,4@���А!?�03�T6�@1n��z�ٿu��o��@��=�4@?�VE��!?n�o�@1n��z�ٿu��o��@��=�4@?�VE��!?n�o�@1n��z�ٿu��o��@��=�4@?�VE��!?n�o�@1n��z�ٿu��o��@��=�4@?�VE��!?n�o�@1n��z�ٿu��o��@��=�4@?�VE��!?n�o�@23B�ٿ�"�o��@�0�#�3@���+r�!?��� i�@����9�ٿ�6�I1]�@߮�)�(4@	�O��!?��Y��_�@k����ٿY��e�@
~+4@�-р��!?���`��@k����ٿY��e�@
~+4@�-р��!?���`��@9yl&�ٿlD��$��@>���#4@D��h�!?q��Е@9yl&�ٿlD��$��@>���#4@D��h�!?q��Е@9yl&�ٿlD��$��@>���#4@D��h�!?q��Е@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@~�T��ٿ������@oiی.4@��d�!?��\rC��@R����ٿ��,W��@%��v;4@@��3�!?�%�	Ϫ�@�_�*T�ٿv=����@}��"�64@�6���!?0ULR*o�@�_�*T�ٿv=����@}��"�64@�6���!?0ULR*o�@��! ��ٿeڻ��@�(�޵G4@� �ӏ!?Oo�����@��! ��ٿeڻ��@�(�޵G4@� �ӏ!?Oo�����@��! ��ٿeڻ��@�(�޵G4@� �ӏ!?Oo�����@����ٿf��+/k�@ �0��34@#����!?��(!<��@����ٿf��+/k�@ �0��34@#����!?��(!<��@����ٿf��+/k�@ �0��34@#����!?��(!<��@ǂ�h�ٿ� 5����@7�П��3@�����!?�8F�\��@ǂ�h�ٿ� 5����@7�П��3@�����!?�8F�\��@A�����ٿJ�íܔ�@�a��%�3@�d�_�!?�"�t�#�@A�����ٿJ�íܔ�@�a��%�3@�d�_�!?�"�t�#�@A�����ٿJ�íܔ�@�a��%�3@�d�_�!?�"�t�#�@'��a�ٿkKPxf�@f�pFm�3@�h��m�!?�ȴhh��@'��a�ٿkKPxf�@f�pFm�3@�h��m�!?�ȴhh��@"ձ�@�ٿ�;�c=p�@L�M��3@�H���!?_�M��ڕ@"ձ�@�ٿ�;�c=p�@L�M��3@�H���!?_�M��ڕ@"ձ�@�ٿ�;�c=p�@L�M��3@�H���!?_�M��ڕ@��Ƿ�ٿ8<x���@u�_� =4@O>TN^�!? pJ�0�@��Ƿ�ٿ8<x���@u�_� =4@O>TN^�!? pJ�0�@��Ƿ�ٿ8<x���@u�_� =4@O>TN^�!? pJ�0�@��Ƿ�ٿ8<x���@u�_� =4@O>TN^�!? pJ�0�@p��k�ٿc�_:�o�@���>84@��Tx�!?!ϡ9�H�@p��k�ٿc�_:�o�@���>84@��Tx�!?!ϡ9�H�@�� �ɚٿ��"&��@jU�
=4@:e��Z�!?�:��O��@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�*�%��ٿ!9��A�@���1<4@y3P�!?�Zi5�z�@�㰽��ٿ�f��G�@����)4@n{&h�!?~yBt/��@�㰽��ٿ�f��G�@����)4@n{&h�!?~yBt/��@�㰽��ٿ�f��G�@����)4@n{&h�!?~yBt/��@�㰽��ٿ�f��G�@����)4@n{&h�!?~yBt/��@�㰽��ٿ�f��G�@����)4@n{&h�!?~yBt/��@�%��ٿX�In>�@����'N4@K��?�!?��~aV��@�%��ٿX�In>�@����'N4@K��?�!?��~aV��@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@��v]��ٿ\�U
B�@�t��Y4@6�9� �!?cvj���@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@�Է���ٿ}
�����@iC�UF4@�q�0n�!?�M CWO�@��[��ٿ�Ij�V�@�ks�>4@X�ۦ�!?�]�)���@��[��ٿ�Ij�V�@�ks�>4@X�ۦ�!?�]�)���@��[��ٿ�Ij�V�@�ks�>4@X�ۦ�!?�]�)���@�a��ٿ$�����@���xy	4@���\�!?�ty�@��@�a��ٿ$�����@���xy	4@���\�!?�ty�@��@�a��ٿ$�����@���xy	4@���\�!?�ty�@��@���ٿ������@�m��(4@�_�ː!?���H��@���ٿ������@�m��(4@�_�ː!?���H��@���ٿ������@�m��(4@�_�ː!?���H��@���ٿ������@�m��(4@�_�ː!?���H��@���ٿ������@�m��(4@�_�ː!?���H��@���ٿ������@�m��(4@�_�ː!?���H��@9II5٘ٿ�Y�)��@�n��!4@�f^��!?����,'�@9II5٘ٿ�Y�)��@�n��!4@�f^��!?����,'�@9II5٘ٿ�Y�)��@�n��!4@�f^��!?����,'�@9II5٘ٿ�Y�)��@�n��!4@�f^��!?����,'�@����ٿX��цG�@�t�M4@0��Y�!?[���\�@����ٿX��цG�@�t�M4@0��Y�!?[���\�@ԣ����ٿnSKhk�@�_�@4@�ʮs��!?�6���@ԣ����ٿnSKhk�@�_�@4@�ʮs��!?�6���@ԣ����ٿnSKhk�@�_�@4@�ʮs��!?�6���@ך]f�ٿw@��#�@�g��&4@|�o�!?���D��@ך]f�ٿw@��#�@�g��&4@|�o�!?���D��@ך]f�ٿw@��#�@�g��&4@|�o�!?���D��@ך]f�ٿw@��#�@�g��&4@|�o�!?���D��@���
J�ٿ;݈V���@Ie">3*4@�gkݴ�!?����6ʕ@���
J�ٿ;݈V���@Ie">3*4@�gkݴ�!?����6ʕ@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@�&.�ٿ���F���@0�Lq�4@��Zqj�!?-8g9�@7Yܾ��ٿ���ӯ��@ִ��O(4@0��e��!?-t�6ʚ�@7Yܾ��ٿ���ӯ��@ִ��O(4@0��e��!?-t�6ʚ�@���<��ٿ)��Bl�@�$��?�3@R�s�!?$�g��q�@�〵�ٿ��0�F�@�*l�w�3@�.A�!?,d�Θ��@�〵�ٿ��0�F�@�*l�w�3@�.A�!?,d�Θ��@�〵�ٿ��0�F�@�*l�w�3@�.A�!?,d�Θ��@�〵�ٿ��0�F�@�*l�w�3@�.A�!?,d�Θ��@��|O	�ٿ��7�\�@/>���3@'�(M��!?������@��|O	�ٿ��7�\�@/>���3@'�(M��!?������@S� �j�ٿ�#[2a�@M�cu�3@9i�Z�!? %}Ut��@S� �j�ٿ�#[2a�@M�cu�3@9i�Z�!? %}Ut��@��W��ٿ�Jʿ�R�@�<�S��3@�e9��!?R~��5��@��E�M�ٿs�䧬��@^^�	4@&�J]r�!?9��Cz{�@��E�M�ٿs�䧬��@^^�	4@&�J]r�!?9��Cz{�@��E�M�ٿs�䧬��@^^�	4@&�J]r�!?9��Cz{�@��E�M�ٿs�䧬��@^^�	4@&�J]r�!?9��Cz{�@��E�M�ٿs�䧬��@^^�	4@&�J]r�!?9��Cz{�@���=�ٿ��g�@ܭ��>4@V�Y�C�!?��9����@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@"�\y*�ٿ0"��r��@E���t�3@���r�!?GD*x�ٕ@O��]�ٿ����$�@��"�x94@���V��!?6OD�-��@O��]�ٿ����$�@��"�x94@���V��!?6OD�-��@O��]�ٿ����$�@��"�x94@���V��!?6OD�-��@O��]�ٿ����$�@��"�x94@���V��!?6OD�-��@�)�6��ٿ�%G�M�@b���8
4@�º��!?1�F�\��@�)�6��ٿ�%G�M�@b���8
4@�º��!?1�F�\��@�,��I�ٿ�:�%+ �@�;���)4@u�uU�!?�ڿ@�,��I�ٿ�:�%+ �@�;���)4@u�uU�!?�ڿ@ё8�S�ٿ<����I�@1Ú\�4@"P��5�!?�O�Z��@ё8�S�ٿ<����I�@1Ú\�4@"P��5�!?�O�Z��@ё8�S�ٿ<����I�@1Ú\�4@"P��5�!?�O�Z��@ё8�S�ٿ<����I�@1Ú\�4@"P��5�!?�O�Z��@k�)W��ٿ�ђ ��@�^,�6$4@�Z2O��!?�7R�Q�@�ȉ��ٿDK�gG��@�<�nP4@�3����!?��1CH�@*�ʲz�ٿ��h�@���f�3@����B�!?�Ɗ����@*�ʲz�ٿ��h�@���f�3@����B�!?�Ɗ����@*�ʲz�ٿ��h�@���f�3@����B�!?�Ɗ����@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@Y��c�ٿH�����@����;�3@+�=��!?�Y�Z�Z�@C�Ξ�ٿ�n��`��@3��o�3@�j٫}�!?��#�c�@C�Ξ�ٿ�n��`��@3��o�3@�j٫}�!?��#�c�@C�Ξ�ٿ�n��`��@3��o�3@�j٫}�!?��#�c�@C�Ξ�ٿ�n��`��@3��o�3@�j٫}�!?��#�c�@�O��ڙٿ�[{�@�@����3@�%+�S�!?�H?�@z��&ʘٿ������@�Ѳ0��3@�k�t�!?��M��@z��&ʘٿ������@�Ѳ0��3@�k�t�!?��M��@z��&ʘٿ������@�Ѳ0��3@�k�t�!?��M��@z��&ʘٿ������@�Ѳ0��3@�k�t�!?��M��@o�+���ٿWcL?d�@k7E�4@�����!?��Xa�>�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@�����ٿ���
�#�@�b�4@�����!?�'Co"�@:7�s�ٿ�NTC�@L/��E4@-����!?�xq��@:7�s�ٿ�NTC�@L/��E4@-����!?�xq��@:7�s�ٿ�NTC�@L/��E4@-����!?�xq��@�B�tМٿi��Õ=�@�g�54@^�A ��!?eXչ�J�@����ٿ�LAN;�@�/�t4@�n*��!?;��3�ɕ@����ٿ�LAN;�@�/�t4@�n*��!?;��3�ɕ@����ٿ�LAN;�@�/�t4@�n*��!?;��3�ɕ@����ٿ�LAN;�@�/�t4@�n*��!?;��3�ɕ@����ٿ�LAN;�@�/�t4@�n*��!?;��3�ɕ@w!�C�ٿ�K�ʐ��@��V�4@����'�!?(t���@w!�C�ٿ�K�ʐ��@��V�4@����'�!?(t���@w!�C�ٿ�K�ʐ��@��V�4@����'�!?(t���@�!�ϔ�ٿ�g�{�s�@���6�24@���FA�!?�����@G�2z%�ٿ�Aן���@�>E�h>4@����,�!?��R�@G�2z%�ٿ�Aן���@�>E�h>4@����,�!?��R�@;�8���ٿ2���=�@y�Jug;4@/�J%U�!?&�l8\�@;�8���ٿ2���=�@y�Jug;4@/�J%U�!?&�l8\�@;�8���ٿ2���=�@y�Jug;4@/�J%U�!?&�l8\�@�_�l�ٿ�Vp<rR�@9@u�4@�O�!?���J�@�_�l�ٿ�Vp<rR�@9@u�4@�O�!?���J�@�_�l�ٿ�Vp<rR�@9@u�4@�O�!?���J�@�A;��ٿ�)�\s��@�{H1�4@�W�
^�!?l����@�A;��ٿ�)�\s��@�{H1�4@�W�
^�!?l����@@T���ٿ2����@�����3@}�X���!?w^b���@@T���ٿ2����@�����3@}�X���!?w^b���@@T���ٿ2����@�����3@}�X���!?w^b���@@T���ٿ2����@�����3@}�X���!?w^b���@@T���ٿ2����@�����3@}�X���!?w^b���@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@Pp���ٿ;ta:f�@�j�@�3@u�!�ѐ!?��\¾�@�&�/�ٿ�v|��@�¯�4@�����!?�\1��@�&�/�ٿ�v|��@�¯�4@�����!?�\1��@�&�/�ٿ�v|��@�¯�4@�����!?�\1��@�&�/�ٿ�v|��@�¯�4@�����!?�\1��@�O���ٿ}D���O�@�N�#4@R��}�!?����1�@�O���ٿ}D���O�@�N�#4@R��}�!?����1�@�O���ٿ}D���O�@�N�#4@R��}�!?����1�@�O���ٿ}D���O�@�N�#4@R��}�!?����1�@��gX,�ٿ�o���!�@b吊4@"�����!?�aN��ѕ@��gX,�ٿ�o���!�@b吊4@"�����!?�aN��ѕ@��gX,�ٿ�o���!�@b吊4@"�����!?�aN��ѕ@��gX,�ٿ�o���!�@b吊4@"�����!?�aN��ѕ@��gX,�ٿ�o���!�@b吊4@"�����!?�aN��ѕ@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@�ҍ�b�ٿ^:�V��@Ū5rn4@B�1Dy�!?�U���@ۖ>�5�ٿ���0#�@�s��3@��jbC�!?7a�n%�@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@w��(�ٿ�40���@(����3@�jP�!?"\3���@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@��/��ٿk��z��@�c_�@4@�*�v�!?b-�.ʕ@2>�,��ٿU�.3�{�@�^=��3@v#~I��!?� -��@2>�,��ٿU�.3�{�@�^=��3@v#~I��!?� -��@2>�,��ٿU�.3�{�@�^=��3@v#~I��!?� -��@2>�,��ٿU�.3�{�@�^=��3@v#~I��!?� -��@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�gC�ٿ��qC�V�@�tG=��3@J09�!?����F�@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@�ظd��ٿ^1d��v�@�B��~�3@e�jhA�!?��	����@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@w��šٿ���)^��@/�Kj�3@�3';d�!?T�PҀ�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@  �A�ٿ|��C��@����.4@tXE��!?�\lneY�@�c>�ٿ�ʶU�q�@:>���3@(i�}<�!?V�	dD�@�c>�ٿ�ʶU�q�@:>���3@(i�}<�!?V�	dD�@�c>�ٿ�ʶU�q�@:>���3@(i�}<�!?V�	dD�@�c>�ٿ�ʶU�q�@:>���3@(i�}<�!?V�	dD�@��bb$�ٿ>�=Z��@�5�&4@ I�Y��!?�mǝr�@��bb$�ٿ>�=Z��@�5�&4@ I�Y��!?�mǝr�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@y+e�ٿ���l�@太�K,4@=��T�!?�X�!�@T�{�n�ٿ�v�F�@�G�G	4@���Mi�!?�N4A�@��W:M�ٿ%&r��@��^�)4@�#��]�!?r&��/�@��W:M�ٿ%&r��@��^�)4@�#��]�!?r&��/�@��W:M�ٿ%&r��@��^�)4@�#��]�!?r&��/�@F�q�ٿ�g�@Z�#U4@��3�T�!?��8�Z�@=ɰ��ٿG��R�@�����%4@��Av�!?�x��Q��@�@ȴ6�ٿ3@h�(��@Ѳ.�?4@ M?J�!?2bhHҕ@�@ȴ6�ٿ3@h�(��@Ѳ.�?4@ M?J�!?2bhHҕ@�@ȴ6�ٿ3@h�(��@Ѳ.�?4@ M?J�!?2bhHҕ@�@ȴ6�ٿ3@h�(��@Ѳ.�?4@ M?J�!?2bhHҕ@�@ȴ6�ٿ3@h�(��@Ѳ.�?4@ M?J�!?2bhHҕ@��R���ٿ��T�@�ގVC4@O�֐!?��H��2�@��R���ٿ��T�@�ގVC4@O�֐!?��H��2�@�P?���ٿ���@�C�9l4@;��G�!?���sG�@���i�ٿɵ�s���@36x��>4@��J稐!?7؝i4�@75t��ٿlHZV��@�a�a4@��|_�!?�'N�@`�?�ٿ������@ �D4@��>��!?��B���@�D�̽�ٿ�68��@ȫ�}�4@��@eE�!?=�[9ϕ@�D�̽�ٿ�68��@ȫ�}�4@��@eE�!?=�[9ϕ@�D�̽�ٿ�68��@ȫ�}�4@��@eE�!?=�[9ϕ@�D�̽�ٿ�68��@ȫ�}�4@��@eE�!?=�[9ϕ@�Sv:�ٿD<U �@��b)'�3@�S�b&�!?ė�@$��@����ٿ��_T��@�/���3@���!?Bբ+�	�@����ٿ��_T��@�/���3@���!?Bբ+�	�@����ٿ��_T��@�/���3@���!?Bբ+�	�@����ٿ��_T��@�/���3@���!?Bբ+�	�@����ٿ��_T��@�/���3@���!?Bբ+�	�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��!ɝٿLZ.u�F�@��`�4@��!#�!?��|X2�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@��5�ٿ����	�@�}��2�3@���b�!?R�]�@ךͱ��ٿM~;۝��@akx\�4@�r���!?ʳ�%�@ךͱ��ٿM~;۝��@akx\�4@�r���!?ʳ�%�@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@�{�]�ٿG����@���3@	�=�z�!?8�����@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@���*d�ٿ����=��@�WHa��3@1��L�!?fhBI�
�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@K�r�ٿ�P4+�@������3@Mu��E�!?���ưR�@Pi�d�ٿq�[����@c�4@��ӎw�!?�)��-ܕ@��� A�ٿ���Na'�@}iJ��"4@��ճ>�!?#{�\��@��� A�ٿ���Na'�@}iJ��"4@��ճ>�!?#{�\��@���d�ٿe��SI�@�V1��34@��R�v�!?��Ŕ��@���d�ٿe��SI�@�V1��34@��R�v�!?��Ŕ��@��;�ٿr� �	��@��l%4@���:�!?<���S��@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@y7UΆ�ٿ0bh����@2A�Q)4@�4ÇX�!?���t5-�@:�#C�ٿ8J�FlE�@� ��=�3@��G2V�!?�%D�CL�@:�#C�ٿ8J�FlE�@� ��=�3@��G2V�!?�%D�CL�@:�#C�ٿ8J�FlE�@� ��=�3@��G2V�!?�%D�CL�@:�#C�ٿ8J�FlE�@� ��=�3@��G2V�!?�%D�CL�@:�#C�ٿ8J�FlE�@� ��=�3@��G2V�!?�%D�CL�@�D |�ٿ�k}���@��FI"�3@��2��!?jw��X�@�C#�ٿm������@%����3@8"�jr�!?�߁���@�C#�ٿm������@%����3@8"�jr�!?�߁���@�?�עٿ�9<|���@͊���3@��e)l�!?�QL��@=����ٿ|g���&�@L1���4@g�����!? � #�"�@_G8�ٿdዃPD�@Ph�6
4@�T�t�!?h��[}�@_G8�ٿdዃPD�@Ph�6
4@�T�t�!?h��[}�@��J�ٿ�0�8;�@w�bk4@�Y���!?���Hٕ@��J�ٿ�0�8;�@w�bk4@�Y���!?���Hٕ@��J�ٿ�0�8;�@w�bk4@�Y���!?���Hٕ@��J�ٿ�0�8;�@w�bk4@�Y���!?���Hٕ@��J�ٿ�0�8;�@w�bk4@�Y���!?���Hٕ@EU� �ٿ�f��9�@I�q�3@������!?�ڰH	�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@٨�P֜ٿv��eA0�@��Ĕ�3@9k��
�!?Ve�I�]�@HIP�ٿ'|�o��@�����3@��d� �!?u\�9�`�@HIP�ٿ'|�o��@�����3@��d� �!?u\�9�`�@HIP�ٿ'|�o��@�����3@��d� �!?u\�9�`�@HIP�ٿ'|�o��@�����3@��d� �!?u\�9�`�@�,�ϥٿ��Y ?��@"�r��3@3A0Ϙ�!?%dg|P�@�,�ϥٿ��Y ?��@"�r��3@3A0Ϙ�!?%dg|P�@�,�ϥٿ��Y ?��@"�r��3@3A0Ϙ�!?%dg|P�@ͩ6���ٿr#� �@>�f4@U�	衐!?�ڿp�@�@��ٿe��2��@�>L��3@8"�琐!?^Su>5��@�@��ٿe��2��@�>L��3@8"�琐!?^Su>5��@�@��ٿe��2��@�>L��3@8"�琐!?^Su>5��@�@��ٿe��2��@�>L��3@8"�琐!?^Su>5��@������ٿ�gjXTq�@����
4@B�C�!?�А�Qȕ@������ٿ�gjXTq�@����
4@B�C�!?�А�Qȕ@������ٿ�gjXTq�@����
4@B�C�!?�А�Qȕ@[=��x�ٿ���?�/�@�Y��4@��FF�!?�H���@[=��x�ٿ���?�/�@�Y��4@��FF�!?�H���@[=��x�ٿ���?�/�@�Y��4@��FF�!?�H���@�bD#�ٿ�����@=O��N4@����!?�H,}Jq�@�bD#�ٿ�����@=O��N4@����!?�H,}Jq�@�bD#�ٿ�����@=O��N4@����!?�H,}Jq�@�bD#�ٿ�����@=O��N4@����!?�H,}Jq�@ʓv�ٿ�n�w��@�'34@��O[�!?�H��D��@�"x�Şٿ�"sI���@%��24@W�Y_X�!?7 ����@�"x�Şٿ�"sI���@%��24@W�Y_X�!?7 ����@�"x�Şٿ�"sI���@%��24@W�Y_X�!?7 ����@���ٿ
������@��'Y�44@�U��!?i�0r�ĕ@z���3�ٿ'~�m��@h�aM�(4@�,dlЏ!?<����@z���3�ٿ'~�m��@h�aM�(4@�,dlЏ!?<����@z���3�ٿ'~�m��@h�aM�(4@�,dlЏ!?<����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@�;Li��ٿ�0�N��@3W�n�4@	6d���!?����@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@���dšٿ���ׂ��@�c2m4@�g�v�!?�#g��7�@��Q1�ٿ��gh�H�@ӝ��6,4@�ѧ��!?�;(:ڕ@��Q1�ٿ��gh�H�@ӝ��6,4@�ѧ��!?�;(:ڕ@��Q1�ٿ��gh�H�@ӝ��6,4@�ѧ��!?�;(:ڕ@�\H�ٿ^j��W��@q�ơ�?4@��wfڐ!?�Qr�q��@�\H�ٿ^j��W��@q�ơ�?4@��wfڐ!?�Qr�q��@$P�&i�ٿ���mn�@C���h!4@��ѐ!?2��ĕ@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@��JZ�ٿ�b����@�a�_4@\#��ߐ!?�1�+f��@�Ck](�ٿv)Z{��@��g�s"4@�F��!?�<a�튕@�Ck](�ٿv)Z{��@��g�s"4@�F��!?�<a�튕@�Ck](�ٿv)Z{��@��g�s"4@�F��!?�<a�튕@�Ck](�ٿv)Z{��@��g�s"4@�F��!?�<a�튕@�Ck](�ٿv)Z{��@��g�s"4@�F��!?�<a�튕@w!�»�ٿH�S�S��@3iG�:4@���3��!?�ժԕ@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�7��ٿY`rl[�@�z�T4@����!?@�w�i�@�%�]k�ٿ�*�'�@yĀ1��3@��qː!?�F;�6�@��e��ٿ�h���@�F��^�3@�Ly�!?q�ԕ�Ǖ@��e��ٿ�h���@�F��^�3@�Ly�!?q�ԕ�Ǖ@��e��ٿ�h���@�F��^�3@�Ly�!?q�ԕ�Ǖ@��e��ٿ�h���@�F��^�3@�Ly�!?q�ԕ�Ǖ@�~�15�ٿ��'H˭�@�R���-4@Y�����!?n�Dd�e�@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@t�=੣ٿ%}��@?Q���3@��΂�!?���`d��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@�60�A�ٿ�+d&��@�#��4@�+>�1�!?t�f��@00R~V�ٿqO�ޯ��@� ��C4@��\12�!?��c�ek�@00R~V�ٿqO�ޯ��@� ��C4@��\12�!?��c�ek�@00R~V�ٿqO�ޯ��@� ��C4@��\12�!?��c�ek�@00R~V�ٿqO�ޯ��@� ��C4@��\12�!?��c�ek�@00R~V�ٿqO�ޯ��@� ��C4@��\12�!?��c�ek�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@R@�UR�ٿ��f�Y�@P�<�R4@�ʗ	�!?�W�9�.�@ã*���ٿ��yt��@>o�54@�75�!?�/�=2B�@ã*���ٿ��yt��@>o�54@�75�!?�/�=2B�@ã*���ٿ��yt��@>o�54@�75�!?�/�=2B�@ã*���ٿ��yt��@>o�54@�75�!?�/�=2B�@�^�,�ٿ��}Y�=�@�]�\�94@����:�!?)#X��@�^�,�ٿ��}Y�=�@�]�\�94@����:�!?)#X��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@��pi:�ٿ)���s�@�����A4@H*Vx�!?h\��}��@o�)/��ٿ-Z'�@�h�L�4@���e�!?_!�:�@o�)/��ٿ-Z'�@�h�L�4@���e�!?_!�:�@���ٿ�|�H�@n��J��3@<�124�!?#Ӽ�A��@���ٿ�|�H�@n��J��3@<�124�!?#Ӽ�A��@	%�Xa�ٿZ�J��@�G��j�3@�d���!?H�q�P �@�)}�ٿ@�A�b��@�d���3@�����!?��pø�@�)}�ٿ@�A�b��@�d���3@�����!?��pø�@�)}�ٿ@�A�b��@�d���3@�����!?��pø�@�)}�ٿ@�A�b��@�d���3@�����!?��pø�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@��).�ٿ�U�,�@8DFB! 4@���w�!?6�HKɃ�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@R �w�ٿ};p�@۷Q#(4@�#�rc�!?�.Lh�@�d��śٿyd��_
�@���GD'4@�nѦ��!?��o6�@�d��śٿyd��_
�@���GD'4@�nѦ��!?��o6�@�d��śٿyd��_
�@���GD'4@�nѦ��!?��o6�@y�$c�ٿ��A�
R�@]^�M�'4@]�>S�!?�k%{��@y�$c�ٿ��A�
R�@]^�M�'4@]�>S�!?�k%{��@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@(� ù�ٿ�B=���@g3�Ur�3@SC��!?��_ͮ�@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��M^��ٿ�yt]	%�@��J��3@]�-��!?����@��qɯ�ٿ�`�': �@*�on(�3@3:EgU�!?ѡې�ȕ@��qɯ�ٿ�`�': �@*�on(�3@3:EgU�!?ѡې�ȕ@��qɯ�ٿ�`�': �@*�on(�3@3:EgU�!?ѡې�ȕ@��qɯ�ٿ�`�': �@*�on(�3@3:EgU�!?ѡې�ȕ@��qɯ�ٿ�`�': �@*�on(�3@3:EgU�!?ѡې�ȕ@YʣL>�ٿ��c,���@���H	4@�]�X�!?�EA{�ŕ@��9"�ٿ�+pY��@���w�3@$�`Y�!?��v[�@��9"�ٿ�+pY��@���w�3@$�`Y�!?��v[�@��9"�ٿ�+pY��@���w�3@$�`Y�!?��v[�@k�Q'��ٿ��z1�k�@B�=9�3@.GK:p�!?�������@k�Q'��ٿ��z1�k�@B�=9�3@.GK:p�!?�������@L�Y���ٿ�=�\�(�@Q����3@Y2o���!?�
�ؕ@L�Y���ٿ�=�\�(�@Q����3@Y2o���!?�
�ؕ@L�Y���ٿ�=�\�(�@Q����3@Y2o���!?�
�ؕ@L�Y���ٿ�=�\�(�@Q����3@Y2o���!?�
�ؕ@������ٿ�=�{M��@ȁ�g4@��?�!? G���@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@���\W�ٿ��T����@��u�94@� ��!?.'���&�@�Vܠ��ٿ,�sN�k�@I��i/4@]׿�Z�!?Jo.:��@�Vܠ��ٿ,�sN�k�@I��i/4@]׿�Z�!?Jo.:��@pK&[�ٿz�UiB�@����r#4@Cw��9�!?�dn^���@pK&[�ٿz�UiB�@����r#4@Cw��9�!?�dn^���@pK&[�ٿz�UiB�@����r#4@Cw��9�!?�dn^���@pK&[�ٿz�UiB�@����r#4@Cw��9�!?�dn^���@fW�ܶ�ٿP�3��@|��i@4@���~ُ!?M��,	�@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@	��Οٿ���!*\�@�Ww�4@�$��(�!?(��Q�ɕ@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@+Ǖ^t�ٿ����3��@���"S94@yJ�G/�!?k6�R8\�@7F����ٿ�h�� �@���v�4@u^�!?�#H��#�@��Ҝ��ٿY���W��@��:rx�3@=i��W�!?ZY�rH�@��ܖٿb�����@)��-O4@�s��o�!?�F�ǳ��@K����ٿ'�
���@���r�4@c�Br2�!?�y���O�@K����ٿ'�
���@���r�4@c�Br2�!?�y���O�@���$x�ٿ��U��@sH24@��KMM�!?�/��@���$x�ٿ��U��@sH24@��KMM�!?�/��@���$x�ٿ��U��@sH24@��KMM�!?�/��@���$x�ٿ��U��@sH24@��KMM�!?�/��@Q��M�ٿRr�ǔ��@{\��H#4@��<K��!?t0Ul���@Q��M�ٿRr�ǔ��@{\��H#4@��<K��!?t0Ul���@Q��M�ٿRr�ǔ��@{\��H#4@��<K��!?t0Ul���@�T��ٿ�R/i�@�bY�3@E�헐!?��f�&�@�T��ٿ�R/i�@�bY�3@E�헐!?��f�&�@�T��ٿ�R/i�@�bY�3@E�헐!?��f�&�@Rc���ٿ%5,�d��@�
���4@<?Wx��!?���f��@�NW��ٿ������@iߜ�+14@H��h�!?��T�l�@�NW��ٿ������@iߜ�+14@H��h�!?��T�l�@�NW��ٿ������@iߜ�+14@H��h�!?��T�l�@GUF��ٿz���4��@|5���4@C�M,|�!?W��@Е@.��D��ٿ
� ����@\����'4@ڞ_�ܐ!?(�Í�ؕ@k�ύ.�ٿ�܍���@����:4@�p���!?V�W����@k�ύ.�ٿ�܍���@����:4@�p���!?V�W����@k�ύ.�ٿ�܍���@����:4@�p���!?V�W����@�qyL�ٿ�G ���@��^�_4@@J��Đ!?�1Q�lȕ@�qyL�ٿ�G ���@��^�_4@@J��Đ!?�1Q�lȕ@�qyL�ٿ�G ���@��^�_4@@J��Đ!?�1Q�lȕ@�qyL�ٿ�G ���@��^�_4@@J��Đ!?�1Q�lȕ@�g�y	�ٿ;&�����@5�ͧs4@��I��!?8峿��@�g�y	�ٿ;&�����@5�ͧs4@��I��!?8峿��@�g�y	�ٿ;&�����@5�ͧs4@��I��!?8峿��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@N�!�	�ٿB\��@e�k4@�s�-y�!?UC�"`��@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@��7��ٿ�� </�@���W'l4@��㛐!?'-� �@����ٿ䱣6��@�O��1:4@�uNym�!?4�E�\��@����ٿ䱣6��@�O��1:4@�uNym�!?4�E�\��@����ٿ䱣6��@�O��1:4@�uNym�!?4�E�\��@=huܖٿS�7zb�@��<��4@\��
�!?��i~J�@�9Jbq�ٿ��=�Z�@����44@���g�!?���9%��@�f��ٿgqL���@ڱ�yAJ4@/&�O�!?F��;��@ʋ|�ٿw����@ÉDv�3@2���!?�N}b��@ʋ|�ٿw����@ÉDv�3@2���!?�N}b��@�Q~�ٿ�\F<l�@����4@���a��!?�˥���@�Q~�ٿ�\F<l�@����4@���a��!?�˥���@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@��G䥡ٿ��c2�@b�O�4@� k�a�!?{��-ŕ@(up�ٿN�;�Hj�@ʬ���4@��"��!?� u Z��@Z��� �ٿ}��
�O�@�`^�4@�I�S��!?!�\��	�@Z��� �ٿ}��
�O�@�`^�4@�I�S��!?!�\��	�@Z��� �ٿ}��
�O�@�`^�4@�I�S��!?!�\��	�@Z��� �ٿ}��
�O�@�`^�4@�I�S��!?!�\��	�@Z��� �ٿ}��
�O�@�`^�4@�I�S��!?!�\��	�@U�Y�ؗٿ�`����@�Qm3��3@���L�!?��\9Fʕ@U�Y�ؗٿ�`����@�Qm3��3@���L�!?��\9Fʕ@U�Y�ؗٿ�`����@�Qm3��3@���L�!?��\9Fʕ@U�Y�ؗٿ�`����@�Qm3��3@���L�!?��\9Fʕ@U ��d�ٿN��"Z0�@�`rT��3@�ww�!??����ؕ@U ��d�ٿN��"Z0�@�`rT��3@�ww�!??����ؕ@U ��d�ٿN��"Z0�@�`rT��3@�ww�!??����ؕ@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@���BG�ٿ����L��@C@�Ԑ�3@��g�b�!?"��Y���@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@Z~�~H�ٿ~����@U?�)4@m>i4H�!?�[�P֊�@�z7�ٿ���]N��@5;3\;4@Y�0�!?�����@�z7�ٿ���]N��@5;3\;4@Y�0�!?�����@�z7�ٿ���]N��@5;3\;4@Y�0�!?�����@�z7�ٿ���]N��@5;3\;4@Y�0�!?�����@�z7�ٿ���]N��@5;3\;4@Y�0�!?�����@<��Z��ٿ�ܯ���@d�X4@W��Q�!?����5��@<��Z��ٿ�ܯ���@d�X4@W��Q�!?����5��@<��Z��ٿ�ܯ���@d�X4@W��Q�!?����5��@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@�~�¡ٿ<�ȥ�(�@�n��Y4@k�Ʉ5�!?��)mE�@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@ؘf��ٿ(v]}W�@X��3@���N=�!?:7[q��@){ >�ٿ�s�u6s�@�k���3@�! H�!?�e��@NfC=��ٿS��i��@�a�	<�3@����L�!?��6	��@NfC=��ٿS��i��@�a�	<�3@����L�!?��6	��@NfC=��ٿS��i��@�a�	<�3@����L�!?��6	��@NfC=��ٿS��i��@�a�	<�3@����L�!?��6	��@NfC=��ٿS��i��@�a�	<�3@����L�!?��6	��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@��6�ٿ���$�@  UE&�3@[|m;.�!?@~X*`��@e�5���ٿ����
��@�Ǣ��4@<y��!?�x�<�@e�5���ٿ����
��@�Ǣ��4@<y��!?�x�<�@tR��ٿ詁O�@0u�A� 4@�v�G&�!?퍼�Օ@tR��ٿ詁O�@0u�A� 4@�v�G&�!?퍼�Օ@tR��ٿ詁O�@0u�A� 4@�v�G&�!?퍼�Օ@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@ap��!�ٿ�y$����@��K*z�3@hz��*�!?YOm�!�@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@<"��J�ٿV;7#�@��Q
nK4@�\�R�!?�[���@�u�ڗ�ٿP��a,d�@jto�4@�j��!? �W���@�u�ڗ�ٿP��a,d�@jto�4@�j��!? �W���@�u�ڗ�ٿP��a,d�@jto�4@�j��!? �W���@�u�ڗ�ٿP��a,d�@jto�4@�j��!? �W���@���/�ٿ����V`�@@�"�Y4@�x4��!?�ɺl(��@���/�ٿ����V`�@@�"�Y4@�x4��!?�ɺl(��@���/�ٿ����V`�@@�"�Y4@�x4��!?�ɺl(��@���/�ٿ����V`�@@�"�Y4@�x4��!?�ɺl(��@�Z�x�ٿl�
���@m���:4@���[�!?C�����@�Z�x�ٿl�
���@m���:4@���[�!?C�����@�Z�x�ٿl�
���@m���:4@���[�!?C�����@�Z�x�ٿl�
���@m���:4@���[�!?C�����@�Z�x�ٿl�
���@m���:4@���[�!?C�����@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@���u�ٿC9����@f��S�4@�=�u:�!?r���Qɕ@��H�"�ٿ�a���l�@ԡU��4@�n���!?����@�����ٿ{D�SO�@1�n�_<4@���?�!?*�`�Ö@ș,��ٿ�%`�z�@�c�d|4@�7��d�!?�"U�@ș,��ٿ�%`�z�@�c�d|4@�7��d�!?�"U�@9P2<�ٿ���j��@�CYt4@f��'S�!?�Nq�[�@9P2<�ٿ���j��@�CYt4@f��'S�!?�Nq�[�@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����աٿGu F�@6	�6�
4@		��Q�!?+TO$��@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@����\�ٿcPG�0��@�$��3@�߻j�!?��(�L�@�#,�S�ٿ�ʟ&�@�0�l("4@��X
�!?d�Y�Bq�@J(��ٿ�j.���@��*��d4@L[��v�!?)�Y��@J(��ٿ�j.���@��*��d4@L[��v�!?)�Y��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@v�6�F�ٿB +�v�@ӤQ��-4@�}K)7�!?p�Xج��@6U����ٿZ.eL�@ȁ|X�+4@N%m�!?b���/�@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�V�AJ�ٿ:2���U�@�x��"4@ ]�{�!?�	��W˕@�7w��ٿ�ڶK�@�b�PM4@|�IX�!?V����ە@�7w��ٿ�ڶK�@�b�PM4@|�IX�!?V����ە@�7w��ٿ�ڶK�@�b�PM4@|�IX�!?V����ە@�7w��ٿ�ڶK�@�b�PM4@|�IX�!?V����ە@�7w��ٿ�ڶK�@�b�PM4@|�IX�!?V����ە@:(sY�ٿ���T�h�@���҂�3@ �N��!?͸�����@:(sY�ٿ���T�h�@���҂�3@ �N��!?͸�����@�C��ٿ�h��
�@�G�>��3@���8g�!?{��4��@�C��ٿ�h��
�@�G�>��3@���8g�!?{��4��@�C��ٿ�h��
�@�G�>��3@���8g�!?{��4��@�C��ٿ�h��
�@�G�>��3@���8g�!?{��4��@�C��ٿ�h��
�@�G�>��3@���8g�!?{��4��@��:h��ٿ�Y:v�w�@�r�	�3@���qh�!?���'AM�@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@i���ٿ���]2��@9���4@��oQ7�!?�	u�<��@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@�U�x�ٿ�R�-�@��]4@�Ġc�!?��h����@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@g���s�ٿ��
J��@3Hn�?4@��C&��!?9���@�+�C&�ٿ�f�F�@Ɓ(4@��u{�!?6}�M�6�@�+�C&�ٿ�f�F�@Ɓ(4@��u{�!?6}�M�6�@�+�C&�ٿ�f�F�@Ɓ(4@��u{�!?6}�M�6�@�Oz,�ٿz2)�hc�@��N�� 4@�@�\v�!?�Ǖ<��@�Oz,�ٿz2)�hc�@��N�� 4@�@�\v�!?�Ǖ<��@�Oz,�ٿz2)�hc�@��N�� 4@�@�\v�!?�Ǖ<��@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@EN`�e�ٿ*r�!���@P�@С+4@����A�!?�k���l�@!���ٿ 'gZA�@X�F��3@Wz-Ӏ�!?�O�Ϲ�@!���ٿ 'gZA�@X�F��3@Wz-Ӏ�!?�O�Ϲ�@!���ٿ 'gZA�@X�F��3@Wz-Ӏ�!?�O�Ϲ�@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@����[�ٿ��R���@��|#4@��髐!?� �N��@�*�B��ٿ���r��@�!4@X�K���!?���Õ@�*�B��ٿ���r��@�!4@X�K���!?���Õ@�*�B��ٿ���r��@�!4@X�K���!?���Õ@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@� ����ٿ�E�G��@�#t�A4@�]�2#�!?E�ҎF�@6q�xޟٿ����T�@�Ԑ��-4@>��D�!?	4�W�@6q�xޟٿ����T�@�Ԑ��-4@>��D�!?	4�W�@BD�x��ٿɋoV)�@Jd<B��3@��n�>�!?��b�+�@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���A�ٿ���@���@!���3@_w�Of�!?��6���@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@���͠ٿ �+��@��=+��3@pfT�!?F�F�&��@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��4l�ٿ��jye��@be ��4@}��!? \[���@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@��K9��ٿle�"Q�@�v�*04@,��Q�!??��`i9�@0���`�ٿ�ڵ�A��@:�6��}4@.3�2K�!?U�����@0���`�ٿ�ڵ�A��@:�6��}4@.3�2K�!?U�����@td
LY�ٿۦf�g��@q�n	L4@���D�!?c�2~��@Vg��`�ٿ�Ct���@8�T^e4@9�^�!?��X!�ɕ@Vg��`�ٿ�Ct���@8�T^e4@9�^�!?��X!�ɕ@Vg��`�ٿ�Ct���@8�T^e4@9�^�!?��X!�ɕ@�J	�U�ٿF�C�@�1��!�3@�w�p��!?8�֔O��@�:wK�ٿ��k�j��@��"��3@d���x�!?.���ו@����X�ٿ"�Ck��@j3 U�3@vHb�)�!?
~) q3�@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@҈���ٿ8Zq$`r�@���+5�3@�?�D�!?��(/>��@#���ٿZ�M�U��@>�;M�14@*Q-m>�!?����F�@#���ٿZ�M�U��@>�;M�14@*Q-m>�!?����F�@#���ٿZ�M�U��@>�;M�14@*Q-m>�!?����F�@#���ٿZ�M�U��@>�;M�14@*Q-m>�!?����F�@#���ٿZ�M�U��@>�;M�14@*Q-m>�!?����F�@AƸ~�ٿ��67��@2<��j4@�žXd�!?[�s�ԕ@AƸ~�ٿ��67��@2<��j4@�žXd�!?[�s�ԕ@AƸ~�ٿ��67��@2<��j4@�žXd�!?[�s�ԕ@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@u��ٿ��f|�1�@"��A�3@yk!m��!? bA�@�yTg�ٿX���@}M;�.4@-�R���!?�7 Q(�@�yTg�ٿX���@}M;�.4@-�R���!?�7 Q(�@-�_`Ŝٿv�J���@c��3@e/�Q�!?t�I�.�@-�_`Ŝٿv�J���@c��3@e/�Q�!?t�I�.�@-�_`Ŝٿv�J���@c��3@e/�Q�!?t�I�.�@}��C=�ٿ0��	��@7�q�4@�Թ5�!?��^��@*K
j��ٿ)$$����@��Ã!4@��ϥZ�!?.*�v��@*K
j��ٿ)$$����@��Ã!4@��ϥZ�!?.*�v��@f �+�ٿ-l^eP�@P3���3@���e�!?%w�&�֕@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@�(�fr�ٿ��^u�+�@i�5�4@���}m�!?��*᫹�@���Ω�ٿ �B ��@f7yW�4@���!?J|�]@�@���Ω�ٿ �B ��@f7yW�4@���!?J|�]@�@��ަi�ٿB��	��@�57��4@�^�)�!?�6P��0�@��ަi�ٿB��	��@�57��4@�^�)�!?�6P��0�@��ަi�ٿB��	��@�57��4@�^�)�!?�6P��0�@}1�̛ٿ2�(1�@��L��3@@&,�'�!?)ߐ���@�P\1�ٿ���V�@�ࢻQ�3@�m#�!?�@�4�͕@�P\1�ٿ���V�@�ࢻQ�3@�m#�!?�@�4�͕@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@ҢP��ٿ&4fY�@`�*[
4@�BP~�!?B[b!K�@��d�ٿ»5܀�@.��Y/4@�9/C�!?Hr�P�ݕ@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�\}�9�ٿ���.C�@3_ӗ�64@L� �^�!?z����@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@�.���ٿ����� �@ǔH-:4@�gO�:�!? @�3�ܕ@qxϹ�ٿ:�F%���@WPG��3@3�T�!?|�t�ϕ@eQDa�ٿ�1a�;��@ٝ�.4@;L�Z&�!?��5l���@eQDa�ٿ�1a�;��@ٝ�.4@;L�Z&�!?��5l���@1�<1�ٿ��[h/�@E�aSr�3@�76~�!?�AraB�@1�<1�ٿ��[h/�@E�aSr�3@�76~�!?�AraB�@1�<1�ٿ��[h/�@E�aSr�3@�76~�!?�AraB�@1�<1�ٿ��[h/�@E�aSr�3@�76~�!?�AraB�@�����ٿ	����@�ܒ��3@�j�b�!?�|��'�@�����ٿ	����@�ܒ��3@�j�b�!?�|��'�@�VH�ٿ8���>��@~��O��3@���t(�!?~�޳/�@�VH�ٿ8���>��@~��O��3@���t(�!?~�޳/�@�	��y�ٿ��t��u�@"�1��3@�΢ #�!?��!(� �@=g�Sq�ٿjj2�#�@��/�
�3@�%Տ!?�F-�C�@�0*m�ٿ��c
���@��≷4@	P���!?�.o��@�0*m�ٿ��c
���@��≷4@	P���!?�.o��@q��p�ٿ�R����@-.�>94@��g1�!?��dÕ@q��p�ٿ�R����@-.�>94@��g1�!?��dÕ@q��p�ٿ�R����@-.�>94@��g1�!?��dÕ@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@9\�f�ٿ���o:��@B=�@�74@A:/�2�!?�=O
��@���8�ٿR*�ޑe�@/`�j�A4@�U\vH�!?q�#��B�@r�t�ٿZ�����@k��/4@G
S�A�!?�c�K��@N<�ٿ6o�$R�@�Y�5
4@�_���!?iȭʽ8�@�1Ŭd�ٿ���G�@��K�#4@���-�!?s�85�6�@�1Ŭd�ٿ���G�@��K�#4@���-�!?s�85�6�@ƣ�ڒ�ٿ�6�[3��@h=a~y�3@eF�=�!?�
�m�ĕ@ƣ�ڒ�ٿ�6�[3��@h=a~y�3@eF�=�!?�
�m�ĕ@ƣ�ڒ�ٿ�6�[3��@h=a~y�3@eF�=�!?�
�m�ĕ@�"���ٿ�i2$��@8sʩ24@�`|�!?D� �@�"���ٿ�i2$��@8sʩ24@�`|�!?D� �@�"���ٿ�i2$��@8sʩ24@�`|�!?D� �@�"���ٿ�i2$��@8sʩ24@�`|�!?D� �@A���/�ٿ%�$��@�,4@����3�!?ׇ2��@A���/�ٿ%�$��@�,4@����3�!?ׇ2��@A���/�ٿ%�$��@�,4@����3�!?ׇ2��@A���/�ٿ%�$��@�,4@����3�!?ׇ2��@��7�ٿ����G��@� ?G)4@��#�!?� ���@h�{9�ٿT:K��V�@?���44@��ck�!?D*�׫��@h�{9�ٿT:K��V�@?���44@��ck�!?D*�׫��@h�{9�ٿT:K��V�@?���44@��ck�!?D*�׫��@h�{9�ٿT:K��V�@?���44@��ck�!?D*�׫��@>����ٿN�kM��@pv�S4@����!?�����@>����ٿN�kM��@pv�S4@����!?�����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@�@��ٿ`X�m�@G�*b�3@�]�d<�!?����@՚�+��ٿͬ�i��@$v��3@��y��!?�M�=ޕ@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�{B���ٿ��G�A�@궧/9�3@b4�!?۫.�̕@�u�^�ٿH���Ld�@�w㭒�3@���X�!?-n6���@�u�^�ٿH���Ld�@�w㭒�3@���X�!?-n6���@�u�^�ٿH���Ld�@�w㭒�3@���X�!?-n6���@���;�ٿj���@*]8V&4@���z�!?n�Yp���@����ٿk�?�gC�@���)4@|�!?d�zn�@eG���ٿ�Bg��@�@Xb{4�4@;����!?1Gy�̕@eG���ٿ�Bg��@�@Xb{4�4@;����!?1Gy�̕@���c�ٿ����O�@
���S4@_>�<�!?��Te��@���c�ٿ����O�@
���S4@_>�<�!?��Te��@���c�ٿ����O�@
���S4@_>�<�!?��Te��@ ��2��ٿj�^p�@�G��"4@�M�Q�!?dÇ봕@�O�.�ٿ>�l���@s�V)�4@3͛�Y�!?�V��d�@�O�.�ٿ>�l���@s�V)�4@3͛�Y�!?�V��d�@�p�ۏ�ٿڌ�X���@vQ�d4@!IRO��!?$�C�3��@�p�ۏ�ٿڌ�X���@vQ�d4@!IRO��!?$�C�3��@�p�ۏ�ٿڌ�X���@vQ�d4@!IRO��!?$�C�3��@�p�ۏ�ٿڌ�X���@vQ�d4@!IRO��!?$�C�3��@�p�ۏ�ٿڌ�X���@vQ�d4@!IRO��!?$�C�3��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@hXi�m�ٿCW��E�@��*f4@JC�Z0�!?Y��"j��@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��8�g�ٿ��� D�@����3@׵ 3E�!?�r�r�ە@��V�Z�ٿɁ�#�U�@� �Y 4@�b��t�!?@SWL軕@��V�Z�ٿɁ�#�U�@� �Y 4@�b��t�!?@SWL軕@������ٿ�Me�b-�@��t!4@�� Y}�!?�qY�R�@������ٿ�Me�b-�@��t!4@�� Y}�!?�qY�R�@A_e���ٿ!P��u�@%:��4@�I5�!?y��_͕@A_e���ٿ!P��u�@%:��4@�I5�!?y��_͕@A_e���ٿ!P��u�@%:��4@�I5�!?y��_͕@A_e���ٿ!P��u�@%:��4@�I5�!?y��_͕@A_e���ٿ!P��u�@%:��4@�I5�!?y��_͕@���D�ٿtz13��@�.�"4@���I��!?r_�It��@�UN�k�ٿ�<��)�@�a���3@>�k�!?��2���@)����ٿ��&���@��?8G4@w��ko�!?����v�@)����ٿ��&���@��?8G4@w��ko�!?����v�@�G&	�ٿ�%�nq�@0�w�-M4@ju5Cl�!?@vb�KT�@�{�DE�ٿ�jbVf��@����&4@&G3,�!?�_���@�{�DE�ٿ�jbVf��@����&4@&G3,�!?�_���@�{�DE�ٿ�jbVf��@����&4@&G3,�!?�_���@�� ��ٿ#�YpC��@��u��?4@��놃�!?�&���@�� ��ٿ#�YpC��@��u��?4@��놃�!?�&���@�� ��ٿ#�YpC��@��u��?4@��놃�!?�&���@�� ��ٿ#�YpC��@��u��?4@��놃�!?�&���@�4��ٿ�f\�_�@oy@r'4@�3�ݞ�!?������@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@�w�kU�ٿ���ψ*�@B�0��4@�4���!?Y��|ѕ@i��l�ٿ��4����@D�`��3@N�f!t�!?*�@�@i��l�ٿ��4����@D�`��3@N�f!t�!?*�@�@3��"�ٿ)w�a|�@Dr����3@��:�!?�j���a�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@ I���ٿ�_�k&��@� ��4@������!?���*q�@^�dDR�ٿqS��h~�@�<�|&4@�O�BX�!?���{���@^�dDR�ٿqS��h~�@�<�|&4@�O�BX�!?���{���@^�dDR�ٿqS��h~�@�<�|&4@�O�BX�!?���{���@Qkɫ�ٿ�����@n�}��%4@YF�P��!?��v��@Qkɫ�ٿ�����@n�}��%4@YF�P��!?��v��@Qkɫ�ٿ�����@n�}��%4@YF�P��!?��v��@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@g�8�ٿ8[8���@�ZA�x4@b���M�!?:�D羕@�'�Q�ٿ��R�L��@*{9�!-4@�"��l�!?�:����@�'�Q�ٿ��R�L��@*{9�!-4@�"��l�!?�:����@�'�Q�ٿ��R�L��@*{9�!-4@�"��l�!?�:����@���KТٿ�����@���4@*q��]�!?s�� �@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�%-$��ٿ����<�@����4@�Ϫ�$�!?@U+�Z��@�B
G(�ٿ2߮�MS�@��oO74@:�0"6�!?(�rF���@�B
G(�ٿ2߮�MS�@��oO74@:�0"6�!?(�rF���@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@."�jO�ٿ�ҿM��@�����D4@�j6@�!?r� �@jW���ٿqO(����@ ��'wB4@�dn}f�!?ʋ�S�ʕ@jW���ٿqO(����@ ��'wB4@�dn}f�!?ʋ�S�ʕ@jW���ٿqO(����@ ��'wB4@�dn}f�!?ʋ�S�ʕ@jW���ٿqO(����@ ��'wB4@�dn}f�!?ʋ�S�ʕ@jW���ٿqO(����@ ��'wB4@�dn}f�!?ʋ�S�ʕ@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@��9Ɵٿ\����@�tp4��3@/�$甐!?�Q�'�@c��*�ٿzV����@!+),4@]�y���!?�Ry԰�@c��*�ٿzV����@!+),4@]�y���!?�Ry԰�@�����ٿV{���@:����3@�� m�!?r�I�cw�@�����ٿV{���@:����3@�� m�!?r�I�cw�@�����ٿV{���@:����3@�� m�!?r�I�cw�@�L�7P�ٿ�c����@���$4@4��MU�!?
a�2ٕ@�L�7P�ٿ�c����@���$4@4��MU�!?
a�2ٕ@�L�7P�ٿ�c����@���$4@4��MU�!?
a�2ٕ@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@a�!�K�ٿ�$�:��@�j��^)4@����+�!?/�ǡֽ�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@���9X�ٿG�u�@�T���34@:�w�!?��<�m�@��y�̝ٿ|�2��A�@6�d��$4@#�ڭ�!?)9XD��@��y�̝ٿ|�2��A�@6�d��$4@#�ڭ�!?)9XD��@��y�̝ٿ|�2��A�@6�d��$4@#�ڭ�!?)9XD��@�c?�*�ٿ2`��0��@>�)l4@��&$-�!?���Y�˕@�c?�*�ٿ2`��0��@>�)l4@��&$-�!?���Y�˕@�c?�*�ٿ2`��0��@>�)l4@��&$-�!?���Y�˕@�c?�*�ٿ2`��0��@>�)l4@��&$-�!?���Y�˕@�c?�*�ٿ2`��0��@>�)l4@��&$-�!?���Y�˕@��F$�ٿ�䭉QP�@w���
4@�"pPM�!?-��k��@��F$�ٿ�䭉QP�@w���
4@�"pPM�!?-��k��@s�ڹ�ٿɗ�Ze��@�b��3@
�?�!?��|;u��@4�1�ߚٿ�]�[���@��B��3@����A�!?��/��@�vƗ��ٿ�6=?��@������3@Y���!?����-��@`���A�ٿ���w��@|wG���3@<���M�!?_Qa�ʕ@`���A�ٿ���w��@|wG���3@<���M�!?_Qa�ʕ@��Мٿ�	Ǌ���@QVt�p!4@B�.�!?]�:���@�t��7�ٿ���|O�@����� 4@�=��S�!?(C�	��@�t��7�ٿ���|O�@����� 4@�=��S�!?(C�	��@�t��7�ٿ���|O�@����� 4@�=��S�!?(C�	��@yT).��ٿ�X U�R�@����4@�NG�!?]P��@�NF/�ٿ��T��@� ���14@�Bv���!? }84�@�NF/�ٿ��T��@� ���14@�Bv���!? }84�@K�:��ٿ)R�Q��@ �IX�4@�pVt�!?�`�Jx��@K�:��ٿ)R�Q��@ �IX�4@�pVt�!?�`�Jx��@K�:��ٿ)R�Q��@ �IX�4@�pVt�!?�`�Jx��@K�:��ٿ)R�Q��@ �IX�4@�pVt�!?�`�Jx��@��3�7�ٿs����@�Z�C4@oe>({�!?�����@1�J��ٿCG�"�(�@�0� �'4@��̎��!?���˕@1�J��ٿCG�"�(�@�0� �'4@��̎��!?���˕@1�J��ٿCG�"�(�@�0� �'4@��̎��!?���˕@1�J��ٿCG�"�(�@�0� �'4@��̎��!?���˕@1�J��ٿCG�"�(�@�0� �'4@��̎��!?���˕@�l���ٿ��8j��@o���E4@G�{4��!?���z�@�l���ٿ��8j��@o���E4@G�{4��!?���z�@;h_���ٿ���rm7�@G�|�e4@b˱E��!?}�X�$f�@�X	�y�ٿ���)Ҥ�@r�E�l4@Nu5b��!?���@�֕@�X	�y�ٿ���)Ҥ�@r�E�l4@Nu5b��!?���@�֕@�X	�y�ٿ���)Ҥ�@r�E�l4@Nu5b��!?���@�֕@Z:�T�ٿxYۍ���@��W��G4@�w���!?�5ΣQ��@Z:�T�ٿxYۍ���@��W��G4@�w���!?�5ΣQ��@Z:�T�ٿxYۍ���@��W��G4@�w���!?�5ΣQ��@Z:�T�ٿxYۍ���@��W��G4@�w���!?�5ΣQ��@Z:�T�ٿxYۍ���@��W��G4@�w���!?�5ΣQ��@���-��ٿ@�^��@�|{s$4@���r�!?=1U�F��@���-��ٿ@�^��@�|{s$4@���r�!?=1U�F��@���-��ٿ@�^��@�|{s$4@���r�!?=1U�F��@���-��ٿ@�^��@�|{s$4@���r�!?=1U�F��@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@�W�b�ٿ?����@�҂ua94@�1e�!?ph44���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@-O�{�ٿR����j�@����4@��u�!?�|V���@�#����ٿ�B��@;�zV�4@�y/z�!?Z��5!��@y����ٿ�S��i�@� 9I>4@o���q�!?
�y���@y����ٿ�S��i�@� 9I>4@o���q�!?
�y���@��I�/�ٿQ~�xD�@�z�ɼ34@�&+7�!?"�C��Õ@4(J	�ٿ2�2l��@#���~I4@��xr$�!?��J%�i�@4(J	�ٿ2�2l��@#���~I4@��xr$�!?��J%�i�@4(J	�ٿ2�2l��@#���~I4@��xr$�!?��J%�i�@ �8i�ٿ����.j�@5c��-4@�T�]\�!?G�O�ߕ@ �8i�ٿ����.j�@5c��-4@�T�]\�!?G�O�ߕ@ �8i�ٿ����.j�@5c��-4@�T�]\�!?G�O�ߕ@��	��ٿ����C�@�z�4@�bl�!?߀|�P{�@��	��ٿ����C�@�z�4@�bl�!?߀|�P{�@��	��ٿ����C�@�z�4@�bl�!?߀|�P{�@��	��ٿ����C�@�z�4@�bl�!?߀|�P{�@4��`˟ٿ!�$�`��@t)�I�3@�<�K�!?�7��Sr�@�I�Ԡٿ��g? ��@ ��/��3@��$F�!?6��Rkו@ɵ�O�ٿF&�n,�@��0��4@���E-�!?0*k��@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@}X"�ٿ�n����@:nS9�4@۝=�`�!?W䝻�0�@P��ٿ��6媀�@�RiC�<4@��t�D�!?넾�֕@�{����ٿU�zn�@&k�-4@K�a�-�!?[�3�Ǖ@V��t}�ٿY��|���@<�Y���3@S �&�!?�muO���@V��t}�ٿY��|���@<�Y���3@S �&�!?�muO���@V��t}�ٿY��|���@<�Y���3@S �&�!?�muO���@V��t}�ٿY��|���@<�Y���3@S �&�!?�muO���@V��t}�ٿY��|���@<�Y���3@S �&�!?�muO���@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@��i��ٿ4�z��2�@�7���4@��V!�!?I���ו@����#�ٿ�w9Z>��@��QT�M4@���/�!?��,��ӕ@����#�ٿ�w9Z>��@��QT�M4@���/�!?��,��ӕ@�9�)�ٿ�tO�>P�@n��@�3@�~R(.�!?��,��&�@�9�)�ٿ�tO�>P�@n��@�3@�~R(.�!?��,��&�@�9�)�ٿ�tO�>P�@n��@�3@�~R(.�!?��,��&�@���b��ٿ_�*���@��F}�4@^�q&�!?��;8g�@���b��ٿ_�*���@��F}�4@^�q&�!?��;8g�@���b��ٿ_�*���@��F}�4@^�q&�!?��;8g�@���b��ٿ_�*���@��F}�4@^�q&�!?��;8g�@���b��ٿ_�*���@��F}�4@^�q&�!?��;8g�@�U�͡ٿ>'՚�#�@_yyۀ�3@Q��6�!?)�q�,�@�U�͡ٿ>'՚�#�@_yyۀ�3@Q��6�!?)�q�,�@R@��q�ٿL�*rP�@��?��4@�b�* �!?��{�@��u��ٿ�Y�����@5�O\��3@c�X�u�!??�bu"ٕ@�6�X�ٿ�i>����@�S��?�3@��{�j�!?��h\���@�6�X�ٿ�i>����@�S��?�3@��{�j�!?��h\���@�6�X�ٿ�i>����@�S��?�3@��{�j�!?��h\���@՛����ٿ`q�q��@4ɦٙ3@�m57W�!?JF5VR��@f��Bלٿ[p��2�@��}yt�3@�_���!?���E��@f��Bלٿ[p��2�@��}yt�3@�_���!?���E��@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@rj�ۚٿ��d�4�@]�Ԛ��3@D@9�@�!?�R�cwڕ@pI��ٿ�����@&�US��3@�����!?�'�;�@pI��ٿ�����@&�US��3@�����!?�'�;�@pI��ٿ�����@&�US��3@�����!?�'�;�@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@���O�ٿ�7N��@ph�Z�3@j}�ǐ!?Jƙi���@5Ib�ٿLk��@���r5�3@�^����!?U?89��@5Ib�ٿLk��@���r5�3@�^����!?U?89��@5Ib�ٿLk��@���r5�3@�^����!?U?89��@5Ib�ٿLk��@���r5�3@�^����!?U?89��@D�lơٿuR����@�{
��3@��R��!?�6$�Fӕ@���Řٿ�ܼ��@~e����3@c�4俐!?)�I���@���Řٿ�ܼ��@~e����3@c�4俐!?)�I���@���Řٿ�ܼ��@~e����3@c�4俐!?)�I���@v#3��ٿ�J����@;�W��4@Y��Đ!?�В�l�@v#3��ٿ�J����@;�W��4@Y��Đ!?�В�l�@�t#{��ٿ���/7�@VBE�54@�ݚ��!?�j��@k�jX�ٿyҷ��k�@�4W�4@&ƌ��!?e��L���@k�jX�ٿyҷ��k�@�4W�4@&ƌ��!?e��L���@k�jX�ٿyҷ��k�@�4W�4@&ƌ��!?e��L���@�	~S�ٿ^�W
�@��>
�3@Yzu#%�!?^��mӕ@�	~S�ٿ^�W
�@��>
�3@Yzu#%�!?^��mӕ@��c��ٿ�������@c{�t��3@r~2-��!?\@��E�@��c��ٿ�������@c{�t��3@r~2-��!?\@��E�@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@r���s�ٿ?�j8�@����3@����i�!?=M=���@SߥK�ٿ�.d+q�@F��M�4@�#_��!?�Y���@�YG�ٿ�a���1�@�p��)4@}&/���!?.�c�@�YG�ٿ�a���1�@�p��)4@}&/���!?.�c�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@tc��E�ٿ��-͍�@yH4
�4@<U湐!?�_�~.�@��F�ߣٿ)� ��f�@�-���3@b�d���!?�n�J�@��F�ߣٿ)� ��f�@�-���3@b�d���!?�n�J�@
��a�ٿ'o|����@=����4@���� �!?'M��@
��a�ٿ'o|����@=����4@���� �!?'M��@
��a�ٿ'o|����@=����4@���� �!?'M��@F�ݥB�ٿ������@
��#4@*�8�!�!?���U�@F�ݥB�ٿ������@
��#4@*�8�!�!?���U�@F�ݥB�ٿ������@
��#4@*�8�!�!?���U�@F�ݥB�ٿ������@
��#4@*�8�!�!?���U�@�y�i��ٿÿc"x�@�����4@�Y�� �!?��A�6�@�y�i��ٿÿc"x�@�����4@�Y�� �!?��A�6�@�����ٿ`��G���@M����4@3d��!?�E+�1,�@5�[�ٿI:��+�@�����3@B�s]ُ!?�q�.G�@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@T�	�ˢٿ+�h�6�@�\�L�3@h+��!?S�[{� �@����o�ٿ)=��$�@ֳ�߅4@[�r<�!?�r��ey�@0���ٿLt����@�D�4@ 0�!?�:�{�~�@0���ٿLt����@�D�4@ 0�!?�:�{�~�@0���ٿLt����@�D�4@ 0�!?�:�{�~�@0���ٿLt����@�D�4@ 0�!?�:�{�~�@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@6ׇ	��ٿ{��T$�@q�+��/4@�\��*�!?�l��(��@���6�ٿ�S�$���@�#�^4@�� P�!?t�H�Y��@7e �M�ٿi�/���@%@�@4@��Z���!?�w���ϕ@c[gi�ٿ_@_u5�@mB��4@�s���!?$���ҕ@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@Iʺ��ٿF�G���@e�5��54@�̊�:�!?æ����@5�����ٿ�O,�q��@���^�74@�6)X5�!?Fƀ���@��+���ٿ���q��@���4@=嬧��!?����ǽ�@��+���ٿ���q��@���4@=嬧��!?����ǽ�@��+���ٿ���q��@���4@=嬧��!?����ǽ�@��+���ٿ���q��@���4@=嬧��!?����ǽ�@��+���ٿ���q��@���4@=嬧��!?����ǽ�@��+���ٿ���q��@���4@=嬧��!?����ǽ�@�vËĜٿww��3v�@t	L�3@֧�Ҭ�!?�3�4ݲ�@�vËĜٿww��3v�@t	L�3@֧�Ҭ�!?�3�4ݲ�@䋗�W�ٿ�~ �r��@Wb244@gQ�{�!?4��@����ٿ7|٤�@p�a��3@�����!?׶P0�@����ٿ7|٤�@p�a��3@�����!?׶P0�@����ٿ7|٤�@p�a��3@�����!?׶P0�@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@^��j�ٿ��=]���@5�9�4@k|�@��!?�/\���@8�M��ٿ�g���@�	^D�3@RR{��!?IJ� �&�@8�M��ٿ�g���@�	^D�3@RR{��!?IJ� �&�@8�M��ٿ�g���@�	^D�3@RR{��!?IJ� �&�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@�7ukA�ٿ�\Aە}�@+"�Mz�3@��m#Y�!?̃D��^�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@#�ٿ�7�7|.�@����[4@ȝ��5�!?f��]A.�@h�$�ٿ9�;����@8�Ї)4@g��!?jh>���@h�$�ٿ9�;����@8�Ї)4@g��!?jh>���@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@@��=��ٿ���$�@s��WC4@�C��Z�!?]��L̕@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@��O�g�ٿ'�%���@
^I[s4@�3�u�!?O*iq��@����ٿ(�����@�P��3@b&qz�!?���O��@����ٿ(�����@�P��3@b&qz�!?���O��@����ٿ(�����@�P��3@b&qz�!?���O��@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�J]j�ٿ%��@���hm�3@V{q��!?�.�ڕ@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�ѲfR�ٿ�>:�@�"G��3@�Jn��!?�$W���@�܃��ٿcycP@\�@L,[�(�3@N�0ݩ�!?v�]�f�@拙�ٿ6�F��@��0�4@|��:�!?/w��\�@拙�ٿ6�F��@��0�4@|��:�!?/w��\�@拙�ٿ6�F��@��0�4@|��:�!?/w��\�@拙�ٿ6�F��@��0�4@|��:�!?/w��\�@拙�ٿ6�F��@��0�4@|��:�!?/w��\�@@8�+��ٿ�X�����@[f���3@
q�%�!?�`TȨ�@@8�+��ٿ�X�����@[f���3@
q�%�!?�`TȨ�@@8�+��ٿ�X�����@[f���3@
q�%�!?�`TȨ�@ �H�+�ٿE�v���@}�tet�3@�v�0�!?�R�
���@ �H�+�ٿE�v���@}�tet�3@�v�0�!?�R�
���@ �H�+�ٿE�v���@}�tet�3@�v�0�!?�R�
���@O����ٿ����nR�@�wY��3@(l!k�!?��k,�@O����ٿ����nR�@�wY��3@(l!k�!?��k,�@O����ٿ����nR�@�wY��3@(l!k�!?��k,�@O����ٿ����nR�@�wY��3@(l!k�!?��k,�@O����ٿ����nR�@�wY��3@(l!k�!?��k,�@��5�ٿ6`q����@��6�3@��T� �!?��8ܰ-�@��.[^�ٿ��T�{�@�����3@9<����!?e2�GG)�@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@��e��ٿ�H]$�L�@�~��3@uuƒW�!?8�ߘ"��@�aX��ٿF�@a$�@�����3@I7f�W�!?�go�:��@�aX��ٿF�@a$�@�����3@I7f�W�!?�go�:��@�aX��ٿF�@a$�@�����3@I7f�W�!?�go�:��@󱻨��ٿ����(�@�dEqu�3@8�����!?0"��8�@󱻨��ٿ����(�@�dEqu�3@8�����!?0"��8�@@^��M�ٿ���Ҫ��@���V�3@x�� ͐!?���9��@@^��M�ٿ���Ҫ��@���V�3@x�� ͐!?���9��@�怨>�ٿ��)�U��@#�	!�4@#�|Ő!?㧘5��@�怨>�ٿ��)�U��@#�	!�4@#�|Ő!?㧘5��@�怨>�ٿ��)�U��@#�	!�4@#�|Ő!?㧘5��@� $��ٿ����+�@ޱ��<#4@� 'd�!?�:]f꩕@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@6��k�ٿgG�x�S�@��.4@Ze>�!?O(�&vĕ@��t�ٿ�38I*�@�wG��4@����!?9?*Aܕ@��t�ٿ�38I*�@�wG��4@����!?9?*Aܕ@��t�ٿ�38I*�@�wG��4@����!?9?*Aܕ@��t�ٿ�38I*�@�wG��4@����!?9?*Aܕ@��t�ٿ�38I*�@�wG��4@����!?9?*Aܕ@*�>�ٿ��Lϓ��@�*��b4@~E�3��!?z�;2��@*�>�ٿ��Lϓ��@�*��b4@~E�3��!?z�;2��@*�>�ٿ��Lϓ��@�*��b4@~E�3��!?z�;2��@*�>�ٿ��Lϓ��@�*��b4@~E�3��!?z�;2��@*�>�ٿ��Lϓ��@�*��b4@~E�3��!?z�;2��@�β�ٿ��S�a�@12��k4@l���ߐ!?�φ!^��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@�
4�>�ٿ���6C�@��i4@j�ъ��!?�*�L��@t�~�D�ٿ�u�4�@{I�B�'4@�N�*:�!?��n�(�@t�~�D�ٿ�u�4�@{I�B�'4@�N�*:�!?��n�(�@t�~�D�ٿ�u�4�@{I�B�'4@�N�*:�!?��n�(�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@�V��ٿ��h��@�9�Ay4@w�\�i�!??mGk=�@��ٿ�<K��@�x
��r4@7�d�*�!?�4F�(�@��ٿ�<K��@�x
��r4@7�d�*�!?�4F�(�@��ٿ�<K��@�x
��r4@7�d�*�!?�4F�(�@�|\�2�ٿ�["��T�@yj;q�&4@X%@?*�!?�1�@�/�@�|\�2�ٿ�["��T�@yj;q�&4@X%@?*�!?�1�@�/�@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@oƴ(��ٿ�������@�,j
c4@"-���!?j��]* �@H�l��ٿn������@�/�(4@��'�U�!?X����@H�l��ٿn������@�/�(4@��'�U�!?X����@H�l��ٿn������@�/�(4@��'�U�!?X����@H�l��ٿn������@�/�(4@��'�U�!?X����@H�l��ٿn������@�/�(4@��'�U�!?X����@H�l��ٿn������@�/�(4@��'�U�!?X����@�]R���ٿ-�:T���@���4@/�,�H�!?�KTJ�@�]R���ٿ-�:T���@���4@/�,�H�!?�KTJ�@�]R���ٿ-�:T���@���4@/�,�H�!?�KTJ�@���H�ٿ&�g4	��@ΈK���3@T+��J�!?�Ĝ�ҕ@���H�ٿ&�g4	��@ΈK���3@T+��J�!?�Ĝ�ҕ@���H�ٿ&�g4	��@ΈK���3@T+��J�!?�Ĝ�ҕ@�^%�3�ٿg��S�@Ӟ����3@�J�Yc�!?��1Gԕ@�^%�3�ٿg��S�@Ӟ����3@�J�Yc�!?��1Gԕ@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@T����ٿR�-��@�����3@�Ny$��!?tf�� ��@�幁�ٿe�ˌ1�@�����3@�E���!?d���ݕ@����ٿ	{�f=*�@\�h�{g4@q�%���!?	�M4�@Vh���ٿ�4����@)6n�JO4@���!?+K��@Vh���ٿ�4����@)6n�JO4@���!?+K��@Vh���ٿ�4����@)6n�JO4@���!?+K��@Vh���ٿ�4����@)6n�JO4@���!?+K��@�'�1,�ٿ��q���@'U�!G4@m�?��!?���A�&�@��8,�ٿ�m`�_�@=/��+4@��/�ߐ!?�T��&�@��8,�ٿ�m`�_�@=/��+4@��/�ߐ!?�T��&�@P{Ao��ٿ��&�d��@�0�4@ ���Ð!?�^�����@P{Ao��ٿ��&�d��@�0�4@ ���Ð!?�^�����@P{Ao��ٿ��&�d��@�0�4@ ���Ð!?�^�����@P{Ao��ٿ��&�d��@�0�4@ ���Ð!?�^�����@���E|�ٿ��GiE#�@�Y%�j�3@��1��!?�^Q��@���E|�ٿ��GiE#�@�Y%�j�3@��1��!?�^Q��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�A��ٿ�/�3�@��_�B�3@�:��ː!?_t��}��@�|�5��ٿ���zx�@�k�[4@��,�ɐ!?<���G�@�|�5��ٿ���zx�@�k�[4@��,�ɐ!?<���G�@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@=��`ڜٿ'"�h4��@������3@
��!?�������@���
��ٿ���yp�@����*�3@�o���!?q�,��P�@���
��ٿ���yp�@����*�3@�o���!?q�,��P�@���
��ٿ���yp�@����*�3@�o���!?q�,��P�@�7褿�ٿ��:	f�@m�n?�<4@�܋u��!?� L�J�@;��A�ٿ��:/G��@y����4@9�ęs�!?g���t�@;��A�ٿ��:/G��@y����4@9�ęs�!?g���t�@;��A�ٿ��:/G��@y����4@9�ęs�!?g���t�@;��A�ٿ��:/G��@y����4@9�ęs�!?g���t�@;��A�ٿ��:/G��@y����4@9�ęs�!?g���t�@��ǡ�ٿ�!50��@�ʿ�*4@�Hq@�!??gϢ]O�@��ǡ�ٿ�!50��@�ʿ�*4@�Hq@�!??gϢ]O�@��ǡ�ٿ�!50��@�ʿ�*4@�Hq@�!??gϢ]O�@�S�=�ٿ�3���@xŕ�94@|ΝgD�!?��g-��@�S�=�ٿ�3���@xŕ�94@|ΝgD�!?��g-��@�S�=�ٿ�3���@xŕ�94@|ΝgD�!?��g-��@�S�=�ٿ�3���@xŕ�94@|ΝgD�!?��g-��@�S�=�ٿ�3���@xŕ�94@|ΝgD�!?��g-��@��X;)�ٿ�N߲��@�j�7�c4@)�Q�A�!?<i����@P�ūܖٿaǡ���@����X4@�dh�J�!?u��eו@P�ūܖٿaǡ���@����X4@�dh�J�!?u��eו@P�ūܖٿaǡ���@����X4@�dh�J�!?u��eו@P�ūܖٿaǡ���@����X4@�dh�J�!?u��eו@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@�pU�ٿD`�%��@�&S��3@+�\�!?�P�8�d�@H�I�ٿo;x��'�@rƝv 4@��;���!?�h;����@H�I�ٿo;x��'�@rƝv 4@��;���!?�h;����@H�I�ٿo;x��'�@rƝv 4@��;���!?�h;����@H�I�ٿo;x��'�@rƝv 4@��;���!?�h;����@l��Šٿ�~�J�@[�Ŵ�+4@2}����!?-6O�O@l��Šٿ�~�J�@[�Ŵ�+4@2}����!?-6O�O@l��Šٿ�~�J�@[�Ŵ�+4@2}����!?-6O�O@��=�ٿ��$�1�@ 5:�3@�w-�|�!?�ј�˕@��=�ٿ��$�1�@ 5:�3@�w-�|�!?�ј�˕@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�`Z?;�ٿ��)%�@�h�4@�z^�N�!?o^5�H�@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@�X��ژٿd}#b�@�Į���3@12�b�!?�#����@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@+4� �ٿ������@� �{t�3@*�V�!?���f��@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@G����ٿ	�����@�+@aq24@�����!?1 w�ޕ@���.�ٿ-<����@2�8vM*4@�v�9�!?6�l;��@���.�ٿ-<����@2�8vM*4@�v�9�!?6�l;��@���.�ٿ-<����@2�8vM*4@�v�9�!?6�l;��@ĩ;T�ٿ>8Wd��@9%m_4@?G�b�!?��t��Е@ĩ;T�ٿ>8Wd��@9%m_4@?G�b�!?��t��Е@ĩ;T�ٿ>8Wd��@9%m_4@?G�b�!?��t��Е@�xz��ٿ����;"�@�;�'�V4@=+`4�!?X�Y��#�@�xz��ٿ����;"�@�;�'�V4@=+`4�!?X�Y��#�@��e\�ٿ���@����Aa4@&߂�A�!?pu���@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@y��eܖٿ�^�ĸ��@�����4@��o�7�!?�"cs�@���*�ٿ��EԌc�@O��;4@�mߙ�!?fT�Vޖ�@���*�ٿ��EԌc�@O��;4@�mߙ�!?fT�Vޖ�@�����ٿ�9�it8�@�\�.4@��˧Ő!?���-j�@%�Ñ�ٿ�B�f��@��s��4@3����!?g���q�@%�Ñ�ٿ�B�f��@��s��4@3����!?g���q�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@��.���ٿ.g�y���@|���(4@��h��!?7Ƨ3r)�@������ٿ|x닣��@�Q]�`�3@J��)�!?������@������ٿ|x닣��@�Q]�`�3@J��)�!?������@������ٿ|x닣��@�Q]�`�3@J��)�!?������@������ٿ|x닣��@�Q]�`�3@J��)�!?������@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@w!���ٿ���%ˣ�@�22�1,4@u_�5�!?���Hɕ@V��ŝٿY� Q���@����3@��x�{�!?�eC9tڕ@V��ŝٿY� Q���@����3@��x�{�!?�eC9tڕ@V��ŝٿY� Q���@����3@��x�{�!?�eC9tڕ@�Q���ٿ�|l~m:�@�5��14@� [�!?�(�ŕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@NW#��ٿ�
=����@��6�4@�|+���!?�-�Kʕ@ݕ���ٿoz�"�@y��;)"4@S�7�!?�z�R��@ݕ���ٿoz�"�@y��;)"4@S�7�!?�z�R��@ݕ���ٿoz�"�@y��;)"4@S�7�!?�z�R��@ݕ���ٿoz�"�@y��;)"4@S�7�!?�z�R��@���b�ٿ:Ik��+�@zY���*4@&(9�-�!?�A�\�ѕ@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@!m�r�ٿ���@Q	�2 4@E{Շ�!?M@S'�@����Z�ٿ��r}/��@{����3@zq�5@�!?����@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@��0�"�ٿF�y����@�Y�"�3@0v���!?p��l-@�@q�L�p�ٿ�h4p�@��ey�3@��RK�!??&���@q�L�p�ٿ�h4p�@��ey�3@��RK�!??&���@q�L�p�ٿ�h4p�@��ey�3@��RK�!??&���@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��|*ͤٿ���-�@���+��3@ߴ�n�!?�-ͷ&�@��e�Ĥٿ�7�9]�@_r8�4@/�d���!?���J�ϕ@��e�Ĥٿ�7�9]�@_r8�4@/�d���!?���J�ϕ@��e�Ĥٿ�7�9]�@_r8�4@/�d���!?���J�ϕ@��e�Ĥٿ�7�9]�@_r8�4@/�d���!?���J�ϕ@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@;-�p �ٿ�~da��@�JS�%�3@F�9dΐ!?S��('�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@��P�ٿ衑�?(�@�@��:4@Y����!?'r�G^�@�U ���ٿ��6%�|�@����54@|�!?_	w�v�@�U ���ٿ��6%�|�@����54@|�!?_	w�v�@��'�ʠٿ�Ӥa�w�@�m�F�74@;�:�|�!?by��E�@��'�ʠٿ�Ӥa�w�@�m�F�74@;�:�|�!?by��E�@7�+� �ٿ[�
���@T50��4@i�÷��!?p��FL��@7�+� �ٿ[�
���@T50��4@i�÷��!?p��FL��@(��&�ٿ3\�~��@dP_�!4@k칐�!?�	�H;ȕ@n��,j�ٿ�p��.P�@�_�N4@�<���!?��z�@Wܵ�r�ٿ��]���@|�ŵ4@��q�K�!?��5�V�@Wܵ�r�ٿ��]���@|�ŵ4@��q�K�!?��5�V�@Wܵ�r�ٿ��]���@|�ŵ4@��q�K�!?��5�V�@Wܵ�r�ٿ��]���@|�ŵ4@��q�K�!?��5�V�@Y�-�ݙٿ��yg�@�6N� 4@�=�x(�!?�>�l��@Y�-�ݙٿ��yg�@�6N� 4@�=�x(�!?�>�l��@Y�-�ݙٿ��yg�@�6N� 4@�=�x(�!?�>�l��@Y�-�ݙٿ��yg�@�6N� 4@�=�x(�!?�>�l��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@:H��A�ٿ��A�U#�@+��r�	4@`o���!?���Z��@%z�ٿg�*$��@~}I�4@���j	�!?��XS%ݕ@%z�ٿg�*$��@~}I�4@���j	�!?��XS%ݕ@����ٿ�/Kaa�@"
�@�4@)�=t�!?�p���@����ٿ�/Kaa�@"
�@�4@)�=t�!?�p���@y���ٿȊ��W��@�{�� "4@6J��p�!?�CAו@y���ٿȊ��W��@�{�� "4@6J��p�!?�CAו@y���ٿȊ��W��@�{�� "4@6J��p�!?�CAו@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@�l���ٿ���}&/�@���Y94@�ޝ�Q�!?�F��Iؕ@sF4\n�ٿ���+p��@��l��4@n���!?�Z�N݉�@;�:V)�ٿ���`���@��p�3�3@\-�i�!?�[�l鬕@;�:V)�ٿ���`���@��p�3�3@\-�i�!?�[�l鬕@�s?A�ٿ�/����@�Ҁ�N<4@��R9�!?E^����@�s?A�ٿ�/����@�Ҁ�N<4@��R9�!?E^����@�s?A�ٿ�/����@�Ҁ�N<4@��R9�!?E^����@�s?A�ٿ�/����@�Ҁ�N<4@��R9�!?E^����@�s?A�ٿ�/����@�Ҁ�N<4@��R9�!?E^����@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�ۇI�ٿF��-��@By��?4@.o�>�!?�:Z0�4�@�I�Q�ٿ|����@Ȉ��@%4@��Pt�!?��n���@�I�Q�ٿ|����@Ȉ��@%4@��Pt�!?��n���@����ٿ6�����@V�IA&/4@1�sß�!?�#,��ڕ@����ٿ6�����@V�IA&/4@1�sß�!?�#,��ڕ@����ٿ6�����@V�IA&/4@1�sß�!?�#,��ڕ@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�5�㐝ٿA|�?_�@Ec��+4@�}�!??s����@�� ��ٿ�mz�A9�@���2�-4@�7��c�!?D�v��ȕ@�� ��ٿ�mz�A9�@���2�-4@�7��c�!?D�v��ȕ@�� ��ٿ�mz�A9�@���2�-4@�7��c�!?D�v��ȕ@�� ��ٿ�mz�A9�@���2�-4@�7��c�!?D�v��ȕ@� ��ٿ� �m(�@S>�JX4@I�⩐!?�x���@� ��ٿ� �m(�@S>�JX4@I�⩐!?�x���@� ��ٿ� �m(�@S>�JX4@I�⩐!?�x���@� ��ٿ� �m(�@S>�JX4@I�⩐!?�x���@� ��ٿ� �m(�@S>�JX4@I�⩐!?�x���@��"�ٿ�^�1�>�@�@Y�=�3@���H�!?qz)���@��"�ٿ�^�1�>�@�@Y�=�3@���H�!?qz)���@��"�ٿ�^�1�>�@�@Y�=�3@���H�!?qz)���@Jr>��ٿ�n"]��@��a�p�3@z%�>�!?��g�x�@Jr>��ٿ�n"]��@��a�p�3@z%�>�!?��g�x�@).è�ٿ�C��t+�@V�o
4@�m����!?.�^d2�@).è�ٿ�C��t+�@V�o
4@�m����!?.�^d2�@��BC�ٿM����@�0bӺ�3@sf�t�!?!���nO�@;���٣ٿo�a��@�c,�`�3@3q�WO�!?�̋_u�@_\��ٿ�5�z���@��� �3@�Ў�h�!?_�Dń��@_\��ٿ�5�z���@��� �3@�Ў�h�!?_�Dń��@_\��ٿ�5�z���@��� �3@�Ў�h�!?_�Dń��@1�*G�ٿf�.+��@���V��3@Nh�*%�!?��L9���@�gf��ٿ��lx�^�@���^�3@�
A"�!?��0�1�@�gf��ٿ��lx�^�@���^�3@�
A"�!?��0�1�@G�޳��ٿm!��3�@�='�4@���Ώ!?�&�/ڎ�@G�޳��ٿm!��3�@�='�4@���Ώ!?�&�/ڎ�@G�޳��ٿm!��3�@�='�4@���Ώ!?�&�/ڎ�@G�޳��ٿm!��3�@�='�4@���Ώ!?�&�/ڎ�@����6�ٿA��AZ��@�~^��3@B�r�=�!?h�?�v|�@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@�a(��ٿP�N���@�WҐ�3@)���i�!?Y��L:��@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@���T�ٿ%H�?�@Ȱa�Q74@���o�!?�#��^%�@6�>��ٿ:Q��}�@��w��$4@C�j�!?�h�d#.�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@�O�ٿ��1��@�� �C4@+��8[�!?1E�9�5�@Buf�E�ٿP�Rk�)�@�|��`4@4L�F�!?/��gϕ@Buf�E�ٿP�Rk�)�@�|��`4@4L�F�!?/��gϕ@Buf�E�ٿP�Rk�)�@�|��`4@4L�F�!?/��gϕ@��$̈�ٿ=���@�҅x�	4@��3�T�!?_�T�@��$̈�ٿ=���@�҅x�	4@��3�T�!?_�T�@��$̈�ٿ=���@�҅x�	4@��3�T�!?_�T�@?h����ٿ�${"���@]-��@4@��x3�!?)z<@Jҕ@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@@���c�ٿ�[�8�@dՖ�)
4@C�>�D�!?����[�@���u��ٿoN�&���@���V!4@	�b�c�!?^�p���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@�+�8=�ٿJ6��@��x�?4@��T�!?V�e���@PL�ܣٿ���Z�@2K�74@A>�
`�!?4@f��ȕ@PL�ܣٿ���Z�@2K�74@A>�
`�!?4@f��ȕ@PL�ܣٿ���Z�@2K�74@A>�
`�!?4@f��ȕ@PL�ܣٿ���Z�@2K�74@A>�
`�!?4@f��ȕ@��ٿcXs����@�0px&4@�9���!?�m{ ��@��ٿcXs����@�0px&4@�9���!?�m{ ��@��ٿcXs����@�0px&4@�9���!?�m{ ��@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@�����ٿ$)r8��@�	(9^.4@�G�j�!?�]��Nŕ@v��R�ٿ�B����@����4@i�C�!?����}�@v��R�ٿ�B����@����4@i�C�!?����}�@dc�Eϛٿ0�A��@�T�#4@����!?��U��q�@dc�Eϛٿ0�A��@�T�#4@����!?��U��q�@dc�Eϛٿ0�A��@�T�#4@����!?��U��q�@.-z��ٿh��ȴ2�@�ze �3@tYm�[�!?�O[�b�@�IK�ٿ���e��@/r�g@�3@T��Z{�!?%_�N]�@�IK�ٿ���e��@/r�g@�3@T��Z{�!?%_�N]�@�IK�ٿ���e��@/r�g@�3@T��Z{�!?%_�N]�@�s{��ٿF�����@��|��3@7ס�N�!?1�>M͈�@�s{��ٿF�����@��|��3@7ס�N�!?1�>M͈�@�p�Y��ٿ?������@��RL�3@��+7X�!?}2sx��@�p�Y��ٿ?������@��RL�3@��+7X�!?}2sx��@�p�Y��ٿ?������@��RL�3@��+7X�!?}2sx��@�p�Y��ٿ?������@��RL�3@��+7X�!?}2sx��@�[���ٿ��}����@-=��I�3@�=�p�!?���1���@�[���ٿ��}����@-=��I�3@�=�p�!?���1���@�[���ٿ��}����@-=��I�3@�=�p�!?���1���@�[���ٿ��}����@-=��I�3@�=�p�!?���1���@�[���ٿ��}����@-=��I�3@�=�p�!?���1���@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@���Gԝٿ~yQ#�@�H���3@k�����!?<��0��@��˓�ٿ#�n����@�5�X�3@8�hPz�!?0/��;l�@��˓�ٿ#�n����@�5�X�3@8�hPz�!?0/��;l�@��˓�ٿ#�n����@�5�X�3@8�hPz�!?0/��;l�@��˓�ٿ#�n����@�5�X�3@8�hPz�!?0/��;l�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@#Fq�q�ٿ�D ���@���d��3@�]�I�!?�<�]�@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@��ן�ٿu�Cy�S�@Q�U�y�3@�^R�w�!?�)���@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@ ���:�ٿ�g猈N�@)g*��3@�A_��!?�!;�@l�?<�ٿ�vp��@P��(4@�1.�K�!?/t_�rٕ@��H��ٿW+am�s�@xTp�[4@��*���!?�v�1q�@ɋ����ٿm��;��@K��d+&4@���&�!?�;I�@ɋ����ٿm��;��@K��d+&4@���&�!?�;I�@ɋ����ٿm��;��@K��d+&4@���&�!?�;I�@ɋ����ٿm��;��@K��d+&4@���&�!?�;I�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@r�ٿ�ozރ�@��
��E4@ȹ��w�!?C�j�@d��]�ٿ��SY�@�����n4@�ʘ�W�!?�x��ɕ@d��]�ٿ��SY�@�����n4@�ʘ�W�!?�x��ɕ@�b���ٿ?�ٵ��@�U�x4@���̔�!?�yS$��@�b���ٿ?�ٵ��@�U�x4@���̔�!?�yS$��@�b���ٿ?�ٵ��@�U�x4@���̔�!?�yS$��@�D72�ٿ�����s�@��T_4@^?��s�!?	�jĕ@�D72�ٿ�����s�@��T_4@^?��s�!?	�jĕ@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@��n娟ٿ��u��@2Ԩ"� 4@�VE��!?b����@¥:d��ٿ(�c��k�@����3@�P��C�!?�~�����@¥:d��ٿ(�c��k�@����3@�P��C�!?�~�����@¥:d��ٿ(�c��k�@����3@�P��C�!?�~�����@¥:d��ٿ(�c��k�@����3@�P��C�!?�~�����@¥:d��ٿ(�c��k�@����3@�P��C�!?�~�����@�"�ۘٿ�z�X^��@��.iE4@ׄ#0�!?L���i�@�-X�ܖٿy��
D�@<é[�H4@�(�!?�Ç�ƕ@�-X�ܖٿy��
D�@<é[�H4@�(�!?�Ç�ƕ@c�1���ٿy+��`$�@A¬�/4@��H�!?�l�aE�@�^";N�ٿ7/��n�@A�M�!?4@|����!?�m���@�^";N�ٿ7/��n�@A�M�!?4@|����!?�m���@
c�`J�ٿ9�u2�@rH�� 4@�_ q�!?!��d�q�@
c�`J�ٿ9�u2�@rH�� 4@�_ q�!?!��d�q�@
c�`J�ٿ9�u2�@rH�� 4@�_ q�!?!��d�q�@
c�`J�ٿ9�u2�@rH�� 4@�_ q�!?!��d�q�@h�)�ٿv*Dc)�@�X�,a4@�}��.�!?'�g�L�@ޜq��ٿ&���y�@<��7�P4@���:P�!?�S-���@ޜq��ٿ&���y�@<��7�P4@���:P�!?�S-���@��O�G�ٿ�M 䣰�@u�?B4@~�@r�!?=�ި��@��O�G�ٿ�M 䣰�@u�?B4@~�@r�!?=�ި��@��O�G�ٿ�M 䣰�@u�?B4@~�@r�!?=�ި��@��O�G�ٿ�M 䣰�@u�?B4@~�@r�!?=�ި��@��O�G�ٿ�M 䣰�@u�?B4@~�@r�!?=�ި��@c/=�C�ٿ���J\�@�$�$*4@���.|�!?��qI���@c/=�C�ٿ���J\�@�$�$*4@���.|�!?��qI���@�Թɢٿ�I�5?��@/�g�q$4@F�s�$�!?��wPٶ�@�Թɢٿ�I�5?��@/�g�q$4@F�s�$�!?��wPٶ�@rf�Պ�ٿ��%e��@ؽ�O�3@ݐ�.�!?��)ȗ�@rf�Պ�ٿ��%e��@ؽ�O�3@ݐ�.�!?��)ȗ�@rf�Պ�ٿ��%e��@ؽ�O�3@ݐ�.�!?��)ȗ�@��Rk,�ٿ9��$��@����3@�Q�n1�!?[�]�`�@��Rk,�ٿ9��$��@����3@�Q�n1�!?[�]�`�@��Rk,�ٿ9��$��@����3@�Q�n1�!?[�]�`�@q[��ٿ�
T���@È�S�3@TD�&�!?�4��^�@�X����ٿ�t]V��@�Nv���3@a�w�!?�T�*9��@�X����ٿ�t]V��@�Nv���3@a�w�!?�T�*9��@�X����ٿ�t]V��@�Nv���3@a�w�!?�T�*9��@7֦xj�ٿ��7�H[�@�lT�?�3@���T(�!?3({��@7֦xj�ٿ��7�H[�@�lT�?�3@���T(�!?3({��@7֦xj�ٿ��7�H[�@�lT�?�3@���T(�!?3({��@7֦xj�ٿ��7�H[�@�lT�?�3@���T(�!?3({��@����ٿ��Q?�@���t�3@����E�!?����٦�@����ٿ��Q?�@���t�3@����E�!?����٦�@����ٿ��Q?�@���t�3@����E�!?����٦�@����ٿ��Q?�@���t�3@����E�!?����٦�@����ٿ��Q?�@���t�3@����E�!?����٦�@��0�ٿ��-E��@˧Ԏ��3@���C�!?NEj%Fٕ@��0�ٿ��-E��@˧Ԏ��3@���C�!?NEj%Fٕ@��0�ٿ��-E��@˧Ԏ��3@���C�!?NEj%Fٕ@��0�ٿ��-E��@˧Ԏ��3@���C�!?NEj%Fٕ@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@[��r{�ٿ�^7�gJ�@����4@�!ZDs�!?=!�7r�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@�ӄ�M�ٿ�Ag��@�	�T"4@��Ud�!?�ZFǢ�@%%R�ٿG'�1�@R*u4@]�M�i�!?�J���@%%R�ٿG'�1�@R*u4@]�M�i�!?�J���@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@����ٿ��2b�c�@K�����3@s�!�{�!?.2
��U�@LaU&�ٿ�`]�VK�@}�,^�3@M���k�!?P�
�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@�@� ��ٿ��zp7��@c&�r@<4@&�*C��!?x���:�@a�(m�ٿ�1��@p+P�+4@�m��	�!?tmz��ݕ@-���Z�ٿ�S�����@5��B4@z|z&M�!?2�����@���T(�ٿ:��Ź��@+M�Z4@�w�>��!?�K~R]{�@���T(�ٿ:��Ź��@+M�Z4@�w�>��!?�K~R]{�@���T(�ٿ:��Ź��@+M�Z4@�w�>��!?�K~R]{�@���T(�ٿ:��Ź��@+M�Z4@�w�>��!?�K~R]{�@-�q;՝ٿ���Y��@5υ�R4@�1UTI�!?<-O�>�@-�q;՝ٿ���Y��@5υ�R4@�1UTI�!?<-O�>�@-�q;՝ٿ���Y��@5υ�R4@�1UTI�!?<-O�>�@-�q;՝ٿ���Y��@5υ�R4@�1UTI�!?<-O�>�@-�q;՝ٿ���Y��@5υ�R4@�1UTI�!?<-O�>�@�?�F��ٿ��H��@U����n4@�G�$t�!?ӘR2���@�?�F��ٿ��H��@U����n4@�G�$t�!?ӘR2���@�?�F��ٿ��H��@U����n4@�G�$t�!?ӘR2���@�f�'M�ٿ��.Uz(�@���N�H4@A�'|�!?���~��@�f�'M�ٿ��.Uz(�@���N�H4@A�'|�!?���~��@�f�'M�ٿ��.Uz(�@���N�H4@A�'|�!?���~��@�f�'M�ٿ��.Uz(�@���N�H4@A�'|�!?���~��@�Ɨg��ٿ���S��@��}�=*4@H�fj�!?t��N�2�@���#��ٿO><(��@���k� 4@�z���!?^#%�@���#��ٿO><(��@���k� 4@�z���!?^#%�@�0�n�ٿ�T�R�@� �c�3@5�*���!?-%�yrZ�@�0�n�ٿ�T�R�@� �c�3@5�*���!?-%�yrZ�@�0�n�ٿ�T�R�@� �c�3@5�*���!?-%�yrZ�@�.�I�ٿg��-8Z�@���FD�3@<���z�!?Bk���p�@�.�I�ٿg��-8Z�@���FD�3@<���z�!?Bk���p�@$d7堜ٿ��Ŵ��@��+3��3@n����!?�#��@$d7堜ٿ��Ŵ��@��+3��3@n����!?�#��@.�T^�ٿC͔���@7��9��3@6�Z��!?����ѕ@�����ٿ�s"ܢ��@�zo 4@
^��!?��;:0�@�����ٿ�s"ܢ��@�zo 4@
^��!?��;:0�@�����ٿ�s"ܢ��@�zo 4@
^��!?��;:0�@�����ٿ�s"ܢ��@�zo 4@
^��!?��;:0�@�����ٿ�s"ܢ��@�zo 4@
^��!?��;:0�@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@�˯B��ٿ���1�.�@�"LAC4@�{󔘐!?3~���̕@b�M�ٿ'0��K�@(��g4@�,��>�!?�D�;��@b�M�ٿ'0��K�@(��g4@�,��>�!?�D�;��@b�M�ٿ'0��K�@(��g4@�,��>�!?�D�;��@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@�;�Q�ٿ(��f��@ĝb�
4@ZeoI�!?�@/*ו@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@8���ΚٿM�!vu[�@�r�7j�3@�ܞj�!?go�dL��@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@=m�F5�ٿ�*�O�^�@9� U)4@�H0s�!?��(��ٕ@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@��Wج�ٿ��P�@/��Q4@"n�h�!?Tw_�{��@�ۆ�:�ٿ��Ό5�@U'X7>^4@��l�!?�c�V�@�ۆ�:�ٿ��Ό5�@U'X7>^4@��l�!?�c�V�@�ۆ�:�ٿ��Ό5�@U'X7>^4@��l�!?�c�V�@�ۆ�:�ٿ��Ό5�@U'X7>^4@��l�!?�c�V�@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@���ٿ��i����@3V�F�4@�ʊ���!?�/�鶕@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@zDqr�ٿ�R����@�ޑ8,%4@����y�!?M����@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@�0�QҠٿ"ڏ�B�@��Tq�4@�~qr2�!?Iay��ܕ@A+�ٿ�����@�7?ٗ�3@����!?I�a����@A+�ٿ�����@�7?ٗ�3@����!?I�a����@A+�ٿ�����@�7?ٗ�3@����!?I�a����@A+�ٿ�����@�7?ٗ�3@����!?I�a����@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@ƞ[>�ٿq�W�@��5�3�3@|�7��!?<9:���@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@���3�ٿ=�$���@�5���4@61��k�!?\#�t�@XU����ٿ�_�tm�@��TxN4@0,�!?� ���@��?!ɣٿ�mY��@���w�4@ٞ�0�!?ӵq��@��?!ɣٿ�mY��@���w�4@ٞ�0�!?ӵq��@��?!ɣٿ�mY��@���w�4@ٞ�0�!?ӵq��@��?!ɣٿ�mY��@���w�4@ٞ�0�!?ӵq��@��?!ɣٿ�mY��@���w�4@ٞ�0�!?ӵq��@>�+y(�ٿ�yYc�@�l�'4@�-;P�!?bh���.�@S&	�ٿW&�s[�@J�kH�!4@���茐!?�~��p��@S&	�ٿW&�s[�@J�kH�!4@���茐!?�~��p��@3%g��ٿ��*ȱ��@����04@dC?���!?��S3b��@3%g��ٿ��*ȱ��@����04@dC?���!?��S3b��@��<N�ٿ�x���@0-˨4@ߌr��!?��0�m�@��<N�ٿ�x���@0-˨4@ߌr��!?��0�m�@��<N�ٿ�x���@0-˨4@ߌr��!?��0�m�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@�~K��ٿz'n���@���yY%4@|�\�!?n���:�@]�z�ڞٿU�ɗXr�@`�BH4@X�_�!?ǚ3�l��@]�z�ڞٿU�ɗXr�@`�BH4@X�_�!?ǚ3�l��@]�z�ڞٿU�ɗXr�@`�BH4@X�_�!?ǚ3�l��@]�z�ڞٿU�ɗXr�@`�BH4@X�_�!?ǚ3�l��@�3�
�ٿ�{��@.ȣw�4@���%^�!?H�� ۉ�@�3�
�ٿ�{��@.ȣw�4@���%^�!?H�� ۉ�@�3�
�ٿ�{��@.ȣw�4@���%^�!?H�� ۉ�@�3�
�ٿ�{��@.ȣw�4@���%^�!?H�� ۉ�@�3�
�ٿ�{��@.ȣw�4@���%^�!?H�� ۉ�@z�6q�ٿ/�q��@�V��Q4@��e�!?h;�wΕ@z�6q�ٿ/�q��@�V��Q4@��e�!?h;�wΕ@z�6q�ٿ/�q��@�V��Q4@��e�!?h;�wΕ@z�6q�ٿ/�q��@�V��Q4@��e�!?h;�wΕ@z�6q�ٿ/�q��@�V��Q4@��e�!?h;�wΕ@��R��ٿ����m��@�%%[44@��}2�!?@�"ɕ@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��D��ٿ�N����@��^�:64@'!1��!?@�Y�^@��M�z�ٿ�h����@v�)�4@��|�%�!?(����@��M�z�ٿ�h����@v�)�4@��|�%�!?(����@��M�z�ٿ�h����@v�)�4@��|�%�!?(����@��M�z�ٿ�h����@v�)�4@��|�%�!?(����@��M�z�ٿ�h����@v�)�4@��|�%�!?(����@�Xs��ٿ�r�p���@���&(�3@��#��!?z�,�pЕ@�Xs��ٿ�r�p���@���&(�3@��#��!?z�,�pЕ@�Xs��ٿ�r�p���@���&(�3@��#��!?z�,�pЕ@�Xs��ٿ�r�p���@���&(�3@��#��!?z�,�pЕ@�*䁋�ٿJ��E2q�@p�B��3@���w�!?�Ye8��@�*䁋�ٿJ��E2q�@p�B��3@���w�!?�Ye8��@��K=�ٿ捚���@�+l6��3@���^�!?\��5Fx�@��K=�ٿ捚���@�+l6��3@���^�!?\��5Fx�@���/��ٿ�U\�;�@��q�3@�4׋�!?-�m3��@Ѕ��j�ٿY��.��@�¢�G�3@�� ���!?�%�~[ŕ@Ѕ��j�ٿY��.��@�¢�G�3@�� ���!?�%�~[ŕ@3�1Z�ٿ�Y�^r�@ƣ���P4@��Ҏ�!?"�`d1�@3�1Z�ٿ�Y�^r�@ƣ���P4@��Ҏ�!?"�`d1�@3�1Z�ٿ�Y�^r�@ƣ���P4@��Ҏ�!?"�`d1�@3�1Z�ٿ�Y�^r�@ƣ���P4@��Ҏ�!?"�`d1�@3�1Z�ٿ�Y�^r�@ƣ���P4@��Ҏ�!?"�`d1�@�!��8�ٿ�p���@���윂4@#ȫ�(�!?���g�5�@D����ٿef�&���@{ŀ[��3@��	0�!?��*~�ٕ@D����ٿef�&���@{ŀ[��3@��	0�!?��*~�ٕ@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�[k6٤ٿ�U�+��@��#�3@\Sb�A�!?��ʓ���@�Bð�ٿ��)���@م���4@��c띐!?ZRY?W�@�Bð�ٿ��)���@م���4@��c띐!?ZRY?W�@�Bð�ٿ��)���@م���4@��c띐!?ZRY?W�@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@W(�OΝٿ��-���@C���84@z5���!?e�{�G��@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@h:�7�ٿƃB���@��rv�4@��q�!?1��c�@s5�Sm�ٿ92�mr�@���
4@��i�!?�dJI'�@s5�Sm�ٿ92�mr�@���
4@��i�!?�dJI'�@s5�Sm�ٿ92�mr�@���
4@��i�!?�dJI'�@u3���ٿ�$����@�E��I4@�*�f�!?@U@��f�@]	�.�ٿ�C1���@M@�B�4@��A�!?�[�a5��@]	�.�ٿ�C1���@M@�B�4@��A�!?�[�a5��@]	�.�ٿ�C1���@M@�B�4@��A�!?�[�a5��@t� 2Ơٿ ����@� �>�4@�^#��!?�6	R(�@t� 2Ơٿ ����@� �>�4@�^#��!?�6	R(�@t� 2Ơٿ ����@� �>�4@�^#��!?�6	R(�@�U��K�ٿ�Lj�;�@�4@�#�g/�!?R�MN��@�U��K�ٿ�Lj�;�@�4@�#�g/�!?R�MN��@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@qי�R�ٿk�R���@]��߁K4@nw9�:�!?2���89�@�]���ٿ����i�@��0j4@�ޜI�!?�ݽ�`�@�]���ٿ����i�@��0j4@�ޜI�!?�ݽ�`�@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@�Y���ٿy-#1-��@�-�L4@ի�'�!?�$w��@I_���ٿ�*�*Q��@>8aTB4@��E�s�!?��,���@I_���ٿ�*�*Q��@>8aTB4@��E�s�!?��,���@I_���ٿ�*�*Q��@>8aTB4@��E�s�!?��,���@I_���ٿ�*�*Q��@>8aTB4@��E�s�!?��,���@��Ꮌ�ٿ��^4��@��]c�4@4^���!?cG��ܕ@��Ꮌ�ٿ��^4��@��]c�4@4^���!?cG��ܕ@��Ꮌ�ٿ��^4��@��]c�4@4^���!?cG��ܕ@��Ꮌ�ٿ��^4��@��]c�4@4^���!?cG��ܕ@	Ă'
�ٿB��U�]�@54�.4@��}r>�!?��5?��@	Ă'
�ٿB��U�]�@54�.4@��}r>�!?��5?��@	Ă'
�ٿB��U�]�@54�.4@��}r>�!?��5?��@	Ă'
�ٿB��U�]�@54�.4@��}r>�!?��5?��@	Ă'
�ٿB��U�]�@54�.4@��}r>�!?��5?��@�?�a�ٿ��n G�@��F��3@��9�!?1
����@�?�a�ٿ��n G�@��F��3@��9�!?1
����@�?�a�ٿ��n G�@��F��3@��9�!?1
����@�?�a�ٿ��n G�@��F��3@��9�!?1
����@�?�a�ٿ��n G�@��F��3@��9�!?1
����@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@�*���ٿ�֨�f�@z��Y��3@؋rW�!?��s2=�@P�`�ٿr�[���@=+BK*�3@��:�!?��5��]�@P�`�ٿr�[���@=+BK*�3@��:�!?��5��]�@�d�H��ٿ,.��U�@a��%4@�zQ�e�!?�o�~���@�d�H��ٿ,.��U�@a��%4@�zQ�e�!?�o�~���@Ū�o�ٿ??�HnZ�@I�)�:84@ׁNUp�!?���r�6�@L�\-֗ٿ�͑����@�
nh.4@gVO�p�!?>3�z;E�@L�\-֗ٿ�͑����@�
nh.4@gVO�p�!?>3�z;E�@L�\-֗ٿ�͑����@�
nh.4@gVO�p�!?>3�z;E�@L�\-֗ٿ�͑����@�
nh.4@gVO�p�!?>3�z;E�@e�p�њٿ1�%g��@��:z14@��TU�!?`E]ưp�@�J�ٿ��ݼ��@�DW�NX4@H�0�d�!?Q��N9�@�J�ٿ��ݼ��@�DW�NX4@H�0�d�!?Q��N9�@�J�ٿ��ݼ��@�DW�NX4@H�0�d�!?Q��N9�@��0��ٿù��
�@l'���3@��H�4�!?K"�N��@��0��ٿù��
�@l'���3@��H�4�!?K"�N��@UmK感ٿS}���@����4@2ɻg�!?��`+���@UmK感ٿS}���@����4@2ɻg�!?��`+���@BUXw(�ٿP%��"L�@&"�:��3@���S�!?3��Z��@���ٿ�/J��Z�@�E4@��K�S�!?�f5�9��@���ٿ�/J��Z�@�E4@��K�S�!?�f5�9��@�T����ٿC^?���@qͿ���3@C���/�!?�iV�G��@�T����ٿC^?���@qͿ���3@C���/�!?�iV�G��@�T����ٿC^?���@qͿ���3@C���/�!?�iV�G��@�T����ٿC^?���@qͿ���3@C���/�!?�iV�G��@�T����ٿC^?���@qͿ���3@C���/�!?�iV�G��@�(�k�ٿ��X	��@�W��3@�X��1�!?�s3iCI�@�(�k�ٿ��X	��@�W��3@�X��1�!?�s3iCI�@�(�k�ٿ��X	��@�W��3@�X��1�!?�s3iCI�@�(�k�ٿ��X	��@�W��3@�X��1�!?�s3iCI�@@�ܦ��ٿ ��tA�@hf�rf�3@t�ؘ�!?���wP�@@�ܦ��ٿ ��tA�@hf�rf�3@t�ؘ�!?���wP�@A_h��ٿH��E���@zM�n=4@;
�+�!?t/�e!ו@A_h��ٿH��E���@zM�n=4@;
�+�!?t/�e!ו@DՐڣٿDf{�}�@�d�u4@�)r2�!?.������@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@��&��ٿ�H��c��@��c)DF4@neX��!?MO!=u��@���Չ�ٿ��]C���@�x*�A4@� ��!?YV�+1l�@���Չ�ٿ��]C���@�x*�A4@� ��!?YV�+1l�@���Չ�ٿ��]C���@�x*�A4@� ��!?YV�+1l�@���Չ�ٿ��]C���@�x*�A4@� ��!?YV�+1l�@���Չ�ٿ��]C���@�x*�A4@� ��!?YV�+1l�@��f���ٿOʼU�@Xj�H4@��I��!?=�M%7��@Qo�j�ٿfm��u�@L�0b9�3@S_�N�!?[$�bՕ@S�L��ٿ�}37��@�
^X�3@��")�!?���ɠ��@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@�G�ɛٿ!��]Z��@��4@d�D�!?T�^�@H�j�ٿ}������@�m���3@	.��b�!?���S�@H�j�ٿ}������@�m���3@	.��b�!?���S�@H�j�ٿ}������@�m���3@	.��b�!?���S�@�^e�,�ٿ5�.Q��@qP%�4@u�>Ð!?�m�`���@�^e�,�ٿ5�.Q��@qP%�4@u�>Ð!?�m�`���@�^e�,�ٿ5�.Q��@qP%�4@u�>Ð!?�m�`���@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@�DU`��ٿ�e3�W��@��� $4@DK�﹐!?:��L��@���i��ٿ��� R�@�d��k4@P"H���!?�7ՉX4�@���i��ٿ��� R�@�d��k4@P"H���!?�7ՉX4�@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@�9�6�ٿG�3�T�@�`�M�4@�]��!?a�ao�͕@Z1<+�ٿ�gې���@ewP>4@�_�ŏ!?�S�M�@Z1<+�ٿ�gې���@ewP>4@�_�ŏ!?�S�M�@Z1<+�ٿ�gې���@ewP>4@�_�ŏ!?�S�M�@! ��ٿbH�~�@�s�'�3@�$	2�!?��ж?�@! ��ٿbH�~�@�s�'�3@�$	2�!?��ж?�@�8s�h�ٿ66b[��@t� 4@�4����!?����m.�@w��ٿ`��lo��@���S�I4@$Q@�!?)�����@5�O�ٿ��$Z�@Q�KK`4@���v�!?�?��*��@5�O�ٿ��$Z�@Q�KK`4@���v�!?�?��*��@5�O�ٿ��$Z�@Q�KK`4@���v�!?�?��*��@5�O�ٿ��$Z�@Q�KK`4@���v�!?�?��*��@5�O�ٿ��$Z�@Q�KK`4@���v�!?�?��*��@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@����ٿ�`�xo��@�܀��o4@���b�!?s�>�@u0Gf��ٿ��9t>�@�5'�M4@oZ�2��!?l�"��@u0Gf��ٿ��9t>�@�5'�M4@oZ�2��!?l�"��@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@s�:N��ٿ�=��X��@�GL�I4@i7XvN�!?�K�k;�@��i��ٿ��iqߔ�@�G���,4@��27�!?��]-b�@��i��ٿ��iqߔ�@�G���,4@��27�!?��]-b�@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@֙��l�ٿ�R�H�f�@!��[!4@v�Z�!?��D ʕ@o��eΙٿ��`����@�П��84@���m|�!?M�'I�@o��eΙٿ��`����@�П��84@���m|�!?M�'I�@ �?Ҿ�ٿ��"���@x��K4@��|s;�!?CC-{��@ �?Ҿ�ٿ��"���@x��K4@��|s;�!?CC-{��@ �?Ҿ�ٿ��"���@x��K4@��|s;�!?CC-{��@}gzX�ٿ0�E`-Q�@�����"4@��&�'�!?A�Q_-��@}gzX�ٿ0�E`-Q�@�����"4@��&�'�!?A�Q_-��@}gzX�ٿ0�E`-Q�@�����"4@��&�'�!?A�Q_-��@j���ٿ�֯���@*�}04@��yA�!?�٦ك��@,�&
8�ٿ2g���@j���4@s%E3�!?tXzP�@,�&
8�ٿ2g���@j���4@s%E3�!?tXzP�@,�&
8�ٿ2g���@j���4@s%E3�!?tXzP�@xsA�F�ٿy9���@,�$V�34@���M�!?~~�l���@xsA�F�ٿy9���@,�$V�34@���M�!?~~�l���@xsA�F�ٿy9���@,�$V�34@���M�!?~~�l���@xsA�F�ٿy9���@,�$V�34@���M�!?~~�l���@�3�`�ٿ���݀�@`�:���3@�w�?G�!?��0���@�3�`�ٿ���݀�@`�:���3@�w�?G�!?��0���@�3�`�ٿ���݀�@`�:���3@�w�?G�!?��0���@mO��Y�ٿc1�Ϋ��@�G���4@p�gF�!?�5p��@mO��Y�ٿc1�Ϋ��@�G���4@p�gF�!?�5p��@mO��Y�ٿc1�Ϋ��@�G���4@p�gF�!?�5p��@mO��Y�ٿc1�Ϋ��@�G���4@p�gF�!?�5p��@mO��Y�ٿc1�Ϋ��@�G���4@p�gF�!?�5p��@����&�ٿ�hGrB��@�gx��3@����B�!?|���@����&�ٿ�hGrB��@�gx��3@����B�!?|���@��	�ҝٿ*�_i�+�@����4@���!?t���ݕ@��	�ҝٿ*�_i�+�@����4@���!?t���ݕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@T=@U�ٿ`}E�@�Cq)t�3@ݝi�7�!?.��0ҕ@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@]*��K�ٿ��z��@�(�~4@�&s���!?/1]���@*�(!�ٿ�d�۔��@I}zb��3@��ɩ��!?�F!�@*�(!�ٿ�d�۔��@I}zb��3@��ɩ��!?�F!�@괙��ٿ۶S۬��@f����3@
#�M�!?�Z�r6V�@괙��ٿ۶S۬��@f����3@
#�M�!?�Z�r6V�@괙��ٿ۶S۬��@f����3@
#�M�!?�Z�r6V�@괙��ٿ۶S۬��@f����3@
#�M�!?�Z�r6V�@�u�5"�ٿ�T�^��@0i4@��]	N�!?^�6i5�@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@n���Y�ٿ"�^:_k�@o2u���3@V���!?�σ5��@F	�B��ٿ[��eK#�@���{�3@�2X�!?x��?��@F	�B��ٿ[��eK#�@���{�3@�2X�!?x��?��@F	�B��ٿ[��eK#�@���{�3@�2X�!?x��?��@l�
��ٿ[?�ң��@��� 24@�1
Χ�!?��Q
	@l�
��ٿ[?�ң��@��� 24@�1
Χ�!?��Q
	@l�
��ٿ[?�ң��@��� 24@�1
Χ�!?��Q
	@l�
��ٿ[?�ң��@��� 24@�1
Χ�!?��Q
	@�ܒI�ٿbZQ.
�@�)�j%�3@s]��J�!?��	�p�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@��ry�ٿ�e���@r��ݜ4@�/{P�!?��l
/�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@�G<ʚٿ�C����@"���3@Jzo�>�!?�r�M&�@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@��;���ٿ1.xNJ=�@�ҿu+�3@�E^L�!?�1#�j��@�du�ٿ(ג�@Jo��)4@����!?��쨕��@0Y��.�ٿW�ޠ���@�����4@�Ē�(�!?���g�Ε@0Y��.�ٿW�ޠ���@�����4@�Ē�(�!?���g�Ε@�U#H��ٿ���d���@I(O��3@�E�4�!?jLh��Ε@���Q�ٿ)��A�@����4@�wq,%�!?�O26�<�@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�c0Ɍ�ٿ�3g�T�@A� �;�3@�oU�!?��݌D��@�⬠ٿ�+$��@P���3@���2�!?���t�@�|�ٿ�0����@_[0��3@D^���!?}&zZH�@Y�[�Y�ٿe�%�)�@S�>r�4@�Lޘ�!?��\�)�@Y�[�Y�ٿe�%�)�@S�>r�4@�Lޘ�!?��\�)�@Y�[�Y�ٿe�%�)�@S�>r�4@�Lޘ�!?��\�)�@Y�[�Y�ٿe�%�)�@S�>r�4@�Lޘ�!?��\�)�@AU� Q�ٿ¹�\"�@m�J�(R4@�D:�!?����O7�@AU� Q�ٿ¹�\"�@m�J�(R4@�D:�!?����O7�@AU� Q�ٿ¹�\"�@m�J�(R4@�D:�!?����O7�@����ٿ��6��@ƌ�@4@6�ޢ�!?�a��W��@����ٿ��6��@ƌ�@4@6�ޢ�!?�a��W��@����ٿ��6��@ƌ�@4@6�ޢ�!?�a��W��@����ٿ��6��@ƌ�@4@6�ޢ�!?�a��W��@n�3~�ٿ?0�l�@�'��:4@���Ma�!?���+�@n�3~�ٿ?0�l�@�'��:4@���Ma�!?���+�@n�3~�ٿ?0�l�@�'��:4@���Ma�!?���+�@n�3~�ٿ?0�l�@�'��:4@���Ma�!?���+�@�A@�	�ٿ��G�@��tk�4@JpRj��!?+X�K�@kDc��ٿ笑z���@��c6�4@��<!?����n�@kDc��ٿ笑z���@��c6�4@��<!?����n�@r	b+�ٿj�dz�@��ظ�3@�:y��!?���ق�@p�ő��ٿ��5�v9�@�6�p�4@�PpD�!?�m�I�@!l�s�ٿb����h�@�9 >4@�����!?�Ӹ%�@!l�s�ٿb����h�@�9 >4@�����!?�Ӹ%�@!l�s�ٿb����h�@�9 >4@�����!?�Ӹ%�@��ߢٿ{A����@���64@W�AJ��!?�� P s�@�q���ٿ_þa���@o^�7��3@��%�8�!?���o|3�@�n���ٿ(�u7���@��`�3@�NHi��!?nA����@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@<A�ٿ$��b��@#�p{�4@.ɬ�a�!?��~��@��gۡٿyHE/�@��60
4@�;�'ΐ!?�=��@��Lf�ٿ�=��@A�E�3@��o\��!?�.���`�@��Lf�ٿ�=��@A�E�3@��o\��!?�.���`�@��Lf�ٿ�=��@A�E�3@��o\��!?�.���`�@uHi�%�ٿIk�'[��@��n_^�3@��"F�!?H�f��˕@uHi�%�ٿIk�'[��@��n_^�3@��"F�!?H�f��˕@Eⱏ��ٿ�ɲVڂ�@�t�aC�3@ �^��!?T����@Eⱏ��ٿ�ɲVڂ�@�t�aC�3@ �^��!?T����@Eⱏ��ٿ�ɲVڂ�@�t�aC�3@ �^��!?T����@&�o�ٿ~�<<��@F*���3@��i-T�!?i��^�;�@&�o�ٿ~�<<��@F*���3@��i-T�!?i��^�;�@&�o�ٿ~�<<��@F*���3@��i-T�!?i��^�;�@&�o�ٿ~�<<��@F*���3@��i-T�!?i��^�;�@&�o�ٿ~�<<��@F*���3@��i-T�!?i��^�;�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@8�G�ٿ����2��@}N�p44@�[��B�!?N��i�@3��Օٿ�0�w�w�@��	94@n��}d�!?4��sY�@3��Օٿ�0�w�w�@��	94@n��}d�!?4��sY�@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@B�×ٿF�B�I��@S���4@�;�w�!?f*n�ߕ@.�`W�ٿ{ȸ<��@�N����3@��w�!?@�	�\��@.�`W�ٿ{ȸ<��@�N����3@��w�!?@�	�\��@&"2I[�ٿ���s�@Ӛ2��3@$C��f�!?��1����@�܋�ٿckQ�e�@�t�2�3@�-[ m�!?Ǐ�Qȕ@�܋�ٿckQ�e�@�t�2�3@�-[ m�!?Ǐ�Qȕ@������ٿ��:�@�	�n�3@�?�?t�!?�0#���@������ٿ��:�@�	�n�3@�?�?t�!?�0#���@������ٿ��:�@�	�n�3@�?�?t�!?�0#���@��s�ٿ��Rf�@��ma�3@X���Z�!?�f�����@��s�ٿ��Rf�@��ma�3@X���Z�!?�f�����@��s�ٿ��Rf�@��ma�3@X���Z�!?�f�����@�uLV��ٿ[U��kd�@�1�p��3@0��)_�!?��9"���@�uLV��ٿ[U��kd�@�1�p��3@0��)_�!?��9"���@�uLV��ٿ[U��kd�@�1�p��3@0��)_�!?��9"���@�uLV��ٿ[U��kd�@�1�p��3@0��)_�!?��9"���@�uLV��ٿ[U��kd�@�1�p��3@0��)_�!?��9"���@S?��ЖٿN$2��Z�@��X�e'4@��dD�!?Yf#6I�@S?��ЖٿN$2��Z�@��X�e'4@��dD�!?Yf#6I�@S?��ЖٿN$2��Z�@��X�e'4@��dD�!?Yf#6I�@S?��ЖٿN$2��Z�@��X�e'4@��dD�!?Yf#6I�@S?��ЖٿN$2��Z�@��X�e'4@��dD�!?Yf#6I�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@��Y�ٿ�`����@����A4@�Z]��!?+��-ܒ�@UQ��%�ٿ�57�Z�@`��W4@��ʥ�!?�.P!;ܕ@UQ��%�ٿ�57�Z�@`��W4@��ʥ�!?�.P!;ܕ@UQ��%�ٿ�57�Z�@`��W4@��ʥ�!?�.P!;ܕ@%�#K��ٿ�e.�@"���d4@�/`1ѐ!?ĉɖ�@�V:�ٿN�*�K�@��~�-�3@O B��!?�9he�ߕ@�V:�ٿN�*�K�@��~�-�3@O B��!?�9he�ߕ@�V:�ٿN�*�K�@��~�-�3@O B��!?�9he�ߕ@^���ٿ8\N!��@�ſ��04@v.�(��!?x���]�@k��<��ٿm0Y9��@�����3@�艙ѐ!?�U(yȕ@.� "�ٿܕ���$�@�� �3@�g��!?Ĵϲ@��@.� "�ٿܕ���$�@�� �3@�g��!?Ĵϲ@��@.� "�ٿܕ���$�@�� �3@�g��!?Ĵϲ@��@.� "�ٿܕ���$�@�� �3@�g��!?Ĵϲ@��@��ia��ٿ�Tzз�@�1$��3@�<��O�!?�r�N��@��ia��ٿ�Tzз�@�1$��3@�<��O�!?�r�N��@��ia��ٿ�Tzз�@�1$��3@�<��O�!?�r�N��@ei�23�ٿ-A�4��@J��fh4@0ý�Q�!?�ҙ"��@ei�23�ٿ-A�4��@J��fh4@0ý�Q�!?�ҙ"��@ei�23�ٿ-A�4��@J��fh4@0ý�Q�!?�ҙ"��@ei�23�ٿ-A�4��@J��fh4@0ý�Q�!?�ҙ"��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@��O	�ٿ�ű���@_�~��64@��B�.�!?oJ�U��@�s�<��ٿ��[�?�@k[9Ut94@V���!�!?*�C?��@�s�<��ٿ��[�?�@k[9Ut94@V���!�!?*�C?��@5z����ٿ O��,�@�4`�r.4@�6E(�!?�p��蜕@5z����ٿ O��,�@�4`�r.4@�6E(�!?�p��蜕@Q�S��ٿ�k#���@Vjq[H4@����X�!?��(��̕@A��$`�ٿ�������@^Fd�W4@�Pm8��!?��Κ�i�@A��$`�ٿ�������@^Fd�W4@�Pm8��!?��Κ�i�@A��$`�ٿ�������@^Fd�W4@�Pm8��!?��Κ�i�@A��$`�ٿ�������@^Fd�W4@�Pm8��!?��Κ�i�@A��$`�ٿ�������@^Fd�W4@�Pm8��!?��Κ�i�@��f��ٿ���J#��@���J4@�=S�!?1��1�@��f��ٿ���J#��@���J4@�=S�!?1��1�@��f��ٿ���J#��@���J4@�=S�!?1��1�@��f��ٿ���J#��@���J4@�=S�!?1��1�@��f��ٿ���J#��@���J4@�=S�!?1��1�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@�T�ٿ����v�@�LsDgP4@�T�X�!?���Qg�@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��x��ٿ^����@��L�84@�%��!?W��~HÕ@��`N�ٿF�5�h��@8��g�*4@Sr�0Ґ!?��1�h��@��`N�ٿF�5�h��@8��g�*4@Sr�0Ґ!?��1�h��@Ĳ�Ga�ٿ$�/W��@���qo
4@�Kb�ʐ!?IX^��֕@Ĳ�Ga�ٿ$�/W��@���qo
4@�Kb�ʐ!?IX^��֕@A�l �ٿ�rf���@n*��D4@�Jd�p�!?� ���@A�l �ٿ�rf���@n*��D4@�Jd�p�!?� ���@�F�G	�ٿ����M��@7�v�3@)��WP�!?����Ε@�F�G	�ٿ����M��@7�v�3@)��WP�!?����Ε@�F�G	�ٿ����M��@7�v�3@)��WP�!?����Ε@�F�G	�ٿ����M��@7�v�3@)��WP�!?����Ε@�?j幥ٿt35��@)�p�3@���*�!?܉��zÕ@�?j幥ٿt35��@)�p�3@���*�!?܉��zÕ@�?j幥ٿt35��@)�p�3@���*�!?܉��zÕ@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@�ª��ٿ"a�K��@ˏ���3@쏁4�!?��n����@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@ �dG�ٿ����A�@H���J�3@���!?��y�@�ɠٿuٞI�@��'�3@vh�9��!?����@�ɠٿuٞI�@��'�3@vh�9��!?����@�ɠٿuٞI�@��'�3@vh�9��!?����@�ɠٿuٞI�@��'�3@vh�9��!?����@�ɠٿuٞI�@��'�3@vh�9��!?����@�ɠٿuٞI�@��'�3@vh�9��!?����@l����ٿ �y���@��mi�3@PgmK^�!?���>�@l����ٿ �y���@��mi�3@PgmK^�!?���>�@l����ٿ �y���@��mi�3@PgmK^�!?���>�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@j��|}�ٿt#)�S�@�� �*�3@p;�}�!?�m" X�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@T:�U^�ٿp�_�#��@=͏�z4@b �H��!?(O�nq�@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@d0��c�ٿoŒ*���@N4��I4@�N|0�!?�j���@�Y�ٿ�뮡�@QT��f4@bm�%�!?�wM�ĕ�@z.�P�ٿx!�H�@h�(g<4@ɬ��+�!?� S'��@z.�P�ٿx!�H�@h�(g<4@ɬ��+�!?� S'��@z.�P�ٿx!�H�@h�(g<4@ɬ��+�!?� S'��@z.�P�ٿx!�H�@h�(g<4@ɬ��+�!?� S'��@������ٿuA��@��?4@�`thC�!?լ��@������ٿuA��@��?4@�`thC�!?լ��@������ٿuA��@��?4@�`thC�!?լ��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�mR�ٿ�d����@fT��!4@[I�&�!?��@��@�&�.�ٿm����@Rm�*�-4@ø�g�!?�3l	�@,�[�ٿ��nL܊�@O'�Z%4@5j����!?0���ȕ@.�;[{�ٿd��LI�@�*���,4@F�7��!?�I?�r��@�a��ٿj���>�@_��mN�3@��L�$�!?����{�@�a��ٿj���>�@_��mN�3@��L�$�!?����{�@�a��ٿj���>�@_��mN�3@��L�$�!?����{�@���?�ٿ�<y�@�1/:4@,���#�!?�o}4X��@���?�ٿ�<y�@�1/:4@,���#�!?�o}4X��@���?�ٿ�<y�@�1/:4@,���#�!?�o}4X��@�9�T�ٿG�iX���@i��KQ4@ ��eQ�!?
�-�?��@v|���ٿ.ϱg���@�bI��4@'E���!?� Q�/��@μ��ٿ�$��F�@ک��+4@�L�i(�!?���"x�@�\�+a�ٿ�\�M7�@�ݪ,1*4@�7��!?�Tu/J��@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@ ċ[��ٿ�p_u�<�@�i5�4@<׸%�!?��?�6�@i�ܤٿ5�x���@�1���4@���4�!?'�N�{��@i�ܤٿ5�x���@�1���4@���4�!?'�N�{��@�{�Ow�ٿ�
�]��@�f�A4@��P �!?"~�(R��@�\��ٿ>��Q��@8�HV��3@�a�!?��;/�@�\��ٿ>��Q��@8�HV��3@�a�!?��;/�@�\��ٿ>��Q��@8�HV��3@�a�!?��;/�@�\��ٿ>��Q��@8�HV��3@�a�!?��;/�@s~X,�ٿ$��v���@����4@�Ud���!?Ƌ�s��@tMA ��ٿTf8O��@���4@C�'��!?#���@tMA ��ٿTf8O��@���4@C�'��!?#���@tMA ��ٿTf8O��@���4@C�'��!?#���@tMA ��ٿTf8O��@���4@C�'��!?#���@tMA ��ٿTf8O��@���4@C�'��!?#���@�k)əٿ�]�GP��@&��-�4@<�"7�!?\d�l<l�@/�%^J�ٿ���(��@��ӈ[4@
�i%��!?P��8�@/�%^J�ٿ���(��@��ӈ[4@
�i%��!?P��8�@/�%^J�ٿ���(��@��ӈ[4@
�i%��!?P��8�@�z��,�ٿ�qS���@,�k�t&4@G����!?v.�$�@�z��,�ٿ�qS���@,�k�t&4@G����!?v.�$�@�L0Y�ٿ����k�@Gp��d�3@�#(6P�!?7;��"�@p��|�ٿӯIhǧ�@�[*�y�3@F�7��!?Ш��R3�@p��|�ٿӯIhǧ�@�[*�y�3@F�7��!?Ш��R3�@p��|�ٿӯIhǧ�@�[*�y�3@F�7��!?Ш��R3�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@���k�ٿ��J��h�@e�"�7�3@�s��!?�W�G�@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@�M�/��ٿu9Ws\�@��~M4@�2��"�!?	��ع��@���E�ٿ��)L�K�@���+	4@�G�<B�!?8�G��@���E�ٿ��)L�K�@���+	4@�G�<B�!?8�G��@���E�ٿ��)L�K�@���+	4@�G�<B�!?8�G��@���E�ٿ��)L�K�@���+	4@�G�<B�!?8�G��@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@�Hp���ٿ�IPtJ�@T���C4@r��Ll�!?%�z�� �@hٱ±�ٿ/&[�B�@�;kP�4@��|���!?��"���@ζ���ٿH��=�B�@�ܵ�g?4@�Z�kd�!?� %I͕@���Z�ٿ��!&�b�@C�gTI4@*��23�!?��5Ǜ'�@���Z�ٿ��!&�b�@C�gTI4@*��23�!?��5Ǜ'�@���Z�ٿ��!&�b�@C�gTI4@*��23�!?��5Ǜ'�@���Z�ٿ��!&�b�@C�gTI4@*��23�!?��5Ǜ'�@���Z�ٿ��!&�b�@C�gTI4@*��23�!?��5Ǜ'�@