�NUMPY v {'descr': '<f8', 'fortran_order': False, 'shape': (3, 10000, 5), }                                                   
������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@�?W:��ٿA��l ��@���I��3@Z�Q�_�!? ���o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@������ٿǞ9] ��@ڸ��  4@� qŏ!?�����o�@y֭#{�ٿOc�T ��@�N�| 4@Kg}��!?q�r��o�@y֭#{�ٿOc�T ��@�N�| 4@Kg}��!?q�r��o�@y֭#{�ٿOc�T ��@�N�| 4@Kg}��!?q�r��o�@:5��y�ٿ�keg ��@iU�g 4@�T๏!?{����o�@:5��y�ٿ�keg ��@iU�g 4@�T๏!?{����o�@:5��y�ٿ�keg ��@iU�g 4@�T๏!?{����o�@:5��y�ٿ�keg ��@iU�g 4@�T๏!?{����o�@:5��y�ٿ�keg ��@iU�g 4@�T๏!?{����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@`/��u�ٿT��c ��@w� 4@�����!?�����o�@@���|�ٿ�w�L ��@Z�  4@�*��a�!?~>���o�@@���|�ٿ�w�L ��@Z�  4@�*��a�!?~>���o�@@���|�ٿ�w�L ��@Z�  4@�*��a�!?~>���o�@7:|hl�ٿ���Q ��@��Og 4@_��#��!?����o�@7:|hl�ٿ���Q ��@��Og 4@_��#��!?����o�@7:|hl�ٿ���Q ��@��Og 4@_��#��!?����o�@�9Ӗn�ٿ�=�X ��@�<{� 4@�$ƨ��!?~���o�@�9Ӗn�ٿ�=�X ��@�<{� 4@�$ƨ��!?~���o�@�9Ӗn�ٿ�=�X ��@�<{� 4@�$ƨ��!?~���o�@�9Ӗn�ٿ�=�X ��@�<{� 4@�$ƨ��!?~���o�@pSтx�ٿ���Y ��@& �l 4@�z ڏ!?^$��o�@pSтx�ٿ���Y ��@& �l 4@�z ڏ!?^$��o�@pSтx�ٿ���Y ��@& �l 4@�z ڏ!?^$��o�@�?	%~�ٿ]�9H ��@2al� 4@��X�ɏ!?>���o�@�?	%~�ٿ]�9H ��@2al� 4@��X�ɏ!?>���o�@�?	%~�ٿ]�9H ��@2al� 4@��X�ɏ!?>���o�@�?	%~�ٿ]�9H ��@2al� 4@��X�ɏ!?>���o�@�?	%~�ٿ]�9H ��@2al� 4@��X�ɏ!?>���o�@QU�z�ٿ���F ��@J��� 4@����!?dp��o�@QU�z�ٿ���F ��@J��� 4@����!?dp��o�@QU�z�ٿ���F ��@J��� 4@����!?dp��o�@g�T�~�ٿ�.�I ��@�/ 4@y�6S��!?|�
��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�C����ٿ��Q ��@�$� 4@^�i��!?r��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�}�Ձ�ٿ:�P ��@+x�� 4@ߐ� �!?�5~��o�@�VZՀ�ٿ1oQ ��@��H 4@�h�*ُ!?'#��o�@�VZՀ�ٿ1oQ ��@��H 4@�h�*ُ!?'#��o�@�����ٿዉM ��@X/  4@*4?���!?�����o�@�����ٿዉM ��@X/  4@*4?���!?�����o�@�[��}�ٿ��DO ��@j�qA 4@d+iK�!?���o�@�[��}�ٿ��DO ��@j�qA 4@d+iK�!?���o�@����~�ٿ9'�O ��@�M�o 4@��o��!?3�M��o�@����~�ٿ9'�O ��@�M�o 4@��o��!?3�M��o�@Ո(�|�ٿzdR ��@��� 4@�xr�s�!?X�a��o�@�\[�ٿ��P ��@D�� 4@	U�m̏!?���o�@�\[�ٿ��P ��@D�� 4@	U�m̏!?���o�@G��}�ٿ*6?W ��@Hh�� 4@>���!?x4���o�@�s�^��ٿW�YT ��@�\2 4@]~ mȏ!?G���o�@sE=�}�ٿ���P ��@
�gR 4@ī亏!?�@��o�@��J~�ٿ]��V ��@��2 4@��;��!?2�d��o�@��J~�ٿ]��V ��@��2 4@��;��!?2�d��o�@��J~�ٿ]��V ��@��2 4@��;��!?2�d��o�@��J~�ٿ]��V ��@��2 4@��;��!?2�d��o�@s�&��ٿ��rT ��@ ;r�  4@t ����!?�ɑ��o�@J��|�ٿ��U ��@�(�  4@�@�mď!?�N0��o�@���x�ٿU��Q ��@��'�  4@؎���!?�����o�@���x�ٿU��Q ��@��'�  4@؎���!?�����o�@��,�|�ٿ�*�R ��@R&M� 4@���>��!?��/��o�@�EZ�y�ٿEu�Q ��@q	�z 4@��5₏!?
����o�@�EZ�y�ٿEu�Q ��@q	�z 4@��5₏!?
����o�@&4��}�ٿ^��M ��@�b�� 4@�=ԅ�!?k���o�@&4��}�ٿ^��M ��@�b�� 4@�=ԅ�!?k���o�@BE�/�ٿ�7K ��@�0g8 4@�>^r��!?�e��o�@]e���ٿ��J ��@�V 4@�[gq��!?ǽ��o�@]e���ٿ��J ��@�V 4@�[gq��!?ǽ��o�@!8jU��ٿ�:H ��@@�� 4@����!?�1��o�@!8jU��ٿ�:H ��@@�� 4@����!?�1��o�@!8jU��ٿ�:H ��@@�� 4@����!?�1��o�@�z�悙ٿ�NH ��@%O/� 4@++S۰�!?
�#��o�@�U��ٿ �E ��@�l�� 4@u�lCˏ!?�`��o�@�U��ٿ �E ��@�l�� 4@u�lCˏ!?�`��o�@v^o<��ٿ��NG ��@�=aQ 4@��ߏ!?MU��o�@v^o<��ٿ��NG ��@�=aQ 4@��ߏ!?MU��o�@v^o<��ٿ��NG ��@�=aQ 4@��ߏ!?MU��o�@�`ק��ٿ�NtG ��@�YS> 4@e�xɳ�!?��O��o�@�`ק��ٿ�NtG ��@�YS> 4@e�xɳ�!?��O��o�@	�#��ٿ�$8J ��@l� 4@�OI6��!?�G��o�@B錇�ٿ� I ��@��y; 4@�La�y�!?\wq��o�@��	3��ٿN��H ��@�R� 4@��t'm�!?�ە��o�@��	3��ٿN��H ��@�R� 4@��t'm�!?�ە��o�@��	3��ٿN��H ��@�R� 4@��t'm�!?�ە��o�@������ٿ�sK ��@�)�� 4@�S�6�!?����o�@������ٿ�sK ��@�)�� 4@�S�6�!?����o�@������ٿ�sK ��@�)�� 4@�S�6�!?����o�@�О��ٿ%[O ��@j�a� 4@�ۼ@E�!?�]���o�@�v|�}�ٿZ�K ��@`�� 4@qz�UP�!?���o�@�ث|�ٿz�M ��@��{� 4@([u��!?�z��o�@�0��|�ٿ%��Q ��@��2� 4@�5�e��!?�-��o�@�0��|�ٿ%��Q ��@��2� 4@�5�e��!?�-��o�@�0��|�ٿ%��Q ��@��2� 4@�5�e��!?�-��o�@�0��|�ٿ%��Q ��@��2� 4@�5�e��!?�-��o�@�x��z�ٿŲ�R ��@?�5 4@ڃ����!?�R���o�@�x��z�ٿŲ�R ��@?�5 4@ڃ����!?�R���o�@V�Y{�ٿm�YP ��@Dx� 4@���ц�!?�;���o�@S�l�t�ٿ�%�P ��@�E� 4@Tl�-��!?K���o�@S�l�t�ٿ�%�P ��@�E� 4@Tl�-��!?K���o�@��jet�ٿ���S ��@le� 4@��"��!?B����o�@�Cv�ٿ�җT ��@��?� 4@����!?:���o�@��_x�ٿU$X ��@"��� 4@n�͂X�!?��5��o�@���w�ٿ�JZV ��@�m� 4@8�9�!?oc$��o�@��!�w�ٿ��U ��@�DJ� 4@���Z�!?0�y��o�@��!�w�ٿ��U ��@�DJ� 4@���Z�!?0�y��o�@/J}v�ٿ�\W ��@hأ 4@o)T_P�!?jo���o�@/J}v�ٿ�\W ��@hأ 4@o)T_P�!?jo���o�@��e]z�ٿE��U ��@a�% 4@�ut�!?oИ��o�@�E<�{�ٿw�#[ ��@9�� 4@��o�!? �.��o�@ʙ<-{�ٿ���X ��@L�]� 4@���|��!?8�p��o�@f�s|�ٿ���X ��@8� 4@���Y��!?i�ۻ�o�@�A�|�ٿ���V ��@L�.� 4@��䨏!?*\Q��o�@�S����ٿs��U ��@D��` 4@l�9�!?
�8��o�@����~�ٿ�)�V ��@���� 4@�\����!?���o�@����~�ٿ�)�V ��@���� 4@�\����!?���o�@�?�y��ٿ9�R ��@cTP� 4@���1�!?YK��o�@2��S��ٿ�|�S ��@ߐ� 4@ÉG��!?��l��o�@2��S��ٿ�|�S ��@ߐ� 4@ÉG��!?��l��o�@2��S��ٿ�|�S ��@ߐ� 4@ÉG��!?��l��o�@�����ٿ�T~S ��@�ޯ 4@	�D�؏!?b"��o�@if�ہ�ٿ�K�U ��@�P� 4@����!?uq��o�@��l��ٿy}�X ��@i2` 4@�#'u�!?����o�@��l��ٿy}�X ��@i2` 4@�#'u�!?����o�@��l��ٿy}�X ��@i2` 4@�#'u�!?����o�@�B���ٿQIX ��@�E�� 4@�tdЏ!?Sˋ��o�@4�[���ٿ�k�X ��@�� 4@�Z���!?���o�@G�ˆ�ٿo�Y ��@0� 4@rQ�^��!?ƭ���o�@�N�"��ٿ���W ��@�U$� 4@����!?�<1��o�@�N�"��ٿ���W ��@�U$� 4@����!?�<1��o�@Ù&��ٿz{�W ��@~Z�� 4@�^�.
�!?(���o�@=�̊�ٿ:�6Y ��@DqT� 4@��(aƏ!?꿋��o�@=�̊�ٿ:�6Y ��@DqT� 4@��(aƏ!?꿋��o�@Q�M��ٿIy[ ��@�&T� 4@�̀ߏ!?9����o�@ы3���ٿ���^ ��@��� 4@�P!�Ϗ!?�$��o�@��Q���ٿ,��[ ��@9J� 4@��!?y���o�@z�=.��ٿ��B] ��@,��� 4@��k�"�!?�$p��o�@߱�R��ٿ���[ ��@�/A� 4@?�A:�!?�9~��o�@߱�R��ٿ���[ ��@�/A� 4@?�A:�!?�9~��o�@߱�R��ٿ���[ ��@�/A� 4@?�A:�!?�9~��o�@߱�R��ٿ���[ ��@�/A� 4@?�A:�!?�9~��o�@F��ٿh�>Y ��@
��� 4@cN�-��!?��o�@@�b�ٿG�yX ��@���� 4@Ӛ�=��!?o�,��o�@@�b�ٿG�yX ��@���� 4@Ӛ�=��!?o�,��o�@{j�m��ٿ96\ ��@��� 4@]QS��!?61&��o�@C�I��ٿ�K�W ��@�+�� 4@��l̏!?U�;��o�@�n���ٿ71�S ��@�Yǣ 4@�"z�!?,���o�@�����ٿ��*V ��@~&�n 4@\&��x�!?$��o�@�TMl��ٿz��Y ��@F0_ 4@������!?F���o�@�-Q���ٿ��X ��@�,�U 4@F����!?��v��o�@t����ٿ��7T ��@ET�S 4@�6$���!?�K���o�@t����ٿ��7T ��@ET�S 4@�6$���!?�K���o�@���Z��ٿ��R ��@�ua 4@)�d��!?����o�@~=�:��ٿ4�Z ��@�^ 4@C.\7�!?6����o�@~=�:��ٿ4�Z ��@�^ 4@C.\7�!?6����o�@~=�:��ٿ4�Z ��@�^ 4@C.\7�!?6����o�@c:⚆�ٿ�>�[ ��@T	�D 4@����!?���o�@#&����ٿg�q] ��@L��a 4@�͚��!?eFں�o�@��E���ٿ�\ ��@�	?z 4@=5G�!?�
���o�@��E���ٿ�\ ��@�	?z 4@=5G�!?�
���o�@siiH��ٿD\�Z ��@?�_ 4@C�z�!?����o�@������ٿ��/Y ��@��, 4@j�F�!?n����o�@�ڀ�ٿ��[ ��@�0d3 4@��qS�!?ɭ{��o�@��.b��ٿY ��@s�' 4@����!?7��o�@�gy��ٿ	��[ ��@�}B 4@;�n�̏!?�Pu��o�@��/��ٿ8�[ ��@��: 4@)����!?�<���o�@�uj~�ٿ�\[ ��@�re� 4@!~(ɏ!?yΜ��o�@Q�dw}�ٿ
��X ��@N� 4@|[�T�!?�!��o�@5�'|�ٿ���Z ��@/� � 4@1�٩��!?����o�@6�+}�ٿZ��V ��@�R� 4@�6;��!?�C&��o�@6�+}�ٿZ��V ��@�R� 4@�6;��!?�C&��o�@dê�~�ٿI�W ��@��� 4@#���!?�	׶�o�@�=E�{�ٿ�V ��@��V� 4@L�d�^�!?45���o�@�؋�}�ٿ;�T ��@J��� 4@��:�S�!? �´�o�@��n�~�ٿU�ZV ��@�ˍ� 4@(�˯Y�!?I{~��o�@ɑ�	��ٿ��cV ��@F0� 4@���i�!?��@��o�@dZ6|��ٿ��Y ��@2�-r 4@���g�!?ݶf��o�@|�~ٿm�<W ��@O�c 4@��>~��!?o�ù�o�@|�~ٿm�<W ��@O�c 4@��>~��!?o�ù�o�@|�~ٿm�<W ��@O�c 4@��>~��!?o�ù�o�@��q��ٿ��Y ��@���+ 4@�:Zt�!?�п��o�@b�$^��ٿ�s.V ��@��� 4@�hi��!?�v���o�@�����ٿ�C�V ��@�G� 4@/V򧍏!?3�C��o�@�����ٿ�C�V ��@�G� 4@/V򧍏!?3�C��o�@�����ٿ�C�V ��@�G� 4@/V򧍏!?3�C��o�@+�'��ٿ�f9W ��@�� 4@�hJ�ԏ!?�����o�@0����ٿ�0�S ��@��kD 4@���s�!?$�@��o�@�� ���ٿ$y<X ��@�� 4@2?��!?^{��o�@�� ���ٿ$y<X ��@�� 4@2?��!?^{��o�@�^����ٿi�MV ��@����  4@�YHϏ!?����o�@C�f�ٿ��U ��@5A 4@�u2�֏!?�����o�@��^H��ٿ�4�W ��@a�c� 4@���&��!?��^��o�@5F����ٿ{�3\ ��@��� 4@���?�!?�����o�@<ǫ���ٿ`�O[ ��@���c 4@�N�P�!?��W��o�@�yȦ�ٿ�8�\ ��@���  4@�)��!?aJi��o�@�~aO��ٿ�A�Y ��@2_y�  4@ò-#�!?]�!��o�@�~aO��ٿ�A�Y ��@2_y�  4@ò-#�!?]�!��o�@f�:.��ٿ��W ��@	w�: 4@M� �؏!?�����o�@I�c֚�ٿ��,T ��@1�d 4@&�(��!?�J��o�@I�c֚�ٿ��,T ��@1�d 4@&�(��!?�J��o�@�~��ٿ�ɢS ��@W�* 4@��Dߦ�!?}���o�@�ͻ;��ٿ�JY ��@H [���3@B��i��!?�Ħ��o�@�ͻ;��ٿ�JY ��@H [���3@B��i��!?�Ħ��o�@�����ٿ�|W ��@�|���3@=�v!?�s��o�@�'~��ٿ��fZ ��@��Q���3@	�vfڏ!?�����o�@X�k��ٿ'U�Y ��@�t�M��3@k�B��!?B����o�@X�k��ٿ'U�Y ��@�t�M��3@k�B��!?B����o�@f�ɸ��ٿg�Y ��@�|����3@M~j�!?�XB��o�@�q#��ٿ�U�X ��@~$�-��3@��!?n�G��o�@�q#��ٿ�U�X ��@~$�-��3@��!?n�G��o�@\�,��ٿ^F�T ��@��+��3@��mGԏ!?����o�@o�𚡙ٿO�>U ��@���  4@�{��!?M�@��o�@�R���ٿ���T ��@�x� 4@���{�!?dQ ��o�@L���ٿ�X ��@ dj� 4@�Z����!?>���o�@_�et�ٿ��mY ��@��3 4@}��)U�!?\y���o�@_�et�ٿ��mY ��@��3 4@}��)U�!?\y���o�@ՙ���ٿDmtZ ��@��X  4@~%�Ə!?����o�@ՙ���ٿDmtZ ��@��X  4@~%�Ə!?����o�@�s=��ٿ��[ ��@c1���3@�O�<�!?���o�@����ٿ�uY ��@4�;���3@o�I7�!?&+��o�@����ٿ�uY ��@4�;���3@o�I7�!?&+��o�@%���̙ٿ�bW ��@��P���3@�zZ֏!?����o�@�.�ϙٿ&8�T ��@�䠚��3@��jɏ!?@A���o�@�.�ϙٿ&8�T ��@�䠚��3@��jɏ!?@A���o�@.LIz��ٿK7]S ��@M�:"��3@����!?����o�@�)as��ٿ!�mT ��@ew!  4@�KD��!?_4��o�@D*"��ٿ�Q2R ��@��� 4@ލ[/��!?��6��o�@Z�����ٿӤP ��@T�z�  4@�v���!?�f*��o�@�?�~��ٿ)�R ��@�ue��3@�vᓏ!?�� ��o�@�?�~��ٿ)�R ��@�ue��3@�vᓏ!?�� ��o�@W�ȁ��ٿxZ�O ��@�ġ���3@]��g�!?�R���o�@�&,X��ٿq�MP ��@�D�� 4@�mt�%�!?��o�@�&,X��ٿq�MP ��@�D�� 4@�mt�%�!?��o�@���t�ٿ���P ��@�Ps 4@�}9Q�!?���o�@���t�ٿ���P ��@�Ps 4@�}9Q�!?���o�@�4KZ`�ٿ5
�O ��@��om 4@;�a�5�!?'�D��o�@d�x�ٿ�fbN ��@��� 4@��w�:�!?�
x��o�@d�x�ٿ�fbN ��@��� 4@��w�:�!?�
x��o�@d�x�ٿ�fbN ��@��� 4@��w�:�!?�
x��o�@��C2��ٿS��O ��@&�M���3@��^�K�!?ȟ��o�@:��.��ٿ���M ��@/ˍW��3@5$��F�!?��U��o�@93��ٿAZ�P ��@�Ӳ��3@&�鐏!?�����o�@���֙ٿ*�Q ��@������3@,�?l�!?p����o�@���֙ٿ*�Q ��@������3@,�?l�!?p����o�@�����ٿ�N ��@k�����3@�4�x�!?�����o�@��υ��ٿ�K5O ��@ə����3@�Ӟ�!?����o�@��υ��ٿ�K5O ��@ə����3@�Ӟ�!?����o�@��υ��ٿ�K5O ��@ə����3@�Ӟ�!?����o�@��υ��ٿ�K5O ��@ə����3@�Ӟ�!?����o�@�g���ٿF�S ��@!{Sb��3@��M���!?����o�@�З��ٿ@�fS ��@�����3@W�U��!?s ���o�@���_�ٿc"X ��@�����3@��7�K�!?rwU��o�@���_�ٿc"X ��@�����3@��7�K�!?rwU��o�@���_�ٿc"X ��@�����3@��7�K�!?rwU��o�@=����ٿ��8^ ��@�9�  4@����\�!?� ���o�@1RC�ٿ�[ ��@[.�D 4@f�/�֏!?0?���o�@1RC�ٿ�[ ��@[.�D 4@f�/�֏!?0?���o�@%#��ٿG��Y ��@�uƏ  4@����̏!?�4��o�@%#��ٿG��Y ��@�uƏ  4@����̏!?�4��o�@\I����ٿ`g\ ��@���D 4@w�򫪏!?P�i��o�@��8��ٿMs�^ ��@�]g���3@'	!!��!?�����o�@�hĄ��ٿ�^\ ��@��;��3@�\�!?�d��o�@<�'Z��ٿءh^ ��@��� 4@7u�!?�/��o�@<�'Z��ٿءh^ ��@��� 4@7u�!?�/��o�@<�'Z��ٿءh^ ��@��� 4@7u�!?�/��o�@xF�#ƙٿ*�O ��@��:���3@��c��!?�j��o�@��ٜ�ٿ�u�N ��@�hu���3@ư���!?�P��o�@��c�f�ٿԣJS ��@� 4@�V{��!?3X��o�@��c�f�ٿԣJS ��@� 4@�V{��!?3X��o�@��c�f�ٿԣJS ��@� 4@�V{��!?3X��o�@��c�f�ٿԣJS ��@� 4@�V{��!?3X��o�@��c�f�ٿԣJS ��@� 4@�V{��!?3X��o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@lr�m�ٿ��Q ��@�f�� 4@uZ؜�!?㮳�o�@�S��'�ٿ;~�J ��@	��{ 4@�6e)O�!?3$��o�@?IϦb�ٿ�>�P ��@n`�F 4@V��c�!?�tY��o�@�X�H��ٿy��Y ��@��\  4@M�-��!?:�V��o�@���g��ٿl�Y ��@���0 4@���[�!?�o��o�@Zw�V~�ٿ4,P^ ��@l1�� 4@���x�!?%:��o�@G H��ٿaBc ��@G�\j 4@=���!?�����o�@���籙ٿ��
[ ��@�V0���3@��7ǋ�!?���o�@f"�C�ٿ��] ��@Ez4���3@X��ԏ!?�B0��o�@���P�ٿZ�k[ ��@��p���3@�/��u�!?����o�@�Q�3��ٿ�эV ��@�e����3@j��ں�!?�����o�@�Q�3��ٿ�эV ��@�e����3@j��ں�!?�����o�@��<��ٿq�Y^ ��@"s���3@y���ޏ!?� N��o�@N�Y��ٿ9�/[ ��@4����3@]J���!?m���o�@N�Y��ٿ9�/[ ��@4����3@]J���!?m���o�@�C���ٿӉ�\ ��@���,��3@��$��!?�����o�@�C���ٿӉ�\ ��@���,��3@��$��!?�����o�@���m�ٿN�[ ��@�/۝��3@�<;�!?Wx���o�@Y01�ٿ�T_ ��@���:��3@t�˭��!?2�w��o�@Wa�n,�ٿ8ZcU ��@7����3@ۿ�֏!?��|��o�@��3f<�ٿ0o�\ ��@ �����3@� ~Տ!?�,��o�@��3f<�ٿ0o�\ ��@ �����3@� ~Տ!?�,��o�@B��Ŭ�ٿd�d ��@1�b���3@u���ޏ!?�"��o�@6��t�ٿ&��` ��@Jc�`��3@u vƏ!?�M!��o�@6��t�ٿ&��` ��@Jc�`��3@u vƏ!?�M!��o�@�����ٿ��c ��@�h� ��3@��P�!?�C-��o�@�����ٿ��c ��@�h� ��3@��P�!?�C-��o�@�����ٿ��c ��@�h� ��3@��P�!?�C-��o�@0�k��ٿ%��m ��@�h"F��3@q#�
�!?Ĳ��o�@0�k��ٿ%��m ��@�h"F��3@q#�
�!?Ĳ��o�@�'Gj��ٿ 9�` ��@X����3@�����!?��@��o�@�'Gj��ٿ 9�` ��@X����3@�����!?��@��o�@۸�%�ٿ�$7i ��@�t!r��3@ �Ne~�!?/�:�o�@���ٿ�8j ��@�ھ���3@�7z��!?HC��o�@�����ٿV�v ��@ڐ�F��3@��ɏ!?jg}#�o�@FN٩�ٿ6Tl ��@�����3@��ҏ!?]�0��o�@FN٩�ٿ6Tl ��@�����3@��ҏ!?]�0��o�@K-Y�D�ٿn|�Y ��@��� 4@V�<L��!?�Y4��o�@K-Y�D�ٿn|�Y ��@��� 4@V�<L��!?�Y4��o�@�)Ѕ��ٿ%fh ��@���> 4@�,Is��!?�L���o�@(˂\ڙٿ�wL� ��@���j 4@F�-���!?�2���o�@}�8 �ٿ*w9| ��@���"��3@��o �!?#׵��o�@}�8 �ٿ*w9| ��@���"��3@��o �!?#׵��o�@����E�ٿ�xWo ��@U[s� 4@�D]�!?�~B��o�@�"Ȍ�ٿA�pR ��@��D; 4@s�꫏!?�]�y�o�@O��E�ٿ�.&b ��@�f\
	 4@�sz�
�!?��˙�o�@o��ٿ�o�x ��@���	 4@�&%�!?��;��o�@�	���ٿ���o ��@ ci	 4@�%��!?u����o�@��C �ٿ;.Z ��@� 4@��2o��!?��5��o�@��C �ٿ;.Z ��@� 4@��2o��!?��5��o�@K�5�ٿ���d ��@�EO#��3@�����!?��P��o�@K�5�ٿ���d ��@�EO#��3@�����!?��P��o�@K�5�ٿ���d ��@�EO#��3@�����!?��P��o�@�x�TٙٿlM7{ ��@�l4A��3@I>�܀�!?G����o�@�H�Nr�ٿp� ��@X�W��3@rqOO��!?��	�o�@ý֚ٿ]��� ��@��}���3@�ox��!?1G4�o�@�'�=֚ٿ�M�u ��@�|Y$��3@#�\؏!?N�TA�o�@5���ٿWa�Y ��@-ӗ���3@4P����!?����o�@P%�:Ùٿ�\ ��@�G|  4@"��2y�!?�n���o�@P%�:Ùٿ�\ ��@�G|  4@"��2y�!?�n���o�@h_��ٿP0| ��@�(�o��3@����X�!?�h>�o�@u'))��ٿr-+v ��@(��d��3@��D>k�!?ɨ%�o�@[��ٿC�:v ��@h^"S 4@�e��O�!?≾��o�@���ٿ��� ��@E�`p 4@�yj��!?߽��o�@����̙ٿ�iFL ��@a����3@uן�W�!?��?
�o�@ް"=.�ٿ~� I ��@�	 4@$�p�!?}�E��o�@�"x���ٿ\�B ��@qp>��3@Л|Y�!?�+ ��o�@�"x���ٿ\�B ��@qp>��3@Л|Y�!?�+ ��o�@]��
z�ٿ�cb8 ��@��� 4@��	5.�!? ���o�@Ήu�Øٿ�G% ��@���` 4@C+|�!?Q,���o�@Ήu�Øٿ�G% ��@���` 4@C+|�!?Q,���o�@Ήu�Øٿ�G% ��@���` 4@C+|�!?Q,���o�@�U����ٿ� 2 ��@���� 4@D��w�!? �ͪ�o�@�U����ٿ� 2 ��@���� 4@D��w�!? �ͪ�o�@g��c�ٿ־8 ��@�4����3@R�jh!?U	���o�@H�� �ٿt2G ��@Z�����3@�5\̏!?�¬��o�@��ޒI�ٿ)��( ��@�9J���3@�²*ԏ!?����o�@YLn�ٿ�(����@`����3@	0�۷�!?�v���o�@��~�s�ٿ�eVE ��@7ك���3@�v@��!?�����o�@��~�s�ٿ�eVE ��@7ك���3@�v@��!?�����o�@��~�s�ٿ�eVE ��@7ك���3@�v@��!?�����o�@�Ge�ٿ�N�f ��@����3@ �i ȏ!?۪���o�@�// �ٿ�O<Z ��@)����3@��1U�!?�0�
�o�@�// �ٿ�O<Z ��@)����3@��1U�!?�0�
�o�@�// �ٿ�O<Z ��@)����3@��1U�!?�0�
�o�@�// �ٿ�O<Z ��@)����3@��1U�!?�0�
�o�@`!澐�ٿk��V ��@T�+���3@���~�!?�2�&�o�@�ʹ"֝ٿ'�P ��@A ��3@���wُ!?�$�o�@ԇo`p�ٿ�i ��@@�4X��3@��o
�!?M���o�@ԇo`p�ٿ�i ��@@�4X��3@��o
�!?M���o�@D���ٿ@~ ��@~C����3@�S�9��!?0rΈ�o�@UX˸��ٿ������@�����3@iA#|E�!?�P>�o�@UX˸��ٿ������@�����3@iA#|E�!?�P>�o�@|��]�ٿC�e����@�JG���3@WB�P�!?���h�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@��}�^�ٿ�UM����@��[�3@�"�@�!?y��'�o�@���-�ٿ!~H���@c�� �3@u95�Ǐ!?e]�G�o�@���-�ٿ!~H���@c�� �3@u95�Ǐ!?e]�G�o�@�^Tp�ٿ�������@N���^�3@E�����!? l��o�@�^Tp�ٿ�������@N���^�3@E�����!? l��o�@����ٿp3�����@ցxB��3@�'�N��!?y���o�@6��_�ٿ�G	 ��@z|s���3@;�꜏!?L����o�@6��_�ٿ�G	 ��@z|s���3@;�꜏!?L����o�@6��_�ٿ�G	 ��@z|s���3@;�꜏!?L����o�@6��_�ٿ�G	 ��@z|s���3@;�꜏!?L����o�@6��_�ٿ�G	 ��@z|s���3@;�꜏!?L����o�@�e#\ҙٿ_�~ ��@�<U�  4@bN�!?����o�@�7��ݞٿݧ
' ��@�Ĩֳ�3@30,��!?(� o�o�@�7��ݞٿݧ
' ��@�Ĩֳ�3@30,��!?(� o�o�@�7��ݞٿݧ
' ��@�Ĩֳ�3@30,��!?(� o�o�@]��y`�ٿ�������@6B����3@�Ft�!?](�Z�o�@M��ۘٿ������@L*�: 4@5�]ޏ!?|��d�o�@��ݼ��ٿ��9����@�at���3@W8S�ȏ!?�:���o�@���ٿ������@��]+ 4@T�e��!?��/�o�@���ٿ������@��]+ 4@T�e��!?��/�o�@],|�ؠٿF�&	���@������3@Y�!4�!?Pi6z�o�@],|�ؠٿF�&	���@������3@Y�!4�!?Pi6z�o�@�>̈́��ٿ�]����@dP��3@/��;N�!?���m�o�@����`�ٿ& ����@��<*B�3@#&h�!?�7��o�@�?��̣ٿ�χ����@MrTS�3@X���!?�J���o�@�?��̣ٿ�χ����@MrTS�3@X���!?�J���o�@�?��̣ٿ�χ����@MrTS�3@X���!?�J���o�@�?��̣ٿ�χ����@MrTS�3@X���!?�J���o�@4�8���ٿ؃ͧ���@���F�3@i�o�z�!?�
S��o�@4�8���ٿ؃ͧ���@���F�3@i�o�z�!?�
S��o�@L~�J�ٿ���K���@��9e�3@ͥ��x�!?Pp~��o�@�o��ٿ~�j����@���,��3@3�Z��!?.5���o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@����ݤٿZ����@���:�3@�&�P��!?ÕC�o�@�n(�ٿU{O����@��R��3@�h3�!?�Q
�o�@d���*�ٿ�I����@A�����3@�]\!J�!?�hn��o�@d���*�ٿ�I����@A�����3@�]\!J�!?�hn��o�@����z�ٿs�U����@�S��3@��[PF�!?+�8q�o�@����z�ٿs�U����@�S��3@��[PF�!?+�8q�o�@����z�ٿs�U����@�S��3@��[PF�!?+�8q�o�@7�TTG�ٿ��.z���@�,Lc�3@��a��!?::���o�@7�TTG�ٿ��.z���@�,Lc�3@��a��!?::���o�@7�TTG�ٿ��.z���@�,Lc�3@��a��!?::���o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@�ɸ�êٿZ�F���@ˬk��3@��hΏ!?'08��o�@]���ٿsp\����@�z���3@��z�!?��g�o�@]���ٿsp\����@�z���3@��z�!?��g�o�@]���ٿsp\����@�z���3@��z�!?��g�o�@]���ٿsp\����@�z���3@��z�!?��g�o�@]���ٿsp\����@�z���3@��z�!?��g�o�@]���ٿsp\����@�z���3@��z�!?��g�o�@iO�ٿ͒�(���@��	|��3@��ӹw�!?)����o�@�_���ٿ��4���@�#o-��3@�rH��!?R�oV�o�@�_���ٿ��4���@�#o-��3@�rH��!?R�oV�o�@�_���ٿ��4���@�#o-��3@�rH��!?R�oV�o�@ִ��ٿ�ۓ~���@kI};��3@+Ңux�!?e����o�@�~����ٿ��\���@�{7yW�3@x�琏!?��W��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@'Z��ٿ��ވ���@��:1�3@�k�F�!?)�b��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@��?�ٿj'L����@J�X[��3@����!?ܷa��o�@'�R9��ٿ�Ɂ����@��۱�3@�/L��!?�#�6�o�@'�R9��ٿ�Ɂ����@��۱�3@�/L��!?�#�6�o�@�$L��ٿl��j���@�qF�H�3@0V�(�!?H>��o�@�$L��ٿl��j���@�qF�H�3@0V�(�!?H>��o�@�$L��ٿl��j���@�qF�H�3@0V�(�!?H>��o�@�޿���ٿC�C  ��@(P?��3@|��.�!?tiq+�o�@�޿���ٿC�C  ��@(P?��3@|��.�!?tiq+�o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@f[��
�ٿ������@�@3C�3@S:V�.�!?�97��o�@?�7t]�ٿ~�y ��@����3@r$���!?�Cϯ�o�@?�7t]�ٿ~�y ��@����3@r$���!?�Cϯ�o�@?�7t]�ٿ~�y ��@����3@r$���!?�Cϯ�o�@z����ٿi�)���@�A��P�3@��p��!?"�zt�o�@�����ٿ������@瑏^�3@X+d��!?'����o�@f�&yߝٿ{��k ��@S����3@� ����!?�aa��o�@f�&yߝٿ{��k ��@S����3@� ����!?�aa��o�@����ٿϨ�f���@1�q�3@h� i��!?G҉�o�@����ٿϨ�f���@1�q�3@h� i��!?G҉�o�@����ٿϨ�f���@1�q�3@h� i��!?G҉�o�@����ٿϨ�f���@1�q�3@h� i��!?G҉�o�@����ٿϨ�f���@1�q�3@h� i��!?G҉�o�@�yX6��ٿIP�����@���?��3@��ޏ!?ޥ�*�o�@�yX6��ٿIP�����@���?��3@��ޏ!?ޥ�*�o�@��*T�ٿ2t8���@pzhh��3@݆�{l�!?��+�o�@��*T�ٿ2t8���@pzhh��3@݆�{l�!?��+�o�@�&���ٿ?�Z���@�ݽO��3@	�2۹�!?���d�o�@�&���ٿ?�Z���@�ݽO��3@	�2۹�!?���d�o�@�/��ٿL(����@#�N�-�3@L�Ī@�!?�G"T�o�@�w���ٿVIW��@�w�! 4@DSR�Џ!?!�l��o�@���!{�ٿ�S����@�[W���3@ϋJM�!?H���o�@���+ �ٿ�o�P���@'`ܓ��3@'�=��!?,����o�@���+ �ٿ�o�P���@'`ܓ��3@'�=��!?,����o�@;�j4դٿ��Ύ ��@Hj2�j�3@�Ϙ;a�!?��A��o�@;�j4դٿ��Ύ ��@Hj2�j�3@�Ϙ;a�!?��A��o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@�B%�N�ٿ{�
 ��@AQȥ�3@�_"z�!?#�b�o�@۔��ٿ�]����@$UGp��3@݂5�T�!?U����o�@۔��ٿ�]����@$UGp��3@݂5�T�!?U����o�@۔��ٿ�]����@$UGp��3@݂5�T�!?U����o�@۔��ٿ�]����@$UGp��3@݂5�T�!?U����o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@'�-M۟ٿ*�4u���@�x}m�3@Gck1v�!?�y�5�o�@29����ٿ��a����@j�40��3@i-P(��!?��S�o�@29����ٿ��a����@j�40��3@i-P(��!?��S�o�@M-���ٿ5e)����@�f����3@#h�Ly�!? 1�o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@}PF�>�ٿuUZ���@���'w�3@*+m�Ï!?��e��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��W6�ٿ��J���@o:��3@�����!?��U��o�@��Ry�ٿcH�����@Hl��M�3@bԩۉ�!?��{W�o�@�Ƅŏ�ٿ���0���@`����3@�XV�!?���o�@�!oj�ٿ��<���@�H�?S�3@�Q�2Տ!?P�j��o�@�!oj�ٿ��<���@�H�?S�3@�Q�2Տ!?P�j��o�@C��6>�ٿ	����@���q��3@�h��!?�9! p�@C��6>�ٿ	����@���q��3@�h��!?�9! p�@C��6>�ٿ	����@���q��3@�h��!?�9! p�@�P�ٿ�l�e��@��e��3@K��᥏!?t�D�p�@������ٿ$,��@A�׵[�3@�!��!?f�y
p�@�!���ٿ����@ð�@��3@���-P�!?j-�Dp�@�!���ٿ����@ð�@��3@���-P�!?j-�Dp�@�!���ٿ����@ð�@��3@���-P�!?j-�Dp�@�!���ٿ����@ð�@��3@���-P�!?j-�Dp�@�!���ٿ����@ð�@��3@���-P�!?j-�Dp�@�łF�ٿ���j���@�ka���3@*���!?�_��o�@�łF�ٿ���j���@�ka���3@*���!?�_��o�@�*�@�ٿ��Q����@	p�i�3@
�:��!?�b��p�@�*�@�ٿ��Q����@	p�i�3@
�:��!?�b��p�@��vE~�ٿ��b��@ԍr�S 4@����!?̻���o�@��vE~�ٿ��b��@ԍr�S 4@����!?̻���o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�)�
4�ٿ��%���@�ְ���3@��h�!?�ʜ�o�@�dX+7�ٿ�&%���@�x�c��3@��btv�!?��8��o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@R�H��ٿ��2��@�%o�3@���I1�!?g(c
�o�@._�uͥٿ�^� ��@�$?�e�3@x�L[X�!?@	��o�@w�/��ٿ�Z[` ��@��S��3@�09L�!?[әh�o�@w�/��ٿ�Z[` ��@��S��3@�09L�!?[әh�o�@w�/��ٿ�Z[` ��@��S��3@�09L�!?[әh�o�@w�/��ٿ�Z[` ��@��S��3@�09L�!?[әh�o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@^Eԗ�ٿAk����@i���6 4@�[�C��!?"�q��o�@�7c?��ٿ�cv]��@z�/m�4@�:�M�!?2>��o�@��yGŗٿ�E���@�d�' 4@�p�.�!?����o�@2̞ٿD�B���@��d�;�3@��?��!?γ9p�@2̞ٿD�B���@��d�;�3@��?��!?γ9p�@2̞ٿD�B���@��d�;�3@��?��!?γ9p�@2̞ٿD�B���@��d�;�3@��?��!?γ9p�@2̞ٿD�B���@��d�;�3@��?��!?γ9p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@� �ٿg����@k��Y��3@3
c�z�!?�T�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@c�ySU�ٿψ����@�}mD�3@S��P�!?��z�p�@������ٿi�����@hd����3@�׌��!?��#\p�@�Z~ޙٿ-'����@��J�{�3@����7�!?���p�@���mZ�ٿ9o�C��@� ���3@��Z,�!?B��D/p�@��"2 �ٿ��ם���@�d����3@�OH�!?(��ap�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@���ɞٿhpF����@��Ea�3@�?��!?��f/.p�@~���Οٿ$t����@M�Eӫ�3@�e�t�!?�[��o�@~���Οٿ$t����@M�Eӫ�3@�e�t�!?�[��o�@����ٿ�q� ��@L��� 4@F��R�!?�f#��o�@����ٿ�q� ��@L��� 4@F��R�!?�f#��o�@.�*�3�ٿ�!^l��@�|�hg4@�`a�a�!?�3A�o�@.�*�3�ٿ�!^l��@�|�hg4@�`a�a�!?�3A�o�@.�*�3�ٿ�!^l��@�|�hg4@�`a�a�!?�3A�o�@�Y��ʤٿ/#:%���@y݆{� 4@C�s�8�!?�.~�o�@wZ�,��ٿ4�����@����3@Nh;�!?#0a�o�@wZ�,��ٿ4�����@����3@Nh;�!?#0a�o�@wZ�,��ٿ4�����@����3@Nh;�!?#0a�o�@wZ�,��ٿ4�����@����3@Nh;�!?#0a�o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@��؞ �ٿ4v���@JIL�$ 4@OM�t��!?� ���o�@�2a�w�ٿڴ�K���@��8� 4@[�d�!?�Ӽ�o�@<�A�	�ٿ�Ϋ�߇�@�{�� 4@���|��!?��aՋo�@<�A�	�ٿ�Ϋ�߇�@�{�� 4@���|��!?��aՋo�@bV����ٿ�S8�և�@�.^� 4@�1r�Ï!?r�ׂo�@��+;J�ٿ�d{f͇�@�����3@��6���!?ݢ��o�@��+;J�ٿ�d{f͇�@�����3@��6���!?ݢ��o�@d�}c(�ٿ�iD����@������3@<��Ï!?N*^y�o�@d�}c(�ٿ�iD����@������3@<��Ï!?N*^y�o�@��p ��ٿQm����@U�[�p 4@�[�Xُ!?H���Wo�@��p ��ٿQm����@U�[�p 4@�[�Xُ!?H���Wo�@��p ��ٿQm����@U�[�p 4@�[�Xُ!?H���Wo�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@{�P&�ٿ�߇���@��A4@�ܠ=}�!?pb���o�@X!�<�ٿ�j2҇�@�.��4@�H�x�!?��jo�@X!�<�ٿ�j2҇�@�.��4@�H�x�!?��jo�@f��h�ٿe\{F���@1p��4@���\�!?��5E6o�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@/Jׂ:�ٿz"m����@G^I4@�2�*
�!?C��Ao�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�@=R�ٿGK�Ї�@��0���3@��ϙ��!?��P�o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�n��{�ٿ\T��@�b��3@�ġ�؏!?<B��o�@�W���ٿ9��,��@��Z(� 4@+��ʏ!?qXj&p�@�W���ٿ9��,��@��Z(� 4@+��ʏ!?qXj&p�@�W���ٿ9��,��@��Z(� 4@+��ʏ!?qXj&p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@���2�ٿQ�g7��@��A� 4@�}��L�!?Z��*p�@XP�D�ٿ�bO/��@f�T���3@�=u��!?ji���o�@XP�D�ٿ�bO/��@f�T���3@�=u��!?ji���o�@XP�D�ٿ�bO/��@f�T���3@�=u��!?ji���o�@46SE�ٿ��n�@sUF4@{��K��!?����.o�@46SE�ٿ��n�@sUF4@{��K��!?����.o�@46SE�ٿ��n�@sUF4@{��K��!?����.o�@J.�K�ٿ��ᨇ�@>2���3@g��ڏ!?�:�{o�@J.�K�ٿ��ᨇ�@>2���3@g��ڏ!?�:�{o�@J.�K�ٿ��ᨇ�@>2���3@g��ڏ!?�:�{o�@J.�K�ٿ��ᨇ�@>2���3@g��ڏ!?�:�{o�@�s}�\�ٿt~�,��@�Q�{+�3@�19���!?9�b��p�@�s}�\�ٿt~�,��@�Q�{+�3@�19���!?9�b��p�@5���o�ٿ�C�Q��@�'#��3@�V��K�!?�3g�p�@F3��ٿn��=N��@���3@�gU7�!?��9̶p�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@���f^�ٿ͇
��@�X�^g�3@��m��!?&6���q�@r�$d��ٿ��@O��@0�eK��3@�#h�ˏ!?&|�;xp�@r�$d��ٿ��@O��@0�eK��3@�#h�ˏ!?&|�;xp�@r�$d��ٿ��@O��@0�eK��3@�#h�ˏ!?&|�;xp�@r�$d��ٿ��@O��@0�eK��3@�#h�ˏ!?&|�;xp�@]c�Zg�ٿ����m��@Ō��3@ꦠ ُ!?�?/g�n�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@�̣�L�ٿ�����@�3n̘�3@���!?O����p�@��	��ٿM��W��@Cܞ?4@�)��X�!?�d� Zp�@��	��ٿM��W��@Cܞ?4@�)��X�!?�d� Zp�@��	��ٿM��W��@Cܞ?4@�)��X�!?�d� Zp�@'�מٿ��eA��@�|��4@�-тR�!?�Wo@�n�@'�מٿ��eA��@�|��4@�-тR�!?�Wo@�n�@'�מٿ��eA��@�|��4@�-тR�!?�Wo@�n�@'�מٿ��eA��@�|��4@�-тR�!?�Wo@�n�@6p4�Ңٿ�'ۇ�@ѳ�@�4@����!?݉lo�@6p4�Ңٿ�'ۇ�@ѳ�@�4@����!?݉lo�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@IC#!e�ٿS.�;���@vV�a��3@��?X�!?��1��p�@�5s�ٿ�Ƒdr��@�)2���3@P���!?�-�I�p�@�5s�ٿ�Ƒdr��@�)2���3@P���!?�-�I�p�@�5s�ٿ�Ƒdr��@�)2���3@P���!?�-�I�p�@�5s�ٿ�Ƒdr��@�)2���3@P���!?�-�I�p�@�5s�ٿ�Ƒdr��@�)2���3@P���!?�-�I�p�@��^�ٿ1��^��@����'4@}���!?�+��n�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@3���a�ٿ� �j��@&�WF{4@zQS��!? ��6xn�@�ޥ�ٿ����{��@�F) 4@���/��!?T�)F}n�@�ޥ�ٿ����{��@�F) 4@���/��!?T�)F}n�@�ޥ�ٿ����{��@�F) 4@���/��!?T�)F}n�@P��`ߗٿ��'J��@��d�k4@��_�!?I��
�o�@P��`ߗٿ��'J��@��d�k4@��_�!?I��
�o�@�m�ٿvd^Ї�@�d�4@
|�V��!?"ٺk�n�@�m�ٿvd^Ї�@�d�4@
|�V��!?"ٺk�n�@�m�ٿvd^Ї�@�d�4@
|�V��!?"ٺk�n�@���ٿ^P����@��_�4@w�(�!?"���4o�@;�$ϧٿ?K����@TH�	4@Ԙ"?h�!?`s��$o�@;�$ϧٿ?K����@TH�	4@Ԙ"?h�!?`s��$o�@;�$ϧٿ?K����@TH�	4@Ԙ"?h�!?`s��$o�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@���\_�ٿA3P���@�W��4@�����!?���vvl�@Ub{Y��ٿ��!F��@j��p�4@�!E!?v�Vqbm�@����l�ٿ4a�L��@B�a4@o��(Ə!?�/R^p�@����l�ٿ4a�L��@B�a4@o��(Ə!?�/R^p�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�1ҟٿ��s��@��\R��3@��v���!?Ͳ��q�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@�~ѧٿO���{��@K�mk��3@Y)��u�!?\��6�o�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@vW̈�ٿ�4���@�]�� 4@����!?yDҊo�@>�=y�ٿ��H�[��@��
��3@�4�zj�!?����lp�@z��$�ٿL&�WQ��@ YZ6��3@(R�@��!?�#�ap�@z��$�ٿL&�WQ��@ YZ6��3@(R�@��!?�#�ap�@ȝ7ƫٿ%kb��@�����3@�?NV��!?	d���o�@ȝ7ƫٿ%kb��@�����3@�?NV��!?	d���o�@F�D[w�ٿp�ԝ��@5�rz� 4@�Lƛh�!? A߀o�@F�D[w�ٿp�ԝ��@5�rz� 4@�Lƛh�!? A߀o�@���Q�ٿeG.⇈�@Qma�3@�hPF�!?:��`lp�@�d��ٿ9$�ϥ��@"˂o�4@9��2��!?�yʟo�@�d��ٿ9$�ϥ��@"˂o�4@9��2��!?�yʟo�@�d��ٿ9$�ϥ��@"˂o�4@9��2��!?�yʟo�@��a��ٿ�c̒���@��Z�4@+0JM��!?��m�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@���)W�ٿ/��~��@M�P4@Hȏ��!?YC?�k�@�O�{P�ٿ1����@�hJ4@wg1�L�!?@.��l�@�O�{P�ٿ1����@�hJ4@wg1�L�!?@.��l�@�O�{P�ٿ1����@�hJ4@wg1�L�!?@.��l�@�O�{P�ٿ1����@�hJ4@wg1�L�!?@.��l�@�6C��ٿ�U7���@������3@��ܤϏ!?�IMoEo�@�6C��ٿ�U7���@������3@��ܤϏ!?�IMoEo�@�6C��ٿ�U7���@������3@��ܤϏ!?�IMoEo�@�6C��ٿ�U7���@������3@��ܤϏ!?�IMoEo�@��1�ٿ8��S���@/.*��4@�����!?��@Al�@�IT��ٿ �h���@���c�4@��ykg�!?D���n�@�IT��ٿ �h���@���c�4@��ykg�!?D���n�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��ٿ�kr���@����; 4@$hɏ!?JV�q�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@��m{�ٿ�n�W��@"�RŚ4@pѥ�!?5(��m�@�%`�ٿ��CJ��@#�4��3@�$�ӏ!?��¿�o�@�%`�ٿ��CJ��@#�4��3@�$�ӏ!?��¿�o�@�%`�ٿ��CJ��@#�4��3@�$�ӏ!?��¿�o�@�%`�ٿ��CJ��@#�4��3@�$�ӏ!?��¿�o�@�%`�ٿ��CJ��@#�4��3@�$�ӏ!?��¿�o�@�@�\�ٿ G&ᦈ�@6t�n�4@�5��J�!?V�W�o�@�@�\�ٿ G&ᦈ�@6t�n�4@�5��J�!?V�W�o�@�K��0�ٿp��2���@ŧ � 4@?g���!?ϓ.�r�@�K��0�ٿp��2���@ŧ � 4@?g���!?ϓ.�r�@�K��0�ٿp��2���@ŧ � 4@?g���!?ϓ.�r�@�K��0�ٿp��2���@ŧ � 4@?g���!?ϓ.�r�@����ٿ~$�ᝈ�@m��,4@|gƥ�!?�]�p�@éB��ٿ��آ��@|;�= 4@��'܏!?aI��k�@�X���ٿCg�����@��T4@3�lǏ!?�E��k�@�%W��ٿ}�~���@tL q��3@�\O���!?��W��l�@�%W��ٿ}�~���@tL q��3@�\O���!?��W��l�@��i�֩ٿ�<��*��@���64@0�C���!?��l�l�@��i�֩ٿ�<��*��@���64@0�C���!?��l�l�@��i�֩ٿ�<��*��@���64@0�C���!?��l�l�@��i�֩ٿ�<��*��@���64@0�C���!?��l�l�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@��0�n�ٿu&�
���@	V��4@�K�Y�!?$�-�q�@-���ٿ�x7��@�Fcw�4@{�ߐC�!?wmh�r�@-���ٿ�x7��@�Fcw�4@{�ߐC�!?wmh�r�@8%�ɥٿ"ҫ��@�R�U�3@�� ��!?�4e#q�@8%�ɥٿ"ҫ��@�R�U�3@�� ��!?�4e#q�@u6�
�ٿ���
/��@�_$/{ 4@>rk��!?�L�j�@u6�
�ٿ���
/��@�_$/{ 4@>rk��!?�L�j�@u6�
�ٿ���
/��@�_$/{ 4@>rk��!?�L�j�@�v�u��ٿk���@�P^��3@X�w?t�!?�3���q�@�v�u��ٿk���@�P^��3@X�w?t�!?�3���q�@�v�u��ٿk���@�P^��3@X�w?t�!?�3���q�@�v�u��ٿk���@�P^��3@X�w?t�!?�3���q�@]�G'��ٿ\� oƊ�@��'��3@�d��Ώ!?p����q�@]�G'��ٿ\� oƊ�@��'��3@�d��Ώ!?p����q�@]�G'��ٿ\� oƊ�@��'��3@�d��Ώ!?p����q�@u�� ��ٿ��'i���@�}��4@hC:�!?��^%/k�@u�� ��ٿ��'i���@�}��4@hC:�!?��^%/k�@u�� ��ٿ��'i���@�}��4@hC:�!?��^%/k�@u�� ��ٿ��'i���@�}��4@hC:�!?��^%/k�@u�� ��ٿ��'i���@�}��4@hC:�!?��^%/k�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@7_&3�ٿQ\6��@��@j4@���{,�!?Oώ�.i�@��P��ٿ�39#h��@ğ+4@�(�+�!? �nCf�@��P��ٿ�39#h��@ğ+4@�(�+�!? �nCf�@��P��ٿ�39#h��@ğ+4@�(�+�!? �nCf�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�H�eޠٿ��<����@7�7a�3@�DՖ0�!?**~�f�@�u�WX�ٿǙK,��@�nKa 4@b1���!?�����b�@�u�WX�ٿǙK,��@�nKa 4@b1���!?�����b�@�u�WX�ٿǙK,��@�nKa 4@b1���!?�����b�@�u�WX�ٿǙK,��@�nKa 4@b1���!?�����b�@]u��ٿ�*q�@+��9u�3@�e��-�!?��QO�S�@]u��ٿ�*q�@+��9u�3@�e��-�!?��QO�S�@]u��ٿ�*q�@+��9u�3@�e��-�!?��QO�S�@]u��ٿ�*q�@+��9u�3@�e��-�!?��QO�S�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�����ٿ��%Y��@���F4@��~p��!?)�i�_b�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@�p,ԗ�ٿ@�g*���@P��s 4@��&X'�!?S�^a\�@J��I�ٿ���K���@��W�;�3@=��z��!?�Zywa�@J��I�ٿ���K���@��W�;�3@=��z��!?�Zywa�@J��I�ٿ���K���@��W�;�3@=��z��!?�Zywa�@J��I�ٿ���K���@��W�;�3@=��z��!?�Zywa�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@���G�ٿ�+�*�@�=�U��3@�w�mŏ!?�h
��a�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�.�3�ٿT��<���@�׬4@v�ycI�!?�ǳ�Hn�@�|@u�ٿ��W��@�$�h4@�����!?Ln�F-l�@�|@u�ٿ��W��@�$�h4@�����!?Ln�F-l�@1���ٿ������@_�� 4@PC?��!?��o�U}�@1���ٿ������@_�� 4@PC?��!?��o�U}�@��1耛ٿ�aʲ~�@��4@x~����!?�-�x:z�@��1耛ٿ�aʲ~�@��4@x~����!?�-�x:z�@��1耛ٿ�aʲ~�@��4@x~����!?�-�x:z�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@P��g�ٿM'��{�@�5ٳ� 4@e�����!?Z*�20}�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@�����ٿ6i&�#x�@�C�� 4@]9P���!?���'�p�@���7��ٿ�B��s�@;�ѯ/�3@�=��!?\�����@���7��ٿ�B��s�@;�ѯ/�3@�=��!?\�����@���7��ٿ�B��s�@;�ѯ/�3@�=��!?\�����@���7��ٿ�B��s�@;�ѯ/�3@�=��!?\�����@�"�
�ٿ[j���w�@��xE 4@(w-n��!?>'ˣw�@�"�
�ٿ[j���w�@��xE 4@(w-n��!?>'ˣw�@�"�
�ٿ[j���w�@��xE 4@(w-n��!?>'ˣw�@�"�
�ٿ[j���w�@��xE 4@(w-n��!?>'ˣw�@��`W֜ٿr�pij}�@+ I74@ �f�!?L��8q�@3�f>7�ٿ��>ɀ�@(d��)4@�/\v��!?�a�K�w�@3�f>7�ٿ��>ɀ�@(d��)4@�/\v��!?�a�K�w�@�%3��ٿ��y�ց�@w��P�3@u�	#ڏ!?����XR�@�%3��ٿ��y�ց�@w��P�3@u�	#ڏ!?����XR�@�%3��ٿ��y�ց�@w��P�3@u�	#ڏ!?����XR�@�%3��ٿ��y�ց�@w��P�3@u�	#ڏ!?����XR�@g��A�ٿ2��{�@|�<p��3@�{d"�!?ѯ&�[B�@g��A�ٿ2��{�@|�<p��3@�{d"�!?ѯ&�[B�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@��$O�ٿ�h1^�@Ŝ�F 4@Y��Ώ!?e��e�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@:���§ٿ	?�iՇ�@�9��+�3@<[؊�!?��,�@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���v��ٿ"#�U��@��丒�3@q��Uw�!?�6a5A��@���x�ٿ��B����@V�t�3@�_r�!?��z�A��@���x�ٿ��B����@V�t�3@�_r�!?��z�A��@���x�ٿ��B����@V�t�3@�_r�!?��z�A��@���x�ٿ��B����@V�t�3@�_r�!?��z�A��@���x�ٿ��B����@V�t�3@�_r�!?��z�A��@'TXa�ٿ�Q4@$��@��Y���3@�X�.�!?f?d¤��@'TXa�ٿ�Q4@$��@��Y���3@�X�.�!?f?d¤��@'TXa�ٿ�Q4@$��@��Y���3@�X�.�!?f?d¤��@u},&�ٿ�D��9��@B��D��3@7q�m�!?�CWY��@�����ٿB;zq��@�#b���3@�6DY܏!? W�$j��@�����ٿB;zq��@�#b���3@�6DY܏!? W�$j��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@���F�ٿ��܋��@�T�3��3@�5G��!?��zP��@\�G�ٿ=�lΘ�@����.�3@l�؏!?��?��@\�G�ٿ=�lΘ�@����.�3@l�؏!?��?��@\�G�ٿ=�lΘ�@����.�3@l�؏!?��?��@G?�_�ٿͩ�ަ�@q�O�+�3@��	��!?Y�f�s�@G?�_�ٿͩ�ަ�@q�O�+�3@��	��!?Y�f�s�@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@��=�ٿ՜]�f��@��dcN�3@�G��!?��2���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@f]��ٿ�]��ٜ�@l���z�3@98�o��!?�,�_���@�H�U��ٿ����@#��+�3@׼-��!?s���@�@�H�U��ٿ����@#��+�3@׼-��!?s���@�@T<�̋ٿe�j���@�*\#�3@z2c狏!?�8y
�@T<�̋ٿe�j���@�*\#�3@z2c狏!?�8y
�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@�D���ٿ��˸�@T�=*�3@�{�!?&�'?ZP�@9�[.2�ٿ����Ų�@��l��3@:<�p�!?>���,�@9�[.2�ٿ����Ų�@��l��3@:<�p�!?>���,�@9�[.2�ٿ����Ų�@��l��3@:<�p�!?>���,�@9�[.2�ٿ����Ų�@��l��3@:<�p�!?>���,�@WR��ٿ
���6��@
�P�"�3@.J�Ri�!?H���
K�@WR��ٿ
���6��@
�P�"�3@.J�Ri�!?H���
K�@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@Ry:�ߧٿ �v��@~u�C��3@�c�݃�!?&�����@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@������ٿ����ө�@U��� 4@����}�!?��J]��@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@��w���ٿڣ�O`��@�
3g 4@���2�!?�����@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@K ��ٿ�����@5CF9��3@`�NNG�!?d(߲�@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@ab7ٿ�:�_O��@㤟�=4@a�~;��!?t°.��@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�'���ٿ��x/���@�o���4@��@�{�!?�w9p�B�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@�bÜٿx��
*��@M�9H14@G�վԏ!?�,��r�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���H�ٿ��u�h��@�ͬH4@SɾRg�!? �M�@���/�ٿ������@�W>W� 4@���Eu�!?���(۩�@O��7�ٿ�3�x��@?!��� 4@H��!x�!?��ɣ�a�@O��7�ٿ�3�x��@?!��� 4@H��!x�!?��ɣ�a�@O��7�ٿ�3�x��@?!��� 4@H��!x�!?��ɣ�a�@O��7�ٿ�3�x��@?!��� 4@H��!x�!?��ɣ�a�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@5�aH:�ٿri����@W�j4@'A��g�!?�j�o�@��P��ٿj���t��@}6��� 4@��y{�!?�@����@��P��ٿj���t��@}6��� 4@��y{�!?�@����@��P��ٿj���t��@}6��� 4@��y{�!?�@����@��P��ٿj���t��@}6��� 4@��y{�!?�@����@T4��i�ٿ��g��@�A�I��3@Ų|³�!?,���C�@T4��i�ٿ��g��@�A�I��3@Ų|³�!?,���C�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@"Up��ٿk��|&��@C�[�� 4@�c���!?�� I�@�v2ǣ�ٿL���E��@�bv}4@��<���!?�
B���@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@Z�=ܨٿ������@�,� 4@H��F��!?���a$y�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@�Bz�ӜٿlNz�׺�@N]脐 4@k�0��!?�D��j�@����ٿ'w�;���@a�)�� 4@��d�G�!?[�����@����ٿ'w�;���@a�)�� 4@��d�G�!?[�����@����ٿ'w�;���@a�)�� 4@��d�G�!?[�����@�~	p��ٿ�9_��@���4@W�!���!?^1����@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@(� �ٿ&us����@S �%� 4@�>���!?G�$���@:��s��ٿQZt��@�?��"4@X��<��!?�y��@:��s��ٿQZt��@�?��"4@X��<��!?�y��@:��s��ٿQZt��@�?��"4@X��<��!?�y��@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@��J3�ٿê�����@��6,� 4@�F��T�!?���M���@�Y�Ik�ٿЏ�!��@@F#C�4@�V�g��!?����8�@�Y�Ik�ٿЏ�!��@@F#C�4@�V�g��!?����8�@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�m3"�ٿ���b��@�%�V� 4@�9,��!?��<h��@�!i�ޥٿĄZ%���@��� 4@�3���!?R���]�@�!i�ޥٿĄZ%���@��� 4@�3���!?R���]�@/f�H�ٿ��f�i��@�K^� 4@��D���!?�]�G7�@/f�H�ٿ��f�i��@�K^� 4@��D���!?�]�G7�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@�N89�ٿ��?��@iG�!~�3@Nj��!?}-.[	E�@O"��ٿ������@9/�U��3@�;$��!?���H�j�@ß�TY�ٿ��a(Ƭ�@�}fg��3@/�G=�!?�\*�b&�@�BM�'�ٿW.�#y�@�f5�3@��-�!?��g�{��@�nū�ٿ�B�ڭq�@�Z�U�3@[�mˮ�!?�O�Z��@�nū�ٿ�B�ڭq�@�Z�U�3@[�mˮ�!?�O�Z��@�e�
��ٿ5��L��@/��3� 4@ }����!?�"zVC�@�]H�Ůٿ�þc�@�y�4@Æ��{�!?;�\^��@�]H�Ůٿ�þc�@�y�4@Æ��{�!?;�\^��@�]H�Ůٿ�þc�@�y�4@Æ��{�!?;�\^��@�]H�Ůٿ�þc�@�y�4@Æ��{�!?;�\^��@�]H�Ůٿ�þc�@�y�4@Æ��{�!?;�\^��@d^�g��ٿ��n��q�@�m;	34@��q|��!?Ɯ$���@d^�g��ٿ��n��q�@�m;	34@��q|��!?Ɯ$���@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@��Q�ٿ��6��@��4@F�*W�!?��3�Q,�@ug�K�ٿ7q$fl�@�RCj��3@奾��!?�����@ug�K�ٿ7q$fl�@�RCj��3@奾��!?�����@ug�K�ٿ7q$fl�@�RCj��3@奾��!?�����@�Tn`�ٿ��齖�@���`j�3@ni9渏!?���s3��@�Tn`�ٿ��齖�@���`j�3@ni9渏!?���s3��@�Tn`�ٿ��齖�@���`j�3@ni9渏!?���s3��@�Tn`�ٿ��齖�@���`j�3@ni9渏!?���s3��@�Tn`�ٿ��齖�@���`j�3@ni9渏!?���s3��@)�HèٿAW�"ˍ�@=�w�D 4@�,��!?!}(���@)�HèٿAW�"ˍ�@=�w�D 4@�,��!?!}(���@)�HèٿAW�"ˍ�@=�w�D 4@�,��!?!}(���@
C��ٿX��N��@�x@H 4@ *g�e�!?�$.�G��@
C��ٿX��N��@�x@H 4@ *g�e�!?�$.�G��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@��L?�ٿ�0��9��@���#��3@ĭ.�Ώ!?��J�b��@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@���K�ٿ�o�x��@�+���3@��؆�!?/�O���@�d�=V�ٿ�b���@��Q 4@ra� `�!?�Οf�9�@��u��ٿ�2*����@���p4@&��g�!?m��yH�@��u��ٿ�2*����@���p4@&��g�!?m��yH�@��u��ٿ�2*����@���p4@&��g�!?m��yH�@�*ǐs�ٿ�r��@*��t�4@��-�`�!?��]a��@O�.���ٿh�%���@�����3@��@H��!?̦&Q\�@O�.���ٿh�%���@�����3@��@H��!?̦&Q\�@�
� 7�ٿCb�R��@7�4w�3@����`�!?{��<'�@�
� 7�ٿCb�R��@7�4w�3@����`�!?{��<'�@�
� 7�ٿCb�R��@7�4w�3@����`�!?{��<'�@�
� 7�ٿCb�R��@7�4w�3@����`�!?{��<'�@�
� 7�ٿCb�R��@7�4w�3@����`�!?{��<'�@jw��v�ٿH��`v�@�M��O 4@/�i�i�!?�8㨈��@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@ߝ �ٿ�9#��p�@r�*�4@�{��f�!?`V��c%�@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@"�߉F�ٿ��B�w�@@
�.4@k|��l�!?h�{��@*LT���ٿޡ=���@r�l� 4@x=�]�!?zn���@=Ze�0�ٿr����@�g�ct4@`���!?p�b�y[�@=Ze�0�ٿr����@�g�ct4@`���!?p�b�y[�@����ٿBL6����@y*}]� 4@����!?�s�&K�@����ٿBL6����@y*}]� 4@����!?�s�&K�@����ٿBL6����@y*}]� 4@����!?�s�&K�@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@2S����ٿ��9����@=�K<-�3@a��e|�!?g=���@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@/e&�,�ٿ30��f�@��PY� 4@+b8w�!?rP��S[�@��O�\�ٿE=7�j��@�gg��3@�=NѰ�!?�GKB��@��O�\�ٿE=7�j��@�gg��3@�=NѰ�!?�GKB��@��O�\�ٿE=7�j��@�gg��3@�=NѰ�!?�GKB��@��O�\�ٿE=7�j��@�gg��3@�=NѰ�!?�GKB��@v�Y��ٿ���Ԑ�@��<��3@;�̽�!?�^���@v�Y��ٿ���Ԑ�@��<��3@;�̽�!?�^���@/��x˲ٿ��с=��@�����3@uPy��!?3(���A�@/��x˲ٿ��с=��@�����3@uPy��!?3(���A�@������ٿ��+:��@RB���3@� �֏!?�~^�F(�@������ٿ��+:��@RB���3@� �֏!?�~^�F(�@������ٿ��+:��@RB���3@� �֏!?�~^�F(�@H�y��ٿ]Z����@�.r1� 4@T���!?� ��2��@H�y��ٿ]Z����@�.r1� 4@T���!?� ��2��@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@$~ƈ�ٿ=[~e@��@�l��A�3@ܤU���!?������@�?x,�ٿش^+���@�3��� 4@|qP���!?��d����@�?x,�ٿش^+���@�3��� 4@|qP���!?��d����@�?x,�ٿش^+���@�3��� 4@|qP���!?��d����@�?x,�ٿش^+���@�3��� 4@|qP���!?��d����@�?x,�ٿش^+���@�3��� 4@|qP���!?��d����@��~��ٿ�)Y�{�@�>���4@oF�y��!?u�h�p�@��~��ٿ�)Y�{�@�>���4@oF�y��!?u�h�p�@��~��ٿ�)Y�{�@�>���4@oF�y��!?u�h�p�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@�*��ٿ�!�0Ҥ�@����� 4@����s�!?��!�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@}��VO�ٿޝ5����@X)��Q4@欰�y�!?���0M9�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@0�ׄ�ٿ�f6���@��F\4@M�?�x�!?�|�d�	�@[����ٿ�&ѭ�@n��"4@7Z��!?C�A*ہ�@[����ٿ�&ѭ�@n��"4@7Z��!?C�A*ہ�@[����ٿ�&ѭ�@n��"4@7Z��!?C�A*ہ�@[����ٿ�&ѭ�@n��"4@7Z��!?C�A*ہ�@w��5��ٿ|ks���@�?_� 4@n��@��!?n��)��@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@��f*b�ٿ郜�1��@Fr��4@���T�!?�:j��&�@]v��ٿ��c�u�@�{Gs 4@:��`�!? �bx�@]v��ٿ��c�u�@�{Gs 4@:��`�!? �bx�@]v��ٿ��c�u�@�{Gs 4@:��`�!? �bx�@d]�;R�ٿ�׼��@��Y!4@�<P�b�!?'<7�e��@d]�;R�ٿ�׼��@��Y!4@�<P�b�!?'<7�e��@d]�;R�ٿ�׼��@��Y!4@�<P�b�!?'<7�e��@�.c�ٿ��b;du�@�f�4@�T�Oڏ!?����g�@�.c�ٿ��b;du�@�f�4@�T�Oڏ!?����g�@�����ٿK�GA{�@����[�3@�}���!?��^�3�@�����ٿK�GA{�@����[�3@�}���!?��^�3�@ǴU
�ٿ�GF�u��@�ڵÎ4@��я!?�,��<I�@ǴU
�ٿ�GF�u��@�ڵÎ4@��я!?�,��<I�@8� g��ٿqgƛ�@���M 4@a��!?�o�:��@8� g��ٿqgƛ�@���M 4@a��!?�o�:��@8� g��ٿqgƛ�@���M 4@a��!?�o�:��@�n4q��ٿ#	����@��u9f�3@�n���!?h-����@�n4q��ٿ#	����@��u9f�3@�n���!?h-����@�n4q��ٿ#	����@��u9f�3@�n���!?h-����@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@j�>@�ٿ�fO���@�!n���3@O�O���!?-�Q�r�@�;{]�ٿ����ω�@n�~�n�3@ O�ˏ!?>�����@C��ٿ��+G��@6R�͚�3@�<�lҏ!?͌�[�%�@C��ٿ��+G��@6R�͚�3@�<�lҏ!?͌�[�%�@C��ٿ��+G��@6R�͚�3@�<�lҏ!?͌�[�%�@C��ٿ��+G��@6R�͚�3@�<�lҏ!?͌�[�%�@C��ٿ��+G��@6R�͚�3@�<�lҏ!?͌�[�%�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@l�J
Ϟٿ@Jɕ"1�@i��: 4@J٤䲏!?)[��U�@4 ���ٿ���+@�@�5�%�3@g�R��!?F�\���@4 ���ٿ���+@�@�5�%�3@g�R��!?F�\���@4 ���ٿ���+@�@�5�%�3@g�R��!?F�\���@4 ���ٿ���+@�@�5�%�3@g�R��!?F�\���@Wr��ٿ3yr>P�@CЛ��3@`u�!?޿�t��@Wr��ٿ3yr>P�@CЛ��3@`u�!?޿�t��@Wr��ٿ3yr>P�@CЛ��3@`u�!?޿�t��@�Q4t��ٿ>�w�R�@��q��3@�k衏�!?wT@�_�@�!��-�ٿ�kP
*�@/hy���3@�2}�_�!?�g�����@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@e�c��ٿ���	{�@@�]���3@��Jv�!?}x��T�@N����ٿ���G�@���pw�3@�Wc|��!?�K��g�@N����ٿ���G�@���pw�3@�Wc|��!?�K��g�@A�:�!�ٿA����@���/4@F�?G�!?j���@A�:�!�ٿA����@���/4@F�?G�!?j���@A�:�!�ٿA����@���/4@F�?G�!?j���@�?��ٿRV����@n�ʀ�4@�\`J��!?~���	�@�?��ٿRV����@n�ʀ�4@�\`J��!?~���	�@t���ٿ�3_�I��@�>w�]�3@|g��Ï!?Y���a�@t���ٿ�3_�I��@�>w�]�3@|g��Ï!?Y���a�@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@Q�����ٿ�u5���@�v���3@��3r�!?�?�9��@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@��-R��ٿVx�k0M�@<�$���3@�����!?:�Oj�@�HA�f�ٿ f�8Sl�@�J��3@gR�\x�!?C�����@�HA�f�ٿ f�8Sl�@�J��3@gR�\x�!?C�����@�HA�f�ٿ f�8Sl�@�J��3@gR�\x�!?C�����@�HA�f�ٿ f�8Sl�@�J��3@gR�\x�!?C�����@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@�CC��ٿƞ:2{t�@DjYZ��3@�w��!?-CCE�~�@����ٿ� 07l�@� �= 4@t��ay�!?���XA�@�+i)Y�ٿ�;���@��8��3@��Zv�!?RV����@�+i)Y�ٿ�;���@��8��3@��Zv�!?RV����@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@�i���ٿARGfq�@�|����3@=��vǏ!?Zp��(��@��՜ٿ�Ҁ�r��@ FT� 4@�k�a�!?ܸ�:v��@��՜ٿ�Ҁ�r��@ FT� 4@�k�a�!?ܸ�:v��@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@rQҪH�ٿN/�6%��@�~��4@�Ə�Q�!?��%�%�@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@!�n&�ٿ;�e��@��z�4@�[1��!?�<�����@d=<�ٿ��.�@�xD#4@u���m�!?B�r�+��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@!�}��ٿ�{�Ny�@�J54@���r�!?�l)�h��@���ߑ�ٿ��B�K�@/�8�H4@�\=�!?���+���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��a�ٿ"�r�r��@�0=Z4@M� �0�!?d$���@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@��S��ٿ�* �[�@}a��H4@(�.�	�!?��d�.��@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@gx���ٿ#�Ѝ�%�@��9���3@H˨팏!?��'u[M�@p�]R�ٿ�cGw���@̨��3@an��c�!?+ff$։�@p�]R�ٿ�cGw���@̨��3@an��c�!?+ff$։�@p�]R�ٿ�cGw���@̨��3@an��c�!?+ff$։�@p�]R�ٿ�cGw���@̨��3@an��c�!?+ff$։�@p�]R�ٿ�cGw���@̨��3@an��c�!?+ff$։�@�l����ٿm��A��@1����3@�a����!?������@�l����ٿm��A��@1����3@�a����!?������@�l����ٿm��A��@1����3@�a����!?������@�l����ٿm��A��@1����3@�a����!?������@�l����ٿm��A��@1����3@�a����!?������@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@w'��*�ٿ�g '�X�@9����3@�k�y�!?w��m�@�I�r��ٿ���V��@��ΔR�3@�u�pv�!?�^���@�I�r��ٿ���V��@��ΔR�3@�u�pv�!?�^���@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�N'�ٿ�����w�@]}v��3@VR74��!?)ˈs�@�pݜٿ����n�@�7J�3@�v'!ԏ!?��b�a��@�pݜٿ����n�@�7J�3@�v'!ԏ!?��b�a��@�pݜٿ����n�@�7J�3@�v'!ԏ!?��b�a��@�Y�%ѩٿ�XZ���@�%!%�3@G��p��!?�ɡ�5��@�Y�%ѩٿ�XZ���@�%!%�3@G��p��!?�ɡ�5��@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@��-��ٿw�a�S��@��	4@����!?M�����@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@�:�S�ٿ���MY��@K�ȋS�3@�RY��!?$�W��@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@���m�ٿ)��B؏�@�G1L� 4@��R��!?[����}�@�2�7ɤٿm������@���
��3@Zl��!?�2:��;�@K���ٿ?R����@y�����3@���Ϗ!?����l��@K���ٿ?R����@y�����3@���Ϗ!?����l��@��1I�ٿ��7���@�Mŝ4@C��[�!?�O@��-�@��1I�ٿ��7���@�Mŝ4@C��[�!?�O@��-�@��1I�ٿ��7���@�Mŝ4@C��[�!?�O@��-�@dT���ٿ^ly{�@5[١Y4@"�`��!?��O�m$�@dT���ٿ^ly{�@5[١Y4@"�`��!?��O�m$�@dT���ٿ^ly{�@5[١Y4@"�`��!?��O�m$�@��^�F�ٿ_�t���@�~��3@��:ߴ�!?&@ϫ_��@��^�F�ٿ_�t���@�~��3@��:ߴ�!?&@ϫ_��@��^�F�ٿ_�t���@�~��3@��:ߴ�!?&@ϫ_��@��^�F�ٿ_�t���@�~��3@��:ߴ�!?&@ϫ_��@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@k��.(�ٿ�A�cy�@\,�T!4@K�2���!?d�<��O�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@�Z���ٿ�rv@�@��;0 4@OY�u��!?(]�8�@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@g�m"�ٿ��x~��@�ۻ� 4@�m�I�!?�m����@-U:D��ٿ�B4���@>��&� 4@�q�,�!?EV�`��@-U:D��ٿ�B4���@>��&� 4@�q�,�!?EV�`��@-U:D��ٿ�B4���@>��&� 4@�q�,�!?EV�`��@-U:D��ٿ�B4���@>��&� 4@�q�,�!?EV�`��@-U:D��ٿ�B4���@>��&� 4@�q�,�!?EV�`��@D1��!�ٿ�����@��F� 4@��>Zs�!?�b��m�@D1��!�ٿ�����@��F� 4@��>Zs�!?�b��m�@�]�ٿP�dYu��@�L��4 4@�$e���!?9-�\� �@�]�ٿP�dYu��@�L��4 4@�$e���!?9-�\� �@�]�ٿP�dYu��@�L��4 4@�$e���!?9-�\� �@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@y��|��ٿf��*���@��mv4@u��w�!?���D7%�@��m�ٿ��Zu�:�@2{1�4@6�䉁�!?qrC�V�@��m�ٿ��Zu�:�@2{1�4@6�䉁�!?qrC�V�@��m�ٿ��Zu�:�@2{1�4@6�䉁�!?qrC�V�@��m�ٿ��Zu�:�@2{1�4@6�䉁�!?qrC�V�@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@b45�ٿ�N�����@��4�4@�Ԅ���!?+�	f��@�����ٿYP�Ko��@a���4@v0�R��!?�4���@�zE���ٿ~�����@��r���3@�L�1�!?2�U��@�zE���ٿ~�����@��r���3@�L�1�!?2�U��@g~�\�ٿx�d��@�lA�� 4@�T���!?�Uh"J�@g~�\�ٿx�d��@�lA�� 4@�T���!?�Uh"J�@g~�\�ٿx�d��@�lA�� 4@�T���!?�Uh"J�@�5��ٿ3N���@D�Q��4@�@���!?/��}�s�@�5��ٿ3N���@D�Q��4@�@���!?/��}�s�@�5��ٿ3N���@D�Q��4@�@���!?/��}�s�@�5��ٿ3N���@D�Q��4@�@���!?/��}�s�@�5��ٿ3N���@D�Q��4@�@���!?/��}�s�@�H`�ٿ�߻���@Q��с 4@$�����!?o0����@�H`�ٿ�߻���@Q��с 4@$�����!?o0����@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@��ٿ=q����@[�-�z 4@' 0z��!?T*�}��@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@& ņ�ٿ�NHl���@�����3@$l2@r�!?�=K%�M�@iTbR�ٿͺ�����@��!� 4@H/U3^�!?��E����@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�l�S~�ٿ�%%S��@����� 4@ٹFB��!?��c��d�@�B�Ϧٿ^��-�@r<�S4@�8��!?5�+V{�@ugP��ٿ�'߾��@O�Z4@�f�⤏!?�9�8�(�@ugP��ٿ�'߾��@O�Z4@�f�⤏!?�9�8�(�@ugP��ٿ�'߾��@O�Z4@�f�⤏!?�9�8�(�@ugP��ٿ�'߾��@O�Z4@�f�⤏!?�9�8�(�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@-��҉�ٿ)	�3��@�G��G4@��͏!?���[�X�@'��0&�ٿ��0<��@E	|�Y 4@����Ï!?Tj�S���@'��0&�ٿ��0<��@E	|�Y 4@����Ï!?Tj�S���@'��0&�ٿ��0<��@E	|�Y 4@����Ï!?Tj�S���@'��0&�ٿ��0<��@E	|�Y 4@����Ï!?Tj�S���@'��0&�ٿ��0<��@E	|�Y 4@����Ï!?Tj�S���@t�����ٿ_·P{��@��Y- 4@�?�p��!?���69\�@�2�L�ٿ(�� �z�@�3� 4@�U7k�!?��p�t�@�2�L�ٿ(�� �z�@�3� 4@�U7k�!?��p�t�@��lh��ٿ���"���@d5#[_ 4@Xg��O�!?��9��|�@��lh��ٿ���"���@d5#[_ 4@Xg��O�!?��9��|�@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@.2 ���ٿ�K��j�@@�r�3@�0��|�!?��y����@���§ٿ�\Y��@@�4��4@�<���!?9�野��@���§ٿ�\Y��@@�4��4@�<���!?9�野��@���§ٿ�\Y��@@�4��4@�<���!?9�野��@���§ٿ�\Y��@@�4��4@�<���!?9�野��@���§ٿ�\Y��@@�4��4@�<���!?9�野��@���§ٿ�\Y��@@�4��4@�<���!?9�野��@ FT��ٿ�6|��@���s4@=�N��!?W"�>J�@ FT��ٿ�6|��@���s4@=�N��!?W"�>J�@ FT��ٿ�6|��@���s4@=�N��!?W"�>J�@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@28���ٿԷW�~�@�uМ4@��s2�!?�i.���@Q��u�ٿhFo�Q�@L����4@�q��ď!?��$5uQ�@���h�ٿ#YXS% �@㽉l4@3'�e�!?wS����@���h�ٿ#YXS% �@㽉l4@3'�e�!?wS����@���h�ٿ#YXS% �@㽉l4@3'�e�!?wS����@A��=��ٿQ�"{���@��ۂ:4@��ޏ!?����z�@A��=��ٿQ�"{���@��ۂ:4@��ޏ!?����z�@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@?���Q�ٿ7��^�,�@c��N4@~���!?i�`F��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@F��}9�ٿ��4睘�@�_��� 4@��s���!?�\� ��@y���ٿ�<���]�@Vؽ�4@�f>���!?����<n�@y���ٿ�<���]�@Vؽ�4@�f>���!?����<n�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@��k�ٿB1���@��� 4@ Z��!?H�%�z;�@�nK�d�ٿ��-_��@S�P(F4@#�ُ!?Nܸ��@Vpk�ٿ6��8~��@�'��3@�d�莏!?�������@Vpk�ٿ6��8~��@�'��3@�d�莏!?�������@Vpk�ٿ6��8~��@�'��3@�d�莏!?�������@I��'R�ٿL�8�5��@�t��4@�K��!?;6���@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@(u,P�ٿ���T���@Г�W��3@}og�V�!?�R'��=�@%k+�ٿ�+Q����@��eF 4@0	Z�!?�T�%I�@%k+�ٿ�+Q����@��eF 4@0	Z�!?�T�%I�@�����ٿ ?&���@�0�4@^�ne��!?QJ���@�����ٿ ?&���@�0�4@^�ne��!?QJ���@�����ٿ ?&���@�0�4@^�ne��!?QJ���@�����ٿ ?&���@�0�4@^�ne��!?QJ���@;^�/�ٿ�\S���@��� 4@��*L�!?�B��3^�@��Q+`�ٿ���C���@��Z�� 4@D���X�!?�{�RtC�@��Q+`�ٿ���C���@��Z�� 4@D���X�!?�{�RtC�@lj��ۨٿ������@�g�� 4@}jO�!?�-��8��@lj��ۨٿ������@�g�� 4@}jO�!?�-��8��@lj��ۨٿ������@�g�� 4@}jO�!?�-��8��@lj��ۨٿ������@�g�� 4@}jO�!?�-��8��@lj��ۨٿ������@�g�� 4@}jO�!?�-��8��@�Iv�F�ٿ(��:�+�@����3@���PA�!?�Vl�\H�@�Iv�F�ٿ(��:�+�@����3@���PA�!?�Vl�\H�@�Iv�F�ٿ(��:�+�@����3@���PA�!?�Vl�\H�@�Iv�F�ٿ(��:�+�@����3@���PA�!?�Vl�\H�@�i' �ٿ���T�@�"����3@�)uT�!?�s�7�(�@�i' �ٿ���T�@�"����3@�)uT�!?�s�7�(�@�i' �ٿ���T�@�"����3@�)uT�!?�s�7�(�@��tӛٿ�3�z��@�61�3@eIM\�!?̉7��K�@qTQm�ٿ����B�@l�-s��3@�U}B�!?���0��@�q37�ٿp+!N@��@^�� *�3@V
�!?Y߅o���@l����ٿ}�&�O�@ tD	��3@��E�!?,��r���@��GJ�ٿ�����@�/���3@�����!?j�9X��@��GJ�ٿ�����@�/���3@�����!?j�9X��@��GJ�ٿ�����@�/���3@�����!?j�9X��@��GJ�ٿ�����@�/���3@�����!?j�9X��@�'��ٿ�:�K��@��.d'�3@�V�v�!?=�����@��\�ٿ�8�����@�Mig 4@�u�N�!?�ue�a+�@" o��ٿ�i����@21�i�3@T�2�R�!?T?��p��@" o��ٿ�i����@21�i�3@T�2�R�!?T?��p��@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@��GV�ٿ�
����@gi[ 4@�,u{��!?t�m�Qq�@к����ٿI�P���@�U[H4@���8�!?eQ���@к����ٿI�P���@�U[H4@���8�!?eQ���@�U봳ٿ�ߝvq�@؎%� 4@�wz9�!?cH@����@�U봳ٿ�ߝvq�@؎%� 4@�wz9�!?cH@����@�U봳ٿ�ߝvq�@؎%� 4@�wz9�!?cH@����@=V���ٿ0+�Ԫ��@�W�d�3@38n&e�!?̜���@=V���ٿ0+�Ԫ��@�W�d�3@38n&e�!?̜���@Fjd��ٿo�L�p�@[�,� 4@r��}�!?��n���@Fjd��ٿo�L�p�@[�,� 4@r��}�!?��n���@Fjd��ٿo�L�p�@[�,� 4@r��}�!?��n���@����}�ٿv�ǭ��@�d;dO4@�@I��!?�U��7��@�Puk�ٿm߽���@DR~��4@#>��i�!?�s��k9�@�Puk�ٿm߽���@DR~��4@#>��i�!?�s��k9�@�Puk�ٿm߽���@DR~��4@#>��i�!?�s��k9�@�Puk�ٿm߽���@DR~��4@#>��i�!?�s��k9�@�ax�ٿթxc��@��ܩ�3@�a���!?���T�@�ax�ٿթxc��@��ܩ�3@�a���!?���T�@�ax�ٿթxc��@��ܩ�3@�a���!?���T�@�ax�ٿթxc��@��ܩ�3@�a���!?���T�@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@�ԙp�ٿ�����@<����3@����!?����(��@ -
m��ٿqt� �J�@ʊ���3@�o��!?C���(�@ -
m��ٿqt� �J�@ʊ���3@�o��!?C���(�@KV(��ٿ���Ib`�@�.��� 4@n_-��!?�4TF=+�@KV(��ٿ���Ib`�@�.��� 4@n_-��!?�4TF=+�@KV(��ٿ���Ib`�@�.��� 4@n_-��!?�4TF=+�@KV(��ٿ���Ib`�@�.��� 4@n_-��!?�4TF=+�@KV(��ٿ���Ib`�@�.��� 4@n_-��!?�4TF=+�@��Һ�ٿ�hq���@��@ԓ 4@:x�=��!?<o���e�@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@�����ٿ�Ԓ�@o�-~�3@�Yġ�!?��aJ��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@S�҈�ٿ9��w�@-C��3@��맏!?�x�7��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@(�)3�ٿ��b�S��@B�.��3@�d���!?�\\/��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@	ݵT�ٿr׌�Y��@�u�� 4@�E�!?lX*��@��(@�ٿ�+h���@�7�8O�3@��z���!?�$3���@��(@�ٿ�+h���@�7�8O�3@��z���!?�$3���@��(@�ٿ�+h���@�7�8O�3@��z���!?�$3���@��(@�ٿ�+h���@�7�8O�3@��z���!?�$3���@��(@�ٿ�+h���@�7�8O�3@��z���!?�$3���@�iัٿ�� ��@�_��� 4@_:���!?�V&�@�iัٿ�� ��@�_��� 4@_:���!?�V&�@�iัٿ�� ��@�_��� 4@_:���!?�V&�@�iัٿ�� ��@�_��� 4@_:���!?�V&�@�iัٿ�� ��@�_��� 4@_:���!?�V&�@�iัٿ�� ��@�_��� 4@_:���!?�V&�@!T����ٿ�rJG�@���}�3@�keky�!?,T�Ā�@!T����ٿ�rJG�@���}�3@�keky�!?,T�Ā�@!T����ٿ�rJG�@���}�3@�keky�!?,T�Ā�@!T����ٿ�rJG�@���}�3@�keky�!?,T�Ā�@!T����ٿ�rJG�@���}�3@�keky�!?,T�Ā�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��R2d�ٿ��u���@�=tSj�3@g��1t�!?���2i�@��[�ٿF%�~[�@�"�[�3@��r�1�!?F��Q�F�@��[�ٿF%�~[�@�"�[�3@��r�1�!?F��Q�F�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@�GE���ٿ�CM�E\�@dQN���3@��T4�!?Yq�E\�@O�߱��ٿ����B�@ �'� 4@�^���!?M�9\�L�@O�߱��ٿ����B�@ �'� 4@�^���!?M�9\�L�@O�߱��ٿ����B�@ �'� 4@�^���!?M�9\�L�@Lƿ?�ٿ���YE"�@&��4@�	� �!?�x����@Lƿ?�ٿ���YE"�@&��4@�	� �!?�x����@��M��ٿϊ	����@��{��4@�&)�ۏ!?H��(�!�@��M��ٿϊ	����@��{��4@�&)�ۏ!?H��(�!�@��M��ٿϊ	����@��{��4@�&)�ۏ!?H��(�!�@��M��ٿϊ	����@��{��4@�&)�ۏ!?H��(�!�@��M��ٿϊ	����@��{��4@�&)�ۏ!?H��(�!�@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@���h�ٿh��IhG�@^&4�4@NOF�ޏ!?NE#F��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@�)���ٿ:�V{�@�_p4@���Ϗ!?��0��@@�#���ٿ�Q(�i��@�Y��C 4@�D�Mj�!?奁��@�N��ٿ�
H��@qO�o4@V��@��!?�,(�'�@�N��ٿ�
H��@qO�o4@V��@��!?�,(�'�@�N��ٿ�
H��@qO�o4@V��@��!?�,(�'�@�N��ٿ�
H��@qO�o4@V��@��!?�,(�'�@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@���E�ٿ�42X��@�P����3@@c#D��!?�T)���@� "��ٿ��@l���@t7� 4@F��뗏!?��#=��@� "��ٿ��@l���@t7� 4@F��뗏!?��#=��@� "��ٿ��@l���@t7� 4@F��뗏!?��#=��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�Gy�A�ٿ��\M��@��^f4@Lwj�k�!?ᵫ� ��@�ŋ��ٿ>&ޡ���@�~�4@d�J���!?Y��X�@�ŋ��ٿ>&ޡ���@�~�4@d�J���!?Y��X�@�ŋ��ٿ>&ޡ���@�~�4@d�J���!?Y��X�@�nFH��ٿ����.g�@�x�) 4@�-�P��!?�23�]��@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@�m�?��ٿ0�:�h��@!�^�Z4@�H�qϏ!?a�=���@a����ٿ#��s��@^�""4@ӱdE��!?��:�y�@a����ٿ#��s��@^�""4@ӱdE��!?��:�y�@a����ٿ#��s��@^�""4@ӱdE��!?��:�y�@a����ٿ#��s��@^�""4@ӱdE��!?��:�y�@F�۷\�ٿ�g�sp��@��h�d 4@�7h:�!?�������@F�۷\�ٿ�g�sp��@��h�d 4@�7h:�!?�������@F�۷\�ٿ�g�sp��@��h�d 4@�7h:�!?�������@F�۷\�ٿ�g�sp��@��h�d 4@�7h:�!?�������@F�۷\�ٿ�g�sp��@��h�d 4@�7h:�!?�������@�����ٿɖ/�I�@{󚼠�3@n�s��!?)��=�@�����ٿɖ/�I�@{󚼠�3@n�s��!?)��=�@����צٿ>��jI[�@�ϣ��3@���j�!?�,fs��@~��ٿ�VUL���@���N��3@��㛺�!?ar8�|�@~��ٿ�VUL���@���N��3@��㛺�!?ar8�|�@~��ٿ�VUL���@���N��3@��㛺�!?ar8�|�@~��ٿ�VUL���@���N��3@��㛺�!?ar8�|�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@(���7�ٿ�qE��@��OgL�3@�cų��!?�	i�B�@39�u�ٿ�!���x�@8(2=�4@d?.���!?t1����@39�u�ٿ�!���x�@8(2=�4@d?.���!?t1����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@��dFЪٿdR�Su�@����� 4@��ĥ�!?aC����@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@x���ٿp�ψ��@���	�4@(M����!?w\�d\,�@�68#�ٿ�'zx��@�;m�4@����ŏ!?w�xW�-�@�68#�ٿ�'zx��@�;m�4@����ŏ!?w�xW�-�@ДaW֡ٿ\�,a���@U���4@����ݏ!?P{-���@ДaW֡ٿ\�,a���@U���4@����ݏ!?P{-���@ДaW֡ٿ\�,a���@U���4@����ݏ!?P{-���@ДaW֡ٿ\�,a���@U���4@����ݏ!?P{-���@�K�ިٿ�&;:�O�@=���4@2�ԕ�!?Tt�W"T�@�K�ިٿ�&;:�O�@=���4@2�ԕ�!?Tt�W"T�@�K�ިٿ�&;:�O�@=���4@2�ԕ�!?Tt�W"T�@�K�ިٿ�&;:�O�@=���4@2�ԕ�!?Tt�W"T�@�K�ިٿ�&;:�O�@=���4@2�ԕ�!?Tt�W"T�@��1�ٿD^K牃�@+�Ch4@m˫&��!?`j�iJ��@��1�ٿD^K牃�@+�Ch4@m˫&��!?`j�iJ��@��1�ٿD^K牃�@+�Ch4@m˫&��!?`j�iJ��@��1�ٿD^K牃�@+�Ch4@m˫&��!?`j�iJ��@��1�ٿD^K牃�@+�Ch4@m˫&��!?`j�iJ��@��S���ٿ��+�E��@/��y��3@�S�K�!?��$x�'�@˭E
E�ٿ��gf� �@X��!P�3@�D7rŏ!?�X�H���@˭E
E�ٿ��gf� �@X��!P�3@�D7rŏ!?�X�H���@˭E
E�ٿ��gf� �@X��!P�3@�D7rŏ!?�X�H���@��l���ٿ2	Vt�r�@-Hi� 4@;���ŏ!?��BY�y�@��l���ٿ2	Vt�r�@-Hi� 4@;���ŏ!?��BY�y�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@
���]�ٿ��A���@�HbO�4@�	����!?��ŠG�@y�0��ٿs�%��z�@x�gH�4@3��	��!?� �����@y�0��ٿs�%��z�@x�gH�4@3��	��!?� �����@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�A����ٿ��.���@��Y� 4@įݳ�!?T��~��@�����ٿ��ﱢ�@�{ҝ 4@(7p�ԏ!?[=���&�@�����ٿ��ﱢ�@�{ҝ 4@(7p�ԏ!?[=���&�@;{^lW�ٿ�z���Z�@ȼ-}��3@��'׏!?�O��QR�@D�Mn2�ٿ��g��t�@Ō�Y��3@k��؏!?�l;���@U7���ٿ��A#�^�@�f�c�3@�c-�`�!??�8��s�@U7���ٿ��A#�^�@�f�c�3@�c-�`�!??�8��s�@��e���ٿ��ɭ���@��ܫ4@-�1Vm�!?�f�9�@��e���ٿ��ɭ���@��ܫ4@-�1Vm�!?�f�9�@m�y�Z�ٿ3��ϧ}�@'Vjv4@p�G�Y�!?�ߐ���@m�y�Z�ٿ3��ϧ}�@'Vjv4@p�G�Y�!?�ߐ���@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@��J���ٿ�-˥P��@ύ�3�4@M)܋��!?sp^Ky�@x�^��ٿ�ɵW��@�S�,J4@Gde��!?TeHk��@x�^��ٿ�ɵW��@�S�,J4@Gde��!?TeHk��@x�^��ٿ�ɵW��@�S�,J4@Gde��!?TeHk��@�Ⱥn�ٿ�-ҽw�@�.'y��3@eT����!?�W�"�@�Ⱥn�ٿ�-ҽw�@�.'y��3@eT����!?�W�"�@�Ⱥn�ٿ�-ҽw�@�.'y��3@eT����!?�W�"�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@�����ٿ�tf�P��@���� 4@'2�Z��!?��)s�@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@"�Y���ٿP:�I׋�@O��-� 4@������!?��ct��@ǿ^���ٿ�NK ��@<�C�Z4@,�w(r�!?G�����@ǿ^���ٿ�NK ��@<�C�Z4@,�w(r�!?G�����@�퇏�ٿ���L\��@�qV�4@7s��t�!?�9{g�@{oU�*�ٿ���	�@��hk4@�"+��!?�3n���@��ֶ&�ٿ��@Ow�H4@I�at�!?�wGQ���@��ֶ&�ٿ��@Ow�H4@I�at�!?�wGQ���@��ֶ&�ٿ��@Ow�H4@I�at�!?�wGQ���@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@�X� ԧٿ��v����@��l�4@
�#���!?�e��3�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@>OX��ٿH5�c|��@M�4� 4@���V��!?�-b�J�@�"3�S�ٿ�G��c�@����g�3@U%u��!?��o1�(�@���b�ٿ�� ���@7�E��3@z��{�!?&ƴcym�@6��qg�ٿ�gECb�@��D���3@0�󚝏!?Iʂu��@6��qg�ٿ�gECb�@��D���3@0�󚝏!?Iʂu��@)/J�ٿ��Ҿ��@m���M�3@]Ech�!?n֛����@)/J�ٿ��Ҿ��@m���M�3@]Ech�!?n֛����@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@6N�Ěٿ�bՐ�@�v,90�3@g[|��!?��LIm��@�]����ٿc�����@ ��A�3@oM��`�!?/E
�a��@�]����ٿc�����@ ��A�3@oM��`�!?/E
�a��@�]����ٿc�����@ ��A�3@oM��`�!?/E
�a��@�]����ٿc�����@ ��A�3@oM��`�!?/E
�a��@GiVã�ٿ����s�@��.5��3@��M]��!?a�����@GiVã�ٿ����s�@��.5��3@��M]��!?a�����@ �९�ٿ*�|��@< � 4@���Ե�!?=�n�qp�@ �९�ٿ*�|��@< � 4@���Ե�!?=�n�qp�@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@��N��ٿ旦��w�@�*u�[4@
�ߞ��!?��#��@�$�*�ٿs��Q�@\�UJ� 4@��'ʏ!?&j��e��@"!rj,�ٿ�ռxE%�@�2ʔ� 4@�k-���!?Sk����@"!rj,�ٿ�ռxE%�@�2ʔ� 4@�k-���!?Sk����@�H�0ޜٿ�l�d�@�H��Y4@M��Q��!?��_�:��@�H�0ޜٿ�l�d�@�H��Y4@M��Q��!?��_�:��@�H�0ޜٿ�l�d�@�H��Y4@M��Q��!?��_�:��@�H�0ޜٿ�l�d�@�H��Y4@M��Q��!?��_�:��@�H�0ޜٿ�l�d�@�H��Y4@M��Q��!?��_�:��@�.F��ٿ�$$]��@���;a4@�g��!?W�-9��@�5P�ٿTlTc��@��C; 4@� 7��!?ew�u���@�5P�ٿTlTc��@��C; 4@� 7��!?ew�u���@�5P�ٿTlTc��@��C; 4@� 7��!?ew�u���@�5P�ٿTlTc��@��C; 4@� 7��!?ew�u���@�r���ٿ}�kB�@O��)4@�H����!?��<����@�r���ٿ}�kB�@O��)4@�H����!?��<����@�r���ٿ}�kB�@O��)4@�H����!?��<����@�r���ٿ}�kB�@O��)4@�H����!?��<����@�r���ٿ}�kB�@O��)4@�H����!?��<����@�r���ٿ}�kB�@O��)4@�H����!?��<����@sd�?�ٿ���t�o�@��u��4@>0���!?|B�蛭�@sd�?�ٿ���t�o�@��u��4@>0���!?|B�蛭�@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@��9��ٿ�X�"��@�1�BS 4@k�bُ!?��/���@(��`r�ٿ�R5���@���4@<�����!?���X%��@(��`r�ٿ�R5���@���4@<�����!?���X%��@r�JƠٿR����@��v� 4@.�WK�!?��,���@U�s�ٿ�Ǫ���@\?�t 4@�w^E�!?������@U�s�ٿ�Ǫ���@\?�t 4@�w^E�!?������@U�s�ٿ�Ǫ���@\?�t 4@�w^E�!?������@U�s�ٿ�Ǫ���@\?�t 4@�w^E�!?������@U�s�ٿ�Ǫ���@\?�t 4@�w^E�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@mm�h�ٿ�b�K��@:cw�} 4@�CZ�i�!?������@m"���ٿd�T0�Z�@�/1� 4@a ��o�!?������@m"���ٿd�T0�Z�@�/1� 4@a ��o�!?������@m"���ٿd�T0�Z�@�/1� 4@a ��o�!?������@m"���ٿd�T0�Z�@�/1� 4@a ��o�!?������@m"���ٿd�T0�Z�@�/1� 4@a ��o�!?������@���e�ٿ����x�@��� 4@* Dr�!?�s�#�@���e�ٿ����x�@��� 4@* Dr�!?�s�#�@���e�ٿ����x�@��� 4@* Dr�!?�s�#�@�+�ٿCQ_P��@�U� 4@9��nY�!?�X�2���@�+�ٿCQ_P��@�U� 4@9��nY�!?�X�2���@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@�,��D�ٿ�W�o��@m�	׷ 4@�E��u�!?v/t��@7[5�ٿ�Vҿ�U�@��o6n 4@�:��V�!?�@Pw,�@7[5�ٿ�Vҿ�U�@��o6n 4@�:��V�!?�@Pw,�@7[5�ٿ�Vҿ�U�@��o6n 4@�:��V�!?�@Pw,�@7[5�ٿ�Vҿ�U�@��o6n 4@�:��V�!?�@Pw,�@7[5�ٿ�Vҿ�U�@��o6n 4@�:��V�!?�@Pw,�@b#j�*�ٿ�۽��>�@3���  4@!���T�!?�lZ�GP�@b#j�*�ٿ�۽��>�@3���  4@!���T�!?�lZ�GP�@b#j�*�ٿ�۽��>�@3���  4@!���T�!?�lZ�GP�@�Aw�h�ٿkz�f� �@N���3@:�˃x�!?�d�Z�@�Aw�h�ٿkz�f� �@N���3@:�˃x�!?�d�Z�@����ٿ��6�4�@�.OO��3@��siT�!?�q�)�~�@�jeP
�ٿl[�K�l�@0�S?��3@a���(�!?v9��)��@S�Uܬٿ�f��Ȏ�@v�k���3@L�\z�!?�y�>I(�@S�Uܬٿ�f��Ȏ�@v�k���3@L�\z�!?�y�>I(�@S�Uܬٿ�f��Ȏ�@v�k���3@L�\z�!?�y�>I(�@S�Uܬٿ�f��Ȏ�@v�k���3@L�\z�!?�y�>I(�@���QH�ٿ3��n�M�@PC�4@�+X�2�!?p:%�c9�@���QH�ٿ3��n�M�@PC�4@�+X�2�!?p:%�c9�@_����ٿ����W�@��C�4@����"�!?���65��@_����ٿ����W�@��C�4@����"�!?���65��@_����ٿ����W�@��C�4@����"�!?���65��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�G\,t�ٿ��
���@���h44@]��༏!?���ݸ��@�1ͳ��ٿ��Uq�@U7)�4@XB�o�!?��w���@�1ͳ��ٿ��Uq�@U7)�4@XB�o�!?��w���@�1ͳ��ٿ��Uq�@U7)�4@XB�o�!?��w���@�1ͳ��ٿ��Uq�@U7)�4@XB�o�!?��w���@�1ͳ��ٿ��Uq�@U7)�4@XB�o�!?��w���@_QFo�ٿ]{���*�@	#o��4@w6�ߞ�!?:��JIo�@_QFo�ٿ]{���*�@	#o��4@w6�ߞ�!?:��JIo�@n��v��ٿ��,�k�@�{+��4@������!?�-T�o��@n��v��ٿ��,�k�@�{+��4@������!?�-T�o��@n��v��ٿ��,�k�@�{+��4@������!?�-T�o��@n��v��ٿ��,�k�@�{+��4@������!?�-T�o��@n��v��ٿ��,�k�@�{+��4@������!?�-T�o��@�];��ٿٚ��L�@t�4@5psď!?�R�B�@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�N�h��ٿ�
���@f3�{z�3@=�tЏ!?݉2��@�o�٪�ٿY;����@�؃O�4@ė�!?������@�o�٪�ٿY;����@�؃O�4@ė�!?������@�o�٪�ٿY;����@�؃O�4@ė�!?������@�o�٪�ٿY;����@�؃O�4@ė�!?������@�o�٪�ٿY;����@�؃O�4@ė�!?������@�o�٪�ٿY;����@�؃O�4@ė�!?������@	P�-(�ٿG�i ��@o#Eǣ 4@���t��!?��Tkt�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@߫���ٿ��9_@�@�=�3�4@�|��"�!?j@��V�@�A���ٿrV��E�@M�F� 4@���Ï!?p�:���@�A���ٿrV��E�@M�F� 4@���Ï!?p�:���@f�'?a�ٿ����8C�@�G�m4@�-��ۏ!?���vL��@f�'?a�ٿ����8C�@�G�m4@�-��ۏ!?���vL��@f�'?a�ٿ����8C�@�G�m4@�-��ۏ!?���vL��@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@�ֱ�b�ٿ׌j ���@��jL�4@>��;��!?�v�r���@��pE!�ٿG6$����@*�U��4@ ��bҏ!?Z��k&&�@��pE!�ٿG6$����@*�U��4@ ��bҏ!?Z��k&&�@��pE!�ٿG6$����@*�U��4@ ��bҏ!?Z��k&&�@��pE!�ٿG6$����@*�U��4@ ��bҏ!?Z��k&&�@��pE!�ٿG6$����@*�U��4@ ��bҏ!?Z��k&&�@HR�s��ٿ�������@�u4@��:�Ǐ!?z9�g��@#���ٿ��m���@���/�4@K{VM��!?�'��G��@#���ٿ��m���@���/�4@K{VM��!?�'��G��@#���ٿ��m���@���/�4@K{VM��!?�'��G��@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��4�:�ٿ��\��@�R�+4@:!}Ș�!?7��H�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@��z�ٿCl|�@�RG�4@Wd��!?u�N��a�@������ٿſ�H�@/١4@���ji�!?�@js��@������ٿſ�H�@/١4@���ji�!?�@js��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@s[t�ٿ`k���@yB�I� 4@ؔ�d3�!?�,�E1��@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@�c
}��ٿ,7��_��@8IO� 4@��'U�!?D���,A�@d&H�ٿ)���u�@����]�3@jI�r�!?�\����@d&H�ٿ)���u�@����]�3@jI�r�!?�\����@ =��B�ٿ(v�9#�@��(��3@$��ʏ!?�P&�N�@ =��B�ٿ(v�9#�@��(��3@$��ʏ!?�P&�N�@��C<�ٿG���c��@�Gպ��3@Q�sL��!?��Oo-��@��C<�ٿG���c��@�Gպ��3@Q�sL��!?��Oo-��@��C<�ٿG���c��@�Gպ��3@Q�sL��!?��Oo-��@vv{g�ٿ��w;*I�@O~+j��3@��S�ŏ!?�,(ED��@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@��F(�ٿ?��@u��@��J̳4@>��֏!?�Z����@`��^=�ٿ�h�0X�@�ͼ24@��b��!?h(�/6�@`��^=�ٿ�h�0X�@�ͼ24@��b��!?h(�/6�@`��^=�ٿ�h�0X�@�ͼ24@��b��!?h(�/6�@`��^=�ٿ�h�0X�@�ͼ24@��b��!?h(�/6�@�R%��ٿ�'�E��@�c��`4@�����!?��Q��@�R%��ٿ�'�E��@�c��`4@�����!?��Q��@�R%��ٿ�'�E��@�c��`4@�����!?��Q��@�R%��ٿ�'�E��@�c��`4@�����!?��Q��@m�!`��ٿP�9j��@=n���4@����!?�D����@m�!`��ٿP�9j��@=n���4@����!?�D����@m�!`��ٿP�9j��@=n���4@����!?�D����@m�!`��ٿP�9j��@=n���4@����!?�D����@m�!`��ٿP�9j��@=n���4@����!?�D����@|mH�,�ٿ�İ��@b�V���3@���z�!?S�e( ��@|mH�,�ٿ�İ��@b�V���3@���z�!?S�e( ��@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@�����ٿ��?��@Ji�.�4@�Q�*o�!?(�iK���@��W\�ٿ�*e(��@Y��}�4@4�ҫ��!?f�"���@��W\�ٿ�*e(��@Y��}�4@4�ҫ��!?f�"���@��W\�ٿ�*e(��@Y��}�4@4�ҫ��!?f�"���@��W\�ٿ�*e(��@Y��}�4@4�ҫ��!?f�"���@��W\�ٿ�*e(��@Y��}�4@4�ҫ��!?f�"���@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@�W�Ԙٿ`tg���@:��4@�	x��!?UR�8R��@#d���ٿ���tk�@x(y 4@�WT ��!?����j*�@#d���ٿ���tk�@x(y 4@�WT ��!?����j*�@#d���ٿ���tk�@x(y 4@�WT ��!?����j*�@8�胟ٿ��MN&�@�[Y4@I��N#�!?�}bY��@8�胟ٿ��MN&�@�[Y4@I��N#�!?�}bY��@8�胟ٿ��MN&�@�[Y4@I��N#�!?�}bY��@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@hr:��ٿU8h	��@n*�� 4@�cw�!?H�|�7]�@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@�j�(��ٿ�K�C���@�1��" 4@�~_�i�!?c�b3f��@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@*�v�ԟٿM��)��@��}�4@M,I�!?�:����@�|~^�ٿ阝l|g�@įmР�3@x��p-�!?�"b��@�|~^�ٿ阝l|g�@įmР�3@x��p-�!?�"b��@�|~^�ٿ阝l|g�@įmР�3@x��p-�!?�"b��@�|~^�ٿ阝l|g�@įmР�3@x��p-�!?�"b��@�|~^�ٿ阝l|g�@įmР�3@x��p-�!?�"b��@^ء-�ٿ�EDI--�@�J?�4@1s!��!?~�W����@^ء-�ٿ�EDI--�@�J?�4@1s!��!?~�W����@�ET;#�ٿ���f�@�ak�� 4@���-Џ!?�� ��@�ET;#�ٿ���f�@�ak�� 4@���-Џ!?�� ��@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@���՛ٿ�ou����@�G�
4@�^[o�!?͐Ǐ�!�@F{��z�ٿeVEkM�@h�:Z� 4@v�+n*�!?�)qZ��@F{��z�ٿeVEkM�@h�:Z� 4@v�+n*�!?�)qZ��@F{��z�ٿeVEkM�@h�:Z� 4@v�+n*�!?�)qZ��@����ٿ
���f�@tq
4@�A\�q�!?�����@����ٿ
���f�@tq
4@�A\�q�!?�����@����ٿ
���f�@tq
4@�A\�q�!?�����@�	A�ٿp%h�2.�@6�M�4@��g��!?1�]`� �@�	A�ٿp%h�2.�@6�M�4@��g��!?1�]`� �@�	A�ٿp%h�2.�@6�M�4@��g��!?1�]`� �@�	A�ٿp%h�2.�@6�M�4@��g��!?1�]`� �@�	A�ٿp%h�2.�@6�M�4@��g��!?1�]`� �@�����ٿ��\����@�eҍ� 4@�2�R�!?��J�t�@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@��<�z�ٿ�����@XA�g�4@�jeΏ!??���p��@�/wu�ٿ�J�a`^�@)�TM4@�%E��!?��/�@���Y�ٿ:rs��/�@
f�n 4@z�Ҟ�!?��lO�@���Y�ٿ:rs��/�@
f�n 4@z�Ҟ�!?��lO�@���Y�ٿ:rs��/�@
f�n 4@z�Ҟ�!?��lO�@�Pg4C�ٿ������@�lb�d 4@�ex2��!?֙�P���@�Pg4C�ٿ������@�lb�d 4@�ex2��!?֙�P���@�Pg4C�ٿ������@�lb�d 4@�ex2��!?֙�P���@�zy�o�ٿo�����@���r6 4@Pr�j��!??�0�%y�@�zy�o�ٿo�����@���r6 4@Pr�j��!??�0�%y�@�zy�o�ٿo�����@���r6 4@Pr�j��!??�0�%y�@�zy�o�ٿo�����@���r6 4@Pr�j��!??�0�%y�@�zy�o�ٿo�����@���r6 4@Pr�j��!??�0�%y�@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�_5.�ٿ0L�A��@�U!� 4@ˬ�!?Cr~����@�e�b�ٿ6��M_�@y:�#��3@���q�!?)be�F�@�e�b�ٿ6��M_�@y:�#��3@���q�!?)be�F�@�e�b�ٿ6��M_�@y:�#��3@���q�!?)be�F�@"V%��ٿ��*E\�@�����3@1ޗ5i�!?Yy�	��@"V%��ٿ��*E\�@�����3@1ޗ5i�!?Yy�	��@"V%��ٿ��*E\�@�����3@1ޗ5i�!?Yy�	��@"V%��ٿ��*E\�@�����3@1ޗ5i�!?Yy�	��@"V%��ٿ��*E\�@�����3@1ޗ5i�!?Yy�	��@W�Z��ٿr������@��*�4@*̔�|�!?���5xS�@W�Z��ٿr������@��*�4@*̔�|�!?���5xS�@W�Z��ٿr������@��*�4@*̔�|�!?���5xS�@W�Z��ٿr������@��*�4@*̔�|�!?���5xS�@w+�
�ٿ�G����@��"T 4@��<�W�!?i�5��@�@w+�
�ٿ�G����@��"T 4@��<�W�!?i�5��@�@d\/P٥ٿ_V��]@�@T[|��3@��ǽ�!?�s���@��R}%�ٿ��Rӑ�@i��wI 4@:w�	؏!?��µ���@��R}%�ٿ��Rӑ�@i��wI 4@:w�	؏!?��µ���@��R}%�ٿ��Rӑ�@i��wI 4@:w�	؏!?��µ���@��R}%�ٿ��Rӑ�@i��wI 4@:w�	؏!?��µ���@��V�T�ٿz�*)�r�@��,���3@��ď!?J2w���@��V�T�ٿz�*)�r�@��,���3@��ď!?J2w���@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@v��Ǧٿ�X����@=e�o� 4@���!?�k�:t�@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@9��M�ٿԵ�����@��q�4�3@ԂY��!?�����@��,�#�ٿ6O$�t�@�T?���3@&�F��!?7� ~B�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@~�2.�ٿ�M����@����3@&E|ď!?ø$�P%�@/��@�ٿ�.�Q���@lԔF�4@���!?4'�IU�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@^��;ӣٿ��>ba+�@�'�74@��)��!?��fk�@�@!џٿ�dŹ��@��=Dp 4@�N4|�!?6�JCe�@!џٿ�dŹ��@��=Dp 4@�N4|�!?6�JCe�@!џٿ�dŹ��@��=Dp 4@�N4|�!?6�JCe�@�4�z�ٿ������@��I�� 4@�	���!?�&54��@�4�z�ٿ������@��I�� 4@�	���!?�&54��@�4�z�ٿ������@��I�� 4@�	���!?�&54��@�4�z�ٿ������@��I�� 4@�	���!?�&54��@�4�z�ٿ������@��I�� 4@�	���!?�&54��@[�VP�ٿ���!��@µ�%l4@�[H��!?!l���@[�VP�ٿ���!��@µ�%l4@�[H��!?!l���@[�VP�ٿ���!��@µ�%l4@�[H��!?!l���@d�
��ٿ������@[z�ʞ 4@�?QJ�!?*��_�@�A];n�ٿr���O�@m��/��3@B׳\��!?<����@�����ٿ��
�F�@PH�+��3@��!?ᵟo�&�@�۾.,�ٿq}�x�(�@PQ�L�4@�B���!?�r�^C��@�#��
�ٿ2'̑�@�Q<4@]��!?G_M�m��@�#��
�ٿ2'̑�@�Q<4@]��!?G_M�m��@�#��
�ٿ2'̑�@�Q<4@]��!?G_M�m��@�#��
�ٿ2'̑�@�Q<4@]��!?G_M�m��@�#��
�ٿ2'̑�@�Q<4@]��!?G_M�m��@β�6�ٿ�ې|� �@�ţb*4@�uB��!?�fHNz�@β�6�ٿ�ې|� �@�ţb*4@�uB��!?�fHNz�@β�6�ٿ�ې|� �@�ţb*4@�uB��!?�fHNz�@β�6�ٿ�ې|� �@�ţb*4@�uB��!?�fHNz�@β�6�ٿ�ې|� �@�ţb*4@�uB��!?�fHNz�@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@��Y�ٿߛ��#Y�@Z��+ �3@��Ɖ�!?��Е��@ݭ���ٿ�� +�T�@Ј;���3@�^���!?*�e���@ݭ���ٿ�� +�T�@Ј;���3@�^���!?*�e���@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@r���a�ٿh�ؠS�@���p��3@��i��!?��I��@2Lk��ٿ��&�@�I� 4@��5���!?9���Q��@2Lk��ٿ��&�@�I� 4@��5���!?9���Q��@2Lk��ٿ��&�@�I� 4@��5���!?9���Q��@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@%���ٿ�����q�@�f��K4@Y�����!?q'���`�@R�h��ٿ`�l�
��@/D�� 4@4B���!?�-~�@R�h��ٿ`�l�
��@/D�� 4@4B���!?�-~�@R�h��ٿ`�l�
��@/D�� 4@4B���!?�-~�@���p��ٿ�fv(���@ �� � 4@��q�l�!?��AW@b�@���p��ٿ�fv(���@ �� � 4@��q�l�!?��AW@b�@���p��ٿ�fv(���@ �� � 4@��q�l�!?��AW@b�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@���§ٿ#!w����@�FP�h�3@�D۳��!?W���,�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@��*'��ٿ}Zក��@A@B��4@�C���!?�����q�@d�L�-�ٿ������@gz�%4@(�Pߏ!?w����@d�L�-�ٿ������@gz�%4@(�Pߏ!?w����@���ٿ�jN{R�@��i�R4@	b��t�!?�Y�K���@���ٿ�jN{R�@��i�R4@	b��t�!?�Y�K���@���ٿ�jN{R�@��i�R4@	b��t�!?�Y�K���@��\u��ٿ1��
�@����4@S�Ѯ�!?�������@��\u��ٿ1��
�@����4@S�Ѯ�!?�������@��\u��ٿ1��
�@����4@S�Ѯ�!?�������@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@��N�9�ٿҍ����@��+4Y4@���؏!?W����w�@�]����ٿ3�4%�g�@�0��>�3@�j���!? ���i��@�.�?�ٿ����$l�@��s��3@��S�!?���b�@�.�?�ٿ����$l�@��s��3@��S�!?���b�@�.�?�ٿ����$l�@��s��3@��S�!?���b�@�.�?�ٿ����$l�@��s��3@��S�!?���b�@�P�Z�ٿ89ʙ�H�@`�2��3@�\���!??�8Na�@�P�Z�ٿ89ʙ�H�@`�2��3@�\���!??�8Na�@�P�Z�ٿ89ʙ�H�@`�2��3@�\���!??�8Na�@�P�Z�ٿ89ʙ�H�@`�2��3@�\���!??�8Na�@����^�ٿ���=�m�@�	'�Z4@P2�붏!?���,cQ�@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@�U��+�ٿl��{��@D`@�} 4@54i��!?��w��@BK�Y��ٿ7�)�Ě�@Sa�2q4@R�ͨ��!?
6
3��@BK�Y��ٿ7�)�Ě�@Sa�2q4@R�ͨ��!?
6
3��@BK�Y��ٿ7�)�Ě�@Sa�2q4@R�ͨ��!?
6
3��@BK�Y��ٿ7�)�Ě�@Sa�2q4@R�ͨ��!?
6
3��@BK�Y��ٿ7�)�Ě�@Sa�2q4@R�ͨ��!?
6
3��@z��.�ٿ��ĭ�@;�i��4@vH���!?��v��@�n~p�ٿ�}O�`�@:�kX4@?Z���!?nsJ
�u�@�n~p�ٿ�}O�`�@:�kX4@?Z���!?nsJ
�u�@�n~p�ٿ�}O�`�@:�kX4@?Z���!?nsJ
�u�@�n~p�ٿ�}O�`�@:�kX4@?Z���!?nsJ
�u�@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@~���ٿ�&~Sq��@���� 4@��ڏ!?�ǪO��@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@1}��8�ٿޔX�4�@������3@�J��!?ow���y�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@�3�u$�ٿV t���@�AM� 4@g�`�!?��	5�,�@x4�.p�ٿ�HA�®�@1��؀4@��u9�!?���}��@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@��@�!�ٿ,��I��@�cd�(4@��>O�!?yd����@N�*�I�ٿ>V��3�@<]�� 4@~*yN��!?4x0pG�@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@�'S�V�ٿ�}���W�@�t�T��3@P��/��!?Y���@��@s���ٿ���1��@S�2j��3@��/ݏ!?�s���D�@s���ٿ���1��@S�2j��3@��/ݏ!?�s���D�@s���ٿ���1��@S�2j��3@��/ݏ!?�s���D�@s���ٿ���1��@S�2j��3@��/ݏ!?�s���D�@�v�2R�ٿ���'#z�@+g�0��3@��U��!?y��n�\�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@����d�ٿ�cC#�}�@�X�[ 4@�k	il�!?�s�K4�@8c�ٿy� M�>�@�Df���3@}?i���!?'P�J��@8c�ٿy� M�>�@�Df���3@}?i���!?'P�J��@8c�ٿy� M�>�@�Df���3@}?i���!?'P�J��@8c�ٿy� M�>�@�Df���3@}?i���!?'P�J��@8c�ٿy� M�>�@�Df���3@}?i���!?'P�J��@Ø�ʩٿW#m��@�Aw� 4@�.���!?s/h�ɼ�@Ø�ʩٿW#m��@�Aw� 4@�.���!?s/h�ɼ�@Ø�ʩٿW#m��@�Aw� 4@�.���!?s/h�ɼ�@Ø�ʩٿW#m��@�Aw� 4@�.���!?s/h�ɼ�@Ø�ʩٿW#m��@�Aw� 4@�.���!?s/h�ɼ�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@�6퀹�ٿw�l��@J�T 4@K����!?�O �s�@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@}#��ٿ��N
n�@"��o 4@�c�%%�!?k{�m��@�pT�`�ٿ��I/�x�@H�	�Q�3@@t��!?��٪O<�@�pT�`�ٿ��I/�x�@H�	�Q�3@@t��!?��٪O<�@�pT�`�ٿ��I/�x�@H�	�Q�3@@t��!?��٪O<�@�pT�`�ٿ��I/�x�@H�	�Q�3@@t��!?��٪O<�@W��b6�ٿ�r'�\o�@�կ ��3@�����!?��R�A"�@W��b6�ٿ�r'�\o�@�կ ��3@�����!?��R�A"�@o8�|�ٿ�V��~�@��Cz-�3@�Mҏ!?��ɠ�r�@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@����ٿ��rL��@�4�| 4@�X2��!?�++���@�g����ٿ��o}��@���S�4@�X�s�!?�˜7�@�g����ٿ��o}��@���S�4@�X�s�!?�˜7�@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@̬��ٿ�QoE��@��߯J 4@�Bo�!?)�[#j��@�1xߓٿ�g�}���@��4@om7M�!?�����&�@�1xߓٿ�g�}���@��4@om7M�!?�����&�@��i�ٿ�a�B���@7�([4@�l��!?��f=�y�@��i�ٿ�a�B���@7�([4@�l��!?��f=�y�@��i�ٿ�a�B���@7�([4@�l��!?��f=�y�@��i�ٿ�a�B���@7�([4@�l��!?��f=�y�@��i�ٿ�a�B���@7�([4@�l��!?��f=�y�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@srA�՟ٿ�3��V�@K�`� 4@r�^�s�!?+_�^�@�7͓��ٿ�c|?r�@�ňMN4@ƍI���!?E�,�@�7͓��ٿ�c|?r�@�ňMN4@ƍI���!?E�,�@�7͓��ٿ�c|?r�@�ňMN4@ƍI���!?E�,�@�7͓��ٿ�c|?r�@�ňMN4@ƍI���!?E�,�@�7͓��ٿ�c|?r�@�ňMN4@ƍI���!?E�,�@vJ>��ٿ�U� ���@e`�4@V��$6�!?��q�Me�@vJ>��ٿ�U� ���@e`�4@V��$6�!?��q�Me�@7�ε��ٿ���{�|�@!D���4@]�DIя!?!��^n��@7�ε��ٿ���{�|�@!D���4@]�DIя!?!��^n��@_��o�ٿ�%̢�l�@�R�� 4@>��ᯏ!?�1�����@y���ˮٿ��H+��@�ּ4@ƈ�!?�ɝ��P�@y���ˮٿ��H+��@�ּ4@ƈ�!?�ɝ��P�@�dp7�ٿDj4����@�gTo4@����ߏ!?���`A�@u(�� �ٿ�����@�ӕ�4@Lz��!?�Bkj\�@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@�9$MU�ٿ��b%���@�1LMu4@�Tz�!?S�1�r��@����
�ٿ^Z@����@�8���4@�W��@�!?�C8#�O�@�Em̙ٿ���?�@��%1��3@����͏!?�o@�?�@[����ٿ�1�<9�@����R�3@�B�ȏ!?@_�;2)�@��*8�ٿ_���}�@���n��3@;%$���!? _ԋ�@El"W'�ٿl)�1n�@�J�Y�3@������!?��J��B�@&ĺߊ�ٿ�I�$�Y�@�V��M 4@x<ה��!?����@���؟ٿ�:��k�@���N� 4@�&����!?�5K��@���؟ٿ�:��k�@���N� 4@�&����!?�5K��@���ٿ��dH�@A��� 4@hj:g�!?DB�m�v�@��EcG�ٿ�Vb�@~�Ţ 4@�3y�!?С�E-�@��EcG�ٿ�Vb�@~�Ţ 4@�3y�!?С�E-�@��EcG�ٿ�Vb�@~�Ţ 4@�3y�!?С�E-�@��EcG�ٿ�Vb�@~�Ţ 4@�3y�!?С�E-�@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@�yZy��ٿ�No-}�@_3F8 4@��m�z�!?t�e���@ξ�[�ٿ؈+Y��@�5<6 4@�;��ۏ!?K�����@ξ�[�ٿ؈+Y��@�5<6 4@�;��ۏ!?K�����@ξ�[�ٿ؈+Y��@�5<6 4@�;��ۏ!?K�����@ξ�[�ٿ؈+Y��@�5<6 4@�;��ۏ!?K�����@ξ�[�ٿ؈+Y��@�5<6 4@�;��ۏ!?K�����@�
?���ٿ-���c�@C�I 4@�JE��!?ߔ[�)��@�
?���ٿ-���c�@C�I 4@�JE��!?ߔ[�)��@�
?���ٿ-���c�@C�I 4@�JE��!?ߔ[�)��@�
?���ٿ-���c�@C�I 4@�JE��!?ߔ[�)��@�J� ��ٿ���a��@��4@�e�X��!? �8mf�@�J� ��ٿ���a��@��4@�e�X��!? �8mf�@�jJ6�ٿ�@p�!��@Hb� 4@�[qۏ!?d=�@�@�F��ٿFVy�3��@��_�� 4@	娏��!?|�у��@�@�F��ٿFVy�3��@��_�� 4@	娏��!?|�у��@�@�F��ٿFVy�3��@��_�� 4@	娏��!?|�у��@�@�F��ٿFVy�3��@��_�� 4@	娏��!?|�у��@�����ٿ^�)Y��@�����4@��|G��!?ၓ>4��@�����ٿ^�)Y��@�����4@��|G��!?ၓ>4��@jKl4�ٿ�_'���@��.�Q�3@
)��!?2�Ą���@jKl4�ٿ�_'���@��.�Q�3@
)��!?2�Ą���@jKl4�ٿ�_'���@��.�Q�3@
)��!?2�Ą���@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@���ӧٿ�-w��@�v[��3@x�MMҏ!?H*����@�׫r�ٿe����@���(4@�;#4��!?��?ȅn�@����ٿ\�����@ �.I4@�O^���!?�Ȫ�Ӝ�@Z���ٿ����@�Iu�4@�7���!?�{w�so�@A�])b�ٿ��]�M�@�?���4@7
��G�!?�� !
��@A�])b�ٿ��]�M�@�?���4@7
��G�!?�� !
��@A�])b�ٿ��]�M�@�?���4@7
��G�!?�� !
��@�^�s�ٿ5�,l��@O#�4@�G�V�!?`I9׉��@�^�s�ٿ5�,l��@O#�4@�G�V�!?`I9׉��@h�X�ٿ1��<��@J>�I}4@����!?�4o�[�@h�X�ٿ1��<��@J>�I}4@����!?�4o�[�@h�X�ٿ1��<��@J>�I}4@����!?�4o�[�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@�b�zR�ٿ����e��@�J��4@�ُG��!?��A�@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@��$���ٿ������@Sn�� 4@%E���!?�mQ��@�6vtΟٿ73��؞�@�nS� 4@]��Ā�!?� :�|�@�!���ٿC6�[�o�@)m�%Z4@��!? ��!��@��̤ٿ�|�O�c�@�oח4@�r�d��!?��:	�@��̤ٿ�|�O�c�@�oח4@�r�d��!?��:	�@��̤ٿ�|�O�c�@�oח4@�r�d��!?��:	�@��̤ٿ�|�O�c�@�oח4@�r�d��!?��:	�@��̤ٿ�|�O�c�@�oח4@�r�d��!?��:	�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@���d�ٿ�㙈n��@��� 4@�1N=��!?����9e�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@nɧ���ٿ �LA��@͸4d} 4@��	#ˏ!?HU��f�@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@$�'���ٿ�(�����@k��3@�����!?~�e!J��@��">:�ٿf�6r��@&�Qϰ�3@&4�ҏ!?���G��@��">:�ٿf�6r��@&�Qϰ�3@&4�ҏ!?���G��@��">:�ٿf�6r��@&�Qϰ�3@&4�ҏ!?���G��@��">:�ٿf�6r��@&�Qϰ�3@&4�ҏ!?���G��@a$�L�ٿk�r��@�4΃4@�HE�!?��2�~�@J|����ٿ��;`���@j@��A�3@o�2؏!?���cK��@J|����ٿ��;`���@j@��A�3@o�2؏!?���cK��@J|����ٿ��;`���@j@��A�3@o�2؏!?���cK��@J|����ٿ��;`���@j@��A�3@o�2؏!?���cK��@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@�3Q��ٿh��iC/�@�(:�r 4@���î�!?@l�ǩ�@G�+��ٿ���a�@�dc�� 4@���΢�!?���@�
�@G�+��ٿ���a�@�dc�� 4@���΢�!?���@�
�@G�+��ٿ���a�@�dc�� 4@���΢�!?���@�
�@G�+��ٿ���a�@�dc�� 4@���΢�!?���@�
�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@���ٿx��I�@;�o: 4@�tȹ�!?փ���@�@nv�K�ٿ�H����@�4@uJd���!?��*'���@u�pR�ٿ���9�@,?�|4@���K��!? ��X��@u�pR�ٿ���9�@,?�|4@���K��!? ��X��@�c\ؚٿsP���@��a 4@��A�!?!>��(�@�c\ؚٿsP���@��a 4@��A�!?!>��(�@�c\ؚٿsP���@��a 4@��A�!?!>��(�@�c\ؚٿsP���@��a 4@��A�!?!>��(�@��"�ٿ�ţ'X��@G�H 4@�X�O��!?WObdB��@��L��ٿ ��h	��@�`w�� 4@>Wӣ��!?_V����@��L��ٿ ��h	��@�`w�� 4@>Wӣ��!?_V����@��L��ٿ ��h	��@�`w�� 4@>Wӣ��!?_V����@��;��ٿg1s���@�2-��4@<xQ�!?��R�!/�@��;��ٿg1s���@�2-��4@<xQ�!?��R�!/�@��;��ٿg1s���@�2-��4@<xQ�!?��R�!/�@\���ٿ1]ZoG��@I�?˵4@@�<�!?�cV��@OV���ٿ�o���@��c�4@���v��!?QxtdN�@OV���ٿ�o���@��c�4@���v��!?QxtdN�@OV���ٿ�o���@��c�4@���v��!?QxtdN�@��t�ٿ�m�t��@#0�4@P���͏!?x��T���@��t�ٿ�m�t��@#0�4@P���͏!?x��T���@��t�ٿ�m�t��@#0�4@P���͏!?x��T���@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@�5Q�H�ٿ��s�2��@�c��4@X�я!?��|.��@	N}�s�ٿ�so�3D�@��.r4@~���Ə!?�kD��@%UbŨٿA�^��@��C4@+l���!?���k��@hb��8�ٿ?a9����@��ΫU4@ٴ����!?u:<���@hb��8�ٿ?a9����@��ΫU4@ٴ����!?u:<���@hb��8�ٿ?a9����@��ΫU4@ٴ����!?u:<���@hb��8�ٿ?a9����@��ΫU4@ٴ����!?u:<���@�8�} �ٿ5R�/^~�@|�&�P4@�����!?�_{q)�@�8�} �ٿ5R�/^~�@|�&�P4@�����!?�_{q)�@�8�} �ٿ5R�/^~�@|�&�P4@�����!?�_{q)�@�8�} �ٿ5R�/^~�@|�&�P4@�����!?�_{q)�@5����ٿPb��k��@h7��6 4@݋�!? ��2�@��	��ٿ�����@mCyc4@i;�Y�!?%KY��*�@��	��ٿ�����@mCyc4@i;�Y�!?%KY��*�@��qn=�ٿ} 'Z���@���W*4@ɷ�ޏ!?F	5���@��qn=�ٿ} 'Z���@���W*4@ɷ�ޏ!?F	5���@��R@�ٿ�V�@�Ӎ�4@���᷏!?T�&
�7�@��R@�ٿ�V�@�Ӎ�4@���᷏!?T�&
�7�@����ٿGiI��@fO� 4@��a��!?�������@r�P�ٿ��	-M�@'68�! 4@�j��|�!?¶jM)�@r�P�ٿ��	-M�@'68�! 4@�j��|�!?¶jM)�@r�P�ٿ��	-M�@'68�! 4@�j��|�!?¶jM)�@����ٿI��|�@-.��U�3@H��l�!?�dXZ�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@��c�ٿ���!���@f -�v�3@(����!?�(C��(�@�X�ٿ�8�Oą�@c�����3@
�ы?�!?��=�.�@�#��@�ٿ�G.{9Y�@�gy�� 4@4r��!?�j�o��@�5�B�ٿiǇ͟�@�[�C�4@���b��!?��mm��@�5�B�ٿiǇ͟�@�[�C�4@���b��!?��mm��@�5�B�ٿiǇ͟�@�[�C�4@���b��!?��mm��@�5�B�ٿiǇ͟�@�[�C�4@���b��!?��mm��@Ŀ�+�ٿq27J�@�f�g�3@�D6��!?"g�GA�@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@eCΣٿ�N�����@�d�ؠ4@��1���!?VC��:��@qď��ٿke.���@	B� 4@�-p��!?X��A-��@qď��ٿke.���@	B� 4@�-p��!?X��A-��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@"Z��ٿ�̏�3%�@8o��3�3@z�޽�!?fp��@��?��ٿg�ʡ�;�@���� 4@��z���!?a����@��?��ٿg�ʡ�;�@���� 4@��z���!?a����@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@	~��ݝٿkge(��@7�E�3@h1q��!?�O!Q�@�D�XѣٿWOU�H��@'��@�3@�oG�e�!?��վ��@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@h�����ٿ��EG��@�	>��3@T�~���!?'�W���@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@D�(SA�ٿޕ�~���@�B� 4@���Ɲ�!?�?r��E�@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�>�V�ٿ/�ܵ��@�ۿ
4@7���z�!?��65��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�`�P�ٿLgB���@�(�@�4@�d#ᕏ!?d'��>��@�����ٿAi�dd��@R#u4L4@��;~��!?�N�P��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@0���ٿ�/鶶��@�M�%4@��)��!?��`��@�KE�۟ٿ�d�Ì�@��.� 4@�o#/��!?�|<�e�@�KE�۟ٿ�d�Ì�@��.� 4@�o#/��!?�|<�e�@�S��ٿ��t���@�z�� 4@��E3��!?H̑�UJ�@�S��ٿ��t���@�z�� 4@��E3��!?H̑�UJ�@&�i���ٿe{���@���Z�3@�`�͏!?^&��@�P�9Ѡٿ�� ���@�8�?�3@wB5���!?����5��@�P�9Ѡٿ�� ���@�8�?�3@wB5���!?����5��@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@}(f9�ٿ����0�@F�m��3@���ҳ�!?L�w��<�@�Q�ٿ>\�"���@M �h��3@�oP2]�!?
��r>.�@���ˤٿ@ܿh2�@q�U� 4@lSm�f�!?d�Vx���@�%�ťٿb���El�@sP�� 4@�?�!?,7�7?��@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@S\�4�ٿt8���@�%����3@�ǥ_?�!?�R�sj�@�K&�ܡٿVF�r"��@n��Ķ�3@�~�^�!?��>���@������ٿ�f,��@����!�3@/XJ�[�!?�t��6�@������ٿ�f,��@����!�3@/XJ�[�!?�t��6�@&�j�J�ٿ'�!Ŗd�@�_�g4@F��8%�!?���mo��@��A���ٿ��l!f�@��T���3@"Uueb�!?�0I�&)�@��A���ٿ��l!f�@��T���3@"Uueb�!?�0I�&)�@���M�ٿo#W���@�oP3��3@h���j�!?wL��@���M�ٿo#W���@�oP3��3@h���j�!?wL��@���M�ٿo#W���@�oP3��3@h���j�!?wL��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@���~l�ٿ��K~��@I�pb�3@SPdZ�!?�j�N��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@o�2�ٿ��a�2��@�e�3@��{J�!?HX}r:��@��8r�ٿ���#F��@�>q�_4@�q噶�!?Y�l���@���R�ٿ�KT�r�@�t�U� 4@��`���!?)�3� �@���R�ٿ�KT�r�@�t�U� 4@��`���!?)�3� �@���R�ٿ�KT�r�@�t�U� 4@��`���!?)�3� �@���R�ٿ�KT�r�@�t�U� 4@��`���!?)�3� �@���R�ٿ�KT�r�@�t�U� 4@��`���!?)�3� �@`�`10�ٿz�{v\��@�( 4@���ߣ�!?��3�@`�`10�ٿz�{v\��@�( 4@���ߣ�!?��3�@`�`10�ٿz�{v\��@�( 4@���ߣ�!?��3�@��dM�ٿ��
_q�@�K�uG4@������!?�V�o�f�@��dM�ٿ��
_q�@�K�uG4@������!?�V�o�f�@��dM�ٿ��
_q�@�K�uG4@������!?�V�o�f�@��dM�ٿ��
_q�@�K�uG4@������!?�V�o�f�@u�ć�ٿsv��#d�@�.`j 4@@9��!?0m��rs�@u�ć�ٿsv��#d�@�.`j 4@@9��!?0m��rs�@u�ć�ٿsv��#d�@�.`j 4@@9��!?0m��rs�@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@P�Ybs�ٿ���gm�@�^����3@1��2
�!?�j���@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@G��i�ٿ���P��@0���� 4@�gVݏ!?��� ��@�f5ƥ�ٿ�Ns"4��@Yomؾ�3@ҦP��!?&��n��@�f5ƥ�ٿ�Ns"4��@Yomؾ�3@ҦP��!?&��n��@�n5ҭ�ٿKBq�m�@�uI��3@��a~��!?��{���@�n5ҭ�ٿKBq�m�@�uI��3@��a~��!?��{���@��{*g�ٿ�=Si?��@5�j�=4@9�W�!?�ϲ�)�@��{*g�ٿ�=Si?��@5�j�=4@9�W�!?�ϲ�)�@��{*g�ٿ�=Si?��@5�j�=4@9�W�!?�ϲ�)�@��{*g�ٿ�=Si?��@5�j�=4@9�W�!?�ϲ�)�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@�7u�ٿ�����@J�p74@�b�!?S,�R�D�@��曧ٿv��M3��@�W�04@�O�k�!?��i�@��曧ٿv��M3��@�W�04@�O�k�!?��i�@��曧ٿv��M3��@�W�04@�O�k�!?��i�@��曧ٿv��M3��@�W�04@�O�k�!?��i�@��曧ٿv��M3��@�W�04@�O�k�!?��i�@Q�k�S�ٿ�=��О�@�ڑ� 4@�ܣ�!?�,��)�@Q�k�S�ٿ�=��О�@�ڑ� 4@�ܣ�!?�,��)�@)a�,:�ٿ&/�E;��@�N;6!4@�|F�Տ!?=��a2�@)a�,:�ٿ&/�E;��@�N;6!4@�|F�Տ!?=��a2�@��Ѱ��ٿ�CA�e��@E��4@}����!?Ŭ܅?��@�L��N�ٿD+��+�@��}��4@b/����!?�b�f�@�@�L��N�ٿD+��+�@��}��4@b/����!?�b�f�@�@�L��N�ٿD+��+�@��}��4@b/����!?�b�f�@�@�L��N�ٿD+��+�@��}��4@b/����!?�b�f�@�@�L��N�ٿD+��+�@��}��4@b/����!?�b�f�@�@�KX��ٿ� Q��k�@�{�_} 4@5�_2��!?n^T�H�@�KX��ٿ� Q��k�@�{�_} 4@5�_2��!?n^T�H�@�KX��ٿ� Q��k�@�{�_} 4@5�_2��!?n^T�H�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@L�7{�ٿ���8fd�@6/o 4@1:[!8�!?�X5��0�@�,��ٿ������@�I|O��3@�)"��!?��6��L�@z�����ٿ�PJ`�l�@J�X͢4@l���!?'�����@z�����ٿ�PJ`�l�@J�X͢4@l���!?'�����@z�����ٿ�PJ`�l�@J�X͢4@l���!?'�����@z�����ٿ�PJ`�l�@J�X͢4@l���!?'�����@	%��I�ٿ�B.�(��@;�Ϧ��3@#�aX�!?�L�� �@	%��I�ٿ�B.�(��@;�Ϧ��3@#�aX�!?�L�� �@	%��I�ٿ�B.�(��@;�Ϧ��3@#�aX�!?�L�� �@�΃�|�ٿ[�D��@X�C`�3@�rw��!?����@�۸N{�ٿ��ĶJ��@�8�x�3@�j���!?~�� ��@}b��ٿ�m�gL��@���2�3@d��fǏ!?�7��i�@}b��ٿ�m�gL��@���2�3@d��fǏ!?�7��i�@}b��ٿ�m�gL��@���2�3@d��fǏ!?�7��i�@���99�ٿ�s�-��@��!�P�3@��P�4�!?=��K�@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@��^��ٿ�  ǡ�@e�ca" 4@N����!?W+x���@�\݋��ٿVz4�G��@X��4@rư�!?]4O����@�\݋��ٿVz4�G��@X��4@rư�!?]4O����@';U��ٿ}p���@??O�D4@dVx!?p^<�_��@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@M�f�T�ٿ�s|�@�@	�� 4@�>M��!?�(��J�@;{���ٿGlTJ��@���	��3@"H^�܏!?{��4��@���;�ٿS��n!�@X���4@x	���!?��[���@���;�ٿS��n!�@X���4@x	���!?��[���@���;�ٿS��n!�@X���4@x	���!?��[���@���;�ٿS��n!�@X���4@x	���!?��[���@���;�ٿS��n!�@X���4@x	���!?��[���@t���ٿZ�'6�@�����4@�q	�!? ��.S��@, +��ٿ���f��@�g	1� 4@�����!?(���@��@, +��ٿ���f��@�g	1� 4@�����!?(���@��@, +��ٿ���f��@�g	1� 4@�����!?(���@��@����ٿ\�Pz�@�B>g]4@\��r�!?	�|1��@����ٿ\�Pz�@�B>g]4@\��r�!?	�|1��@����ٿ\�Pz�@�B>g]4@\��r�!?	�|1��@zX}�d�ٿ�X3�Q�@gR
�n4@�㣛��!?�w`�W��@zX}�d�ٿ�X3�Q�@gR
�n4@�㣛��!?�w`�W��@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@K��)�ٿ0q��J�@�,t���3@���Y�!?x)/���@4}��?�ٿ��O���@�aB\�3@AP(+�!?@�An�]�@4}��?�ٿ��O���@�aB\�3@AP(+�!?@�An�]�@4}��?�ٿ��O���@�aB\�3@AP(+�!?@�An�]�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@$����ٿ��7���@F%*4W4@n���l�!?t@']i}�@H����ٿ Z�W��@�v
���3@3��l�!?�EZ���@H����ٿ Z�W��@�v
���3@3��l�!?�EZ���@H����ٿ Z�W��@�v
���3@3��l�!?�EZ���@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@&A���ٿ��<�?�@ì/�[�3@�ޘ���!?�)�����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@�	��ٿH��˲��@8�겍4@)�<=�!?�Hh����@��Be�ٿK��b���@1�}�4@�K�@�!?qG2a��@I'����ٿ�b�(�x�@A�|� 4@�o�ja�!?�d6V���@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@E�`?�ٿ���)��@j��{U 4@
�p�e�!?�	Vje�@-U��G�ٿO�h"��@�f0� 4@�0�p��!?c���5�@-U��G�ٿO�h"��@�f0� 4@�0�p��!?c���5�@�����ٿ%����:�@.���� 4@P�L�Ə!?��F��@�����ٿ%����:�@.���� 4@P�L�Ə!?��F��@�����ٿ%����:�@.���� 4@P�L�Ə!?��F��@�����ٿ%����:�@.���� 4@P�L�Ə!?��F��@�����ٿ%����:�@.���� 4@P�L�Ə!?��F��@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@ب�uǢٿ����7��@Y�b7� 4@�����!?��fW-�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@�����ٿ,��9��@�u*�� 4@�MEA�!?��lO�@j�őx�ٿv��*�l�@9K��}�3@�5hr�!?h�R`��@j�őx�ٿv��*�l�@9K��}�3@�5hr�!?h�R`��@j�őx�ٿv��*�l�@9K��}�3@�5hr�!?h�R`��@j�őx�ٿv��*�l�@9K��}�3@�5hr�!?h�R`��@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@{ÌȆ�ٿ���U��@x�x,�3@F����!?
�j֜�@���1J�ٿD�HI�i�@Y|��3@	?
�ڏ!?�(����@���1J�ٿD�HI�i�@Y|��3@	?
�ڏ!?�(����@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@[��ѡٿ�{�8��@Ė�P�3@�*79��!?�n�[���@`���ƨٿ��~2;��@׍�4@� ��!?����@`���ƨٿ��~2;��@׍�4@� ��!?����@`���ƨٿ��~2;��@׍�4@� ��!?����@5��Ԭٿ��.)x��@sR�`R4@�`�J��!?X"��@ؚ�<��ٿ�a�P�@�j A��3@�����!?y�"��@ؚ�<��ٿ�a�P�@�j A��3@�����!?y�"��@ؚ�<��ٿ�a�P�@�j A��3@�����!?y�"��@�I�0j�ٿ�����@��]4@nP�.��!?,g"�@�I�0j�ٿ�����@��]4@nP�.��!?,g"�@�I�0j�ٿ�����@��]4@nP�.��!?,g"�@�I�0j�ٿ�����@��]4@nP�.��!?,g"�@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@	�o.�ٿś��5]�@��� 9 4@�r*���!?�����@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@�pv��ٿ�}Qh�@P�MO 4@�J�h�!?�C�7���@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@"�i|ԥٿ��Q�@�YiL 4@��2�͏!?����ܨ�@H*~d�ٿ�e�U�{�@Y��?' 4@v.ő��!?�Uw�`��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@C�'��ٿ�O�5�;�@
���3@i1=ҏ!?�U�S��@�?�ٿ�φ��_�@\��I"�3@��N���!?��Ց�@�?�ٿ�φ��_�@\��I"�3@��N���!?��Ց�@�?�ٿ�φ��_�@\��I"�3@��N���!?��Ց�@j�$���ٿY��v�@�q�h9�3@��V�!?oi��f�@j�$���ٿY��v�@�q�h9�3@��V�!?oi��f�@j�$���ٿY��v�@�q�h9�3@��V�!?oi��f�@{���ٿ�(�����@;-�Ea�3@���S�!?�Hd�u��@{���ٿ�(�����@;-�Ea�3@���S�!?�Hd�u��@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@.R~��ٿ�ވ��L�@zov�4@Iv.���!?g�/�@���֞ٿ@>���@���z4@�Y�똏!?#���%��@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@I�a���ٿ~�8���@��o4@�c���!?�%(`�<�@	��=��ٿN;>-�@C-���3@�y�B�!?	��G3	�@���^�ٿ�"�!ް�@�� 4@��tu�!?%cbӾ��@Un���ٿ+قM��@Ld�� 4@�y�8��!?ϐ����@Un���ٿ+قM��@Ld�� 4@�y�8��!?ϐ����@m7ꓖ�ٿ�F�o���@~p��a4@@A�ޏ!?���u���@m7ꓖ�ٿ�F�o���@~p��a4@@A�ޏ!?���u���@m7ꓖ�ٿ�F�o���@~p��a4@@A�ޏ!?���u���@dLҥ�ٿ��wX��@�S�.�4@R�ҏ�!?bM;X�^�@+T�Ec�ٿ|�G����@ȑ�4� 4@&ȏ!?Z}�t;�@+T�Ec�ٿ|�G����@ȑ�4� 4@&ȏ!?Z}�t;�@�;���ٿ�J�(��@�ꅲ	4@�rWa؏!?��2�@�;���ٿ�J�(��@�ꅲ	4@�rWa؏!?��2�@�;���ٿ�J�(��@�ꅲ	4@�rWa؏!?��2�@�;���ٿ�J�(��@�ꅲ	4@�rWa؏!?��2�@3�T��ٿ�3R~D��@k����3@d[���!?e+|�.;�@3�T��ٿ�3R~D��@k����3@d[���!?e+|�.;�@tJ��4�ٿ��u��:�@;���� 4@�6��!?{�7� h�@tJ��4�ٿ��u��:�@;���� 4@�6��!?{�7� h�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@B;c���ٿ��*|��@��Z 4@E��ð�!?��[�/v�@j�;��ٿ	J�&8`�@����o 4@gcW���!?36�A}}�@j�;��ٿ	J�&8`�@����o 4@gcW���!?36�A}}�@j�;��ٿ	J�&8`�@����o 4@gcW���!?36�A}}�@Sf$¢ٿ÷��D�@�S4@z��~��!?GU�16��@Sf$¢ٿ÷��D�@�S4@z��~��!?GU�16��@Sf$¢ٿ÷��D�@�S4@z��~��!?GU�16��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@���ٿ�<j��@�V�� 4@��ݜ�!?!���r��@[=�x�ٿYڷf��@��� ��3@��{J��!?$ufD��@[=�x�ٿYڷf��@��� ��3@��{J��!?$ufD��@[=�x�ٿYڷf��@��� ��3@��{J��!?$ufD��@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@w��-0�ٿRI$�p�@�q~��4@�n�!?�������@
xN/��ٿ��|���@Y��� 4@A�L���!?��Z�LI�@
xN/��ٿ��|���@Y��� 4@A�L���!?��Z�LI�@v�3�~�ٿ1��a*�@��2�� 4@������!?8�N~;6�@v�3�~�ٿ1��a*�@��2�� 4@������!?8�N~;6�@�T<��ٿ'�	s2�@s��6 4@9:�h��!?��!lc��@?����ٿº�]��@���4@h��]��!?w�Y�s�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@P~���ٿ���Z��@?���z4@�x���!?ye)_�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�<�ŝٿ�J���@�4u	4@�{�`�!?�|P�,�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�U��}�ٿX��ztW�@-�/ 4@!��!?����4�@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@�Ni��ٿH�@*/\�@���4@ړ�8z�!?mJ{�i��@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@p-�.�ٿIu����@�Z�`��3@�[;���!?z��)�5�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@��͐�ٿ�X���H�@Ɨ�4@W���!?j�*�	�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@����ٿ�|([��@
P S]4@F�p�!?�<��*�@�1���ٿ�Zt�L�@��վ� 4@�x�(��!?�ʥq<V�@�1���ٿ�Zt�L�@��վ� 4@�x�(��!?�ʥq<V�@�1���ٿ�Zt�L�@��վ� 4@�x�(��!?�ʥq<V�@�1���ٿ�Zt�L�@��վ� 4@�x�(��!?�ʥq<V�@�ӑ�ٿ�l(,��@����	 4@�X�J�!?H�2{��@�ӑ�ٿ�l(,��@����	 4@�X�J�!?H�2{��@�ӑ�ٿ�l(,��@����	 4@�X�J�!?H�2{��@Z[�ٿw�o��@K���� 4@���+��!?7�����@Z[�ٿw�o��@K���� 4@���+��!?7�����@Z[�ٿw�o��@K���� 4@���+��!?7�����@Z[�ٿw�o��@K���� 4@���+��!?7�����@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@��j!�ٿ��ǵ�@�#��4@vaĲ�!?YT��>��@c�v���ٿry����@m�"S 4@F��d��!?{���l�@c�v���ٿry����@m�"S 4@F��d��!?{���l�@c�v���ٿry����@m�"S 4@F��d��!?{���l�@c�v���ٿry����@m�"S 4@F��d��!?{���l�@Z��ٿ��Ĝ��@鞫2k 4@�1H��!?�ܤ���@Z��ٿ��Ĝ��@鞫2k 4@�1H��!?�ܤ���@�(b�Q�ٿ�:K�Z��@�g��
�3@��>Wޏ!?>����@�(b�Q�ٿ�:K�Z��@�g��
�3@��>Wޏ!?>����@�(b�Q�ٿ�:K�Z��@�g��
�3@��>Wޏ!?>����@�(b�Q�ٿ�:K�Z��@�g��
�3@��>Wޏ!?>����@�(b�Q�ٿ�:K�Z��@�g��
�3@��>Wޏ!?>����@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@E ����ٿ�bq�ռ�@�����3@�b)��!?�1�~;T�@x�%�ٿ�m��@�˗�,4@e����!?���մ��@}z`��ٿ`#9W��@��z�� 4@���Bُ!?��_�R�@^R� �ٿ�:�)��@���H��3@Da�,��!?�0�����@^R� �ٿ�:�)��@���H��3@Da�,��!?�0�����@�'���ٿ8p���@�%?{�3@?a��!?LM^m>��@>�l��ٿ����@�Im�v�3@{<}��!?Z�z~9�@>�l��ٿ����@�Im�v�3@{<}��!?Z�z~9�@>�l��ٿ����@�Im�v�3@{<}��!?Z�z~9�@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@v~ ʵ�ٿ��1���@���\�4@�0PՏ!?�C��@u^3x�ٿ-��${�@uQP*4@'_�Q��!?����^�@u^3x�ٿ-��${�@uQP*4@'_�Q��!?����^�@u^3x�ٿ-��${�@uQP*4@'_�Q��!?����^�@u^3x�ٿ-��${�@uQP*4@'_�Q��!?����^�@u^3x�ٿ-��${�@uQP*4@'_�Q��!?����^�@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@�vCH�ٿ���Pc�@\A�f4@ �ϤC�!?O,����@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@G13��ٿr�pu��@��I�4@��[��!? $��Y(�@t��t�ٿ�n���@�q|� 4@z�Ⱥ�!?7��#��@t��t�ٿ�n���@�q|� 4@z�Ⱥ�!?7��#��@t��t�ٿ�n���@�q|� 4@z�Ⱥ�!?7��#��@t��t�ٿ�n���@�q|� 4@z�Ⱥ�!?7��#��@���O�ٿ�c�P�p�@fOC�"4@	"|Џ!?��!8]8�@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@�M���ٿ�5�GP�@G �	 4@Pg��̏!?$ϡI��@��J쓠ٿ���o�@��I�04@��܇�!?q�"Ԭ�@9�6�i�ٿ�$Y�}�@��,[�4@쭶>��!?' ,�@���a �ٿ���|Y�@@N��4@:/n���!?2�63��@���a �ٿ���|Y�@@N��4@:/n���!?2�63��@�aa�ٿ�D��@�:i�4@7��zԏ!?sw���@s�E��ٿDd�JH��@�2��b4@�����!?�ϱ�D��@s�E��ٿDd�JH��@�2��b4@�����!?�ϱ�D��@Z���1�ٿw������@!�}k4@o4�?я!?���D$��@Z���1�ٿw������@!�}k4@o4�?я!?���D$��@Z���1�ٿw������@!�}k4@o4�?я!?���D$��@�)�\��ٿH*�=�@١՞� 4@ �)��!?6r�����@y���8�ٿ�==���@_��O��3@�;�$+�!?(f�-�A�@���vצٿ����o�@����3@q�$f�!?k1 ��3�@���vצٿ����o�@����3@q�$f�!?k1 ��3�@���vצٿ����o�@����3@q�$f�!?k1 ��3�@�f,M��ٿiʤ����@N�@�3@�@%r��!?�59(r��@�f,M��ٿiʤ����@N�@�3@�@%r��!?�59(r��@�f,M��ٿiʤ����@N�@�3@�@%r��!?�59(r��@iH+T�ٿi��Zx��@m��L��3@��*S��!?V�q�zn�@iH+T�ٿi��Zx��@m��L��3@��*S��!?V�q�zn�@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@=[ƽ4�ٿ�,����@���.� 4@��n;�!?u��#���@�'�&��ٿ��J�*��@r?f� 4@V��-я!?4Mص���@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@�$��t�ٿ�oا��@���*4@�:�$��!?���g�@C%���ٿŞ�����@y�� 4@q��%��!?%�;#H�@C%���ٿŞ�����@y�� 4@q��%��!?%�;#H�@�����ٿ�ͥ�e��@��^��3@X���!?�P.��@�����ٿ�ͥ�e��@��^��3@X���!?�P.��@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@��N��ٿ��P����@o�O>��3@r��h�!?�>�u]�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@G<ބt�ٿ�v2�
�@O��?4@���t�!?����JI�@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@�;��,�ٿR�;Z�@�쬏4@fr~���!?�	�A���@���I*�ٿ��Й�5�@�߇(4@N�ʏ!?�v%��@���I*�ٿ��Й�5�@�߇(4@N�ʏ!?�v%��@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@��(��ٿJuw�@�e�4@A��X�!?��6hX\�@2b\9{�ٿ�u$��I�@%
�y� 4@�_���!?䋯Q�D�@2b\9{�ٿ�u$��I�@%
�y� 4@�_���!?䋯Q�D�@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@핆�h�ٿ�N����@��[Q� 4@���h�!?$11m��@s�2�ٿG�D5��@u�W�4@Q��v�!?��&�o�@���ٿ$�ҁڣ�@��*S 4@n�z.ҏ!?��܁Q�@���ٿ$�ҁڣ�@��*S 4@n�z.ҏ!?��܁Q�@�s�P��ٿ�E�)V�@C��� �3@��%f�!?:��O��@�s�P��ٿ�E�)V�@C��� �3@��%f�!?:��O��@6�"J<�ٿ��y��9�@��̺��3@T�<HI�!?�Ä�dG�@�� �ٿI9oxH��@�a?�� 4@/�i;�!?]�)�z��@�� �ٿI9oxH��@�a?�� 4@/�i;�!?]�)�z��@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@��ٿ�m7Cd��@���7� 4@�'i�}�!?��T@.5�@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@L�be�ٿB8m�а�@2�6� 4@�T�p�!?H��/���@rjC��ٿ��!o���@�&��� 4@�YOm��!?��R%X�@rjC��ٿ��!o���@�&��� 4@�YOm��!?��R%X�@rjC��ٿ��!o���@�&��� 4@�YOm��!?��R%X�@rjC��ٿ��!o���@�&��� 4@�YOm��!?��R%X�@rjC��ٿ��!o���@�&��� 4@�YOm��!?��R%X�@C;��V�ٿ����@��\W4@�`�n��!?� ����@C;��V�ٿ����@��\W4@�`�n��!?� ����@���ȯٿUp#�K��@�1��4@d��-��!?l�1%F��@���ȯٿUp#�K��@�1��4@d��-��!?l�1%F��@���ȯٿUp#�K��@�1��4@d��-��!?l�1%F��@��Mt�ٿ���
=��@z{Z�� 4@4���ӏ!?]5��]��@��Mt�ٿ���
=��@z{Z�� 4@4���ӏ!?]5��]��@��Mt�ٿ���
=��@z{Z�� 4@4���ӏ!?]5��]��@�8gp�ٿ�w�y��@Qx 4@@m�z��!?"���u�@�U�Y�ٿ��>�B�@��V;4@;��y�!?PV�����@�U�Y�ٿ��>�B�@��V;4@;��y�!?PV�����@�U�Y�ٿ��>�B�@��V;4@;��y�!?PV�����@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@`d�/�ٿ�ƅ��@���b�4@= MÏ!?Vl��>�@��f�u�ٿk��ۂ��@�XĎ 4@� h"�!?w���)��@��f�u�ٿk��ۂ��@�XĎ 4@� h"�!?w���)��@��f�u�ٿk��ۂ��@�XĎ 4@� h"�!?w���)��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@�x�s�ٿf������@u�tO� 4@�d�׏!?���!R��@C��^�ٿ�tX���@��u��4@� C��!?���H��@C��^�ٿ�tX���@��u��4@� C��!?���H��@bU�Ѫٿӷ0�'��@�6O�4@TK;�Ϗ!?1?+`�O�@�wS�C�ٿ,��X���@�P�o� 4@�/��!?�Neg�@�wS�C�ٿ,��X���@�P�o� 4@�/��!?�Neg�@�wS�C�ٿ,��X���@�P�o� 4@�/��!?�Neg�@�wS�C�ٿ,��X���@�P�o� 4@�/��!?�Neg�@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@	��=f�ٿ�L�m�y�@׿�P4@� (���!?��1}��@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@��8�ٿq�&��i�@P:� 4@F*����!?�'t�h�@�#�ٿ�J�t���@�s��n�3@���!?�����@s(�ڽ�ٿ�Vߤ��@�YF 4@���zϏ!?�I��!r�@s(�ڽ�ٿ�Vߤ��@�YF 4@���zϏ!?�I��!r�@s(�ڽ�ٿ�Vߤ��@�YF 4@���zϏ!?�I��!r�@s(�ڽ�ٿ�Vߤ��@�YF 4@���zϏ!?�I��!r�@Z���}�ٿ�<�%��@_J��. 4@:p*t��!?��-yJ�@Z���}�ٿ�<�%��@_J��. 4@:p*t��!?��-yJ�@^3�{�ٿ���/��@��� 4@��Qʩ�!?$ǭ���@���	�ٿ_4��߱�@��R�N4@��D'Џ!?��f[�@���	�ٿ_4��߱�@��R�N4@��D'Џ!?��f[�@���	�ٿ_4��߱�@��R�N4@��D'Џ!?��f[�@X����ٿ!�c���@�S��� 4@��N��!?\3ύ/�@X����ٿ!�c���@�S��� 4@��N��!?\3ύ/�@X����ٿ!�c���@�S��� 4@��N��!?\3ύ/�@X����ٿ!�c���@�S��� 4@��N��!?\3ύ/�@X����ٿ!�c���@�S��� 4@��N��!?\3ύ/�@��a�>�ٿĘ$�h6�@^�Lx4@C'~�|�!?o�̐�n�@��a�>�ٿĘ$�h6�@^�Lx4@C'~�|�!?o�̐�n�@��a�>�ٿĘ$�h6�@^�Lx4@C'~�|�!?o�̐�n�@��a�>�ٿĘ$�h6�@^�Lx4@C'~�|�!?o�̐�n�@��a�>�ٿĘ$�h6�@^�Lx4@C'~�|�!?o�̐�n�@ ��&��ٿ�����@�#�%4@H���h�!?\E\�'��@ ��&��ٿ�����@�#�%4@H���h�!?\E\�'��@ ��&��ٿ�����@�#�%4@H���h�!?\E\�'��@ ��&��ٿ�����@�#�%4@H���h�!?\E\�'��@ ��&��ٿ�����@�#�%4@H���h�!?\E\�'��@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@6��k@�ٿF���w�@Yt�6 4@�9��!?0�����@L�t�j�ٿ �$!���@cm^��3@��d���!?���`�@L�t�j�ٿ �$!���@cm^��3@��d���!?���`�@L�t�j�ٿ �$!���@cm^��3@��d���!?���`�@L�t�j�ٿ �$!���@cm^��3@��d���!?���`�@L�t�j�ٿ �$!���@cm^��3@��d���!?���`�@}���ٿm�����@��5��3@����R�!?������@�nwH�ٿW���Z�@_�2��3@�d�W��!?�"h��@�nwH�ٿW���Z�@_�2��3@�d�W��!?�"h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@?��)�ٿ���X�@�����3@g�tЏ!?位�h��@�բ	�ٿ_�v*�@So��L�3@f>�g�!?P� ���@�բ	�ٿ_�v*�@So��L�3@f>�g�!?P� ���@�բ	�ٿ_�v*�@So��L�3@f>�g�!?P� ���@�բ	�ٿ_�v*�@So��L�3@f>�g�!?P� ���@�`�*ܛٿ�q;�G�@P+�x7 4@�ۤ���!?��5�4�@�`�*ܛٿ�q;�G�@P+�x7 4@�ۤ���!?��5�4�@�N�VרٿL秸\�@D�̝��3@�ڎŏ!?��XÅ�@�N�VרٿL秸\�@D�̝��3@�ڎŏ!?��XÅ�@�N�VרٿL秸\�@D�̝��3@�ڎŏ!?��XÅ�@�N�VרٿL秸\�@D�̝��3@�ڎŏ!?��XÅ�@-X�íٿ;�0�A�@LC1�v�3@Ĕ/�l�!?�#AU��@-X�íٿ;�0�A�@LC1�v�3@Ĕ/�l�!?�#AU��@-X�íٿ;�0�A�@LC1�v�3@Ĕ/�l�!?�#AU��@�:���ٿ��f�2H�@�l.x��3@G���!?�����@�:���ٿ��f�2H�@�l.x��3@G���!?�����@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@�_���ٿH�ZH�@�����3@,F����!?�  >��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@*Cu;�ٿa-���@�P�Q4@��{��!?��C��@
����ٿ����F�@U/)y 4@��!?��wX��@
����ٿ����F�@U/)y 4@��!?��wX��@
����ٿ����F�@U/)y 4@��!?��wX��@
����ٿ����F�@U/)y 4@��!?��wX��@*2��T�ٿ9y��@��=��3@Ƌ-�!?Ak�%[�@*2��T�ٿ9y��@��=��3@Ƌ-�!?Ak�%[�@*2��T�ٿ9y��@��=��3@Ƌ-�!?Ak�%[�@����ٿW+ �l�@���WO�3@�|#��!?:})�@����ٿW+ �l�@���WO�3@�|#��!?:})�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�5�_�ٿ��`2��@�f��W�3@<�'�ۏ!?��&��1�@�1��>�ٿ!�Rt[��@����4@9�b���!?7s�>*�@�1��>�ٿ!�Rt[��@����4@9�b���!?7s�>*�@�1��>�ٿ!�Rt[��@����4@9�b���!?7s�>*�@�1��>�ٿ!�Rt[��@����4@9�b���!?7s�>*�@�1��>�ٿ!�Rt[��@����4@9�b���!?7s�>*�@��Aܱٿ�oM^�@�[,֫�3@��ק�!?�q����@��Aܱٿ�oM^�@�[,֫�3@��ק�!?�q����@��Aܱٿ�oM^�@�[,֫�3@��ק�!?�q����@��Aܱٿ�oM^�@�[,֫�3@��ק�!?�q����@�[{��ٿ�n�d���@�y̅G 4@�T� ��!?Js��@�[{��ٿ�n�d���@�y̅G 4@�T� ��!?Js��@�[{��ٿ�n�d���@�y̅G 4@�T� ��!?Js��@�[{��ٿ�n�d���@�y̅G 4@�T� ��!?Js��@�[{��ٿ�n�d���@�y̅G 4@�T� ��!?Js��@q�v�ٿ/�N�}��@r��{$4@�VL�!?��N�s�@q�v�ٿ/�N�}��@r��{$4@�VL�!?��N�s�@q�v�ٿ/�N�}��@r��{$4@�VL�!?��N�s�@q�v�ٿ/�N�}��@r��{$4@�VL�!?��N�s�@�A{�]�ٿ��u��@M�"�� 4@�@�[�!?�Sbn��@�A{�]�ٿ��u��@M�"�� 4@�@�[�!?�Sbn��@�A{�]�ٿ��u��@M�"�� 4@�@�[�!?�Sbn��@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@��HD8�ٿ���h�@w�S=��3@ `a��!?H~�����@5��w��ٿBiQ�D��@�nP4@��s���!?T�ؽ5�@��M��ٿ`6�D)�@LN�Z4@���z�!?^�?Q3��@�|5֧ٿ��Bd���@gp�k� 4@ϫ|qq�!?�ؕ���@�|5֧ٿ��Bd���@gp�k� 4@ϫ|qq�!?�ؕ���@G�Ǫ��ٿs:*U���@�5Y�4@��4�!?Y=a��@��P
y�ٿ�!��@NBUǡ4@!��6\�!?R<Zo��@a�ۋ�ٿ|�o�ե�@�f�^�4@��]��!?7���g��@a�ۋ�ٿ|�o�ե�@�f�^�4@��]��!?7���g��@a�ۋ�ٿ|�o�ե�@�f�^�4@��]��!?7���g��@a�ۋ�ٿ|�o�ե�@�f�^�4@��]��!?7���g��@ȭ�ٿ�){l��@��wL4@Yy�>��!?�K�lH��@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@
x�ٿ��|)ϸ�@%��4@��ޏ!?���� 5�@��h�ٿM�#v���@{)�d�4@c3a��!?ZZ0����@���x��ٿWu�k�@mQӨ04@P��	�!?�ȵ��@���x��ٿWu�k�@mQӨ04@P��	�!?�ȵ��@���x��ٿWu�k�@mQӨ04@P��	�!?�ȵ��@E�O<�ٿE	]q�@z4��� 4@+�4�!?,W�
Yp�@E�O<�ٿE	]q�@z4��� 4@+�4�!?,W�
Yp�@E�O<�ٿE	]q�@z4��� 4@+�4�!?,W�
Yp�@E�O<�ٿE	]q�@z4��� 4@+�4�!?,W�
Yp�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@�-����ٿ�M�*��@G���4@��D�!?�M��ww�@ٛF���ٿZ����N�@똢� 4@S��p9�!?%�>П�@ٛF���ٿZ����N�@똢� 4@S��p9�!?%�>П�@ٛF���ٿZ����N�@똢� 4@S��p9�!?%�>П�@ʓ�=ͪٿ<Nb�>��@�m1�P�3@m��׏!?���]y�@H ˺�ٿ�,杂�@`��4@@�K/�!?��(Z�O�@H ˺�ٿ�,杂�@`��4@@�K/�!?��(Z�O�@H ˺�ٿ�,杂�@`��4@@�K/�!?��(Z�O�@H ˺�ٿ�,杂�@`��4@@�K/�!?��(Z�O�@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@�d�`y�ٿӜjZ|5�@��a� 4@��)��!?���%��@C�Z(^�ٿ�Q��O�@�-�3@K� Ȭ�!?��H���@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@=��ϝٿ�,6;��@�g���3@�4�곏!?��cL�@��2ۜٿ��Ic�e�@���d�3@�H�-��!?�k�o46�@��2ۜٿ��Ic�e�@���d�3@�H�-��!?�k�o46�@��2ۜٿ��Ic�e�@���d�3@�H�-��!?�k�o46�@���;�ٿ<��z�@���8�3@����u�!?vh����@���;�ٿ<��z�@���8�3@����u�!?vh����@���;�ٿ<��z�@���8�3@����u�!?vh����@���;�ٿ<��z�@���8�3@����u�!?vh����@���;�ٿ<��z�@���8�3@����u�!?vh����@�XD(��ٿ�Hў��@�t(���3@C�;Bt�!?�8x��@�XD(��ٿ�Hў��@�t(���3@C�;Bt�!?�8x��@�XD(��ٿ�Hў��@�t(���3@C�;Bt�!?�8x��@�XD(��ٿ�Hў��@�t(���3@C�;Bt�!?�8x��@�XD(��ٿ�Hў��@�t(���3@C�;Bt�!?�8x��@��C��ٿ�����u�@I����3@P��!?��9���@��C��ٿ�����u�@I����3@P��!?��9���@��C��ٿ�����u�@I����3@P��!?��9���@��C��ٿ�����u�@I����3@P��!?��9���@�T_��ٿ�gD�nG�@�u[�� 4@ ��L��!?=Bt'��@�O�B��ٿG���@�&<Z�4@�
l���!?81ş��@�O�B��ٿG���@�&<Z�4@�
l���!?81ş��@�fwD̩ٿ��+M��@�s�4@
�s9�!?������@����B�ٿ����=3�@��� 4@�"~�o�!?�`�N�A�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@������ٿ�m9�<�@+�h��4@m [{�!?�d��4�@˖K��ٿC�_��7�@y�:�4@xכֿ�!?�-�oP8�@˖K��ٿC�_��7�@y�:�4@xכֿ�!?�-�oP8�@˖K��ٿC�_��7�@y�:�4@xכֿ�!?�-�oP8�@˖K��ٿC�_��7�@y�:�4@xכֿ�!?�-�oP8�@3�=��ٿP��Ҷ��@�u��d4@��Z�!?�7 Z.��@3�=��ٿP��Ҷ��@�u��d4@��Z�!?�7 Z.��@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@t0�ٿ��,gkD�@�M]�� 4@�3\��!?�d_}�@��P��ٿ%(u���@O�%� 4@\��̏!?^jٜ�$�@��P��ٿ%(u���@O�%� 4@\��̏!?^jٜ�$�@'���#�ٿF�a=�@��Js�3@�(�:��!?V!���@'���#�ٿF�a=�@��Js�3@�(�:��!?V!���@'���#�ٿF�a=�@��Js�3@�(�:��!?V!���@M��\�ٿ��v��@�ҭ 4@�,Zu�!??Xf.��@L��殛ٿ:M�i�F�@���UF 4@��s�~�!?weR%
�@L��殛ٿ:M�i�F�@���UF 4@��s�~�!?weR%
�@ϸw�ٿy
���@pw�4` 4@�b�c��!?ϡ^Y�%�@ϸw�ٿy
���@pw�4` 4@�b�c��!?ϡ^Y�%�@�P��ٿ<�7}u�@���4@d�h��!?u�/����@�P��ٿ<�7}u�@���4@d�h��!?u�/����@�P��ٿ<�7}u�@���4@d�h��!?u�/����@�P��ٿ<�7}u�@���4@d�h��!?u�/����@�P��ٿ<�7}u�@���4@d�h��!?u�/����@�P��ٿ<�7}u�@���4@d�h��!?u�/����@n��$�ٿٮ5s��@e��~�3@h�R���!?�R����@n��$�ٿٮ5s��@e��~�3@h�R���!?�R����@n��$�ٿٮ5s��@e��~�3@h�R���!?�R����@n��$�ٿٮ5s��@e��~�3@h�R���!?�R����@n��$�ٿٮ5s��@e��~�3@h�R���!?�R����@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@��ٿ$pk/��@~��4@Au�妏!?%��Y��@�~s�Ʃٿ�̖�,�@ ��m84@ٍ�ҏ!?
�QI���@�~s�Ʃٿ�̖�,�@ ��m84@ٍ�ҏ!?
�QI���@�~s�Ʃٿ�̖�,�@ ��m84@ٍ�ҏ!?
�QI���@�~s�Ʃٿ�̖�,�@ ��m84@ٍ�ҏ!?
�QI���@� ��&�ٿ2�q���@K?5�� 4@B%r�l�!?������@� ��&�ٿ2�q���@K?5�� 4@B%r�l�!?������@]R :�ٿ�������@��S� 4@�Ї0K�!?�^,g���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@��[�ѝٿ͖���@�n%� 4@y��!R�!?�r	���@�����ٿ���r�@{��^ 4@��U��!?�njފ�@��*�ٿ�LG��(�@(!�{4@)��0��!?��� ��@��*�ٿ�LG��(�@(!�{4@)��0��!?��� ��@��*�ٿ�LG��(�@(!�{4@)��0��!?��� ��@L�f�K�ٿ�
,m&%�@�c�5a 4@�	;��!?�B�M[��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@ �"77�ٿ�p/*<!�@��a�
 4@|37��!?c�q=��@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@E���\�ٿD��T �@���b� 4@˪T�!?~�#jZo�@����ٿ�;����@�Ƌ��4@��+���!?>����+�@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@~JḴ�ٿ����D@�@UG4*4@8� ��!?�nN���@��tɰ�ٿ�"u��k�@XR�9Z�3@4y �ӏ!?��y��@��tɰ�ٿ�"u��k�@XR�9Z�3@4y �ӏ!?��y��@��tɰ�ٿ�"u��k�@XR�9Z�3@4y �ӏ!?��y��@�f����ٿ~���oY�@�+-/�3@�X?��!?3���hs�@�f����ٿ~���oY�@�+-/�3@�X?��!?3���hs�@�f����ٿ~���oY�@�+-/�3@�X?��!?3���hs�@�f����ٿ~���oY�@�+-/�3@�X?��!?3���hs�@�f����ٿ~���oY�@�+-/�3@�X?��!?3���hs�@r9�רٿ�6d����@��2��3@���!?�|����@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@:c1�{�ٿ��P�=n�@&����3@#A��!?��"<��@�KVEśٿZ���@����q 4@�51��!?.��f�@�KVEśٿZ���@����q 4@�51��!?.��f�@�KVEśٿZ���@����q 4@�51��!?.��f�@�KVEśٿZ���@����q 4@�51��!?.��f�@��9{<�ٿ `|�>�@<R�D�4@�vn��!?j��bR�@�c����ٿ=�n0P�@���) 4@+��劏!?6˶B~q�@�c����ٿ=�n0P�@���) 4@+��劏!?6˶B~q�@@	��ٿ��E�?^�@S�+�4@�}>�Q�!?,��E�v�@@	��ٿ��E�?^�@S�+�4@�}>�Q�!?,��E�v�@���˦ٿ|m�}���@#}M 4@�6�P�!?�hQ���@.#쪑�ٿ �	���@-T�<4@��E�c�!?hI�K�@.#쪑�ٿ �	���@-T�<4@��E�c�!?hI�K�@`׍�өٿi(�5���@���P� 4@:.�x��!?2_�Xu��@`׍�өٿi(�5���@���P� 4@:.�x��!?2_�Xu��@`׍�өٿi(�5���@���P� 4@:.�x��!?2_�Xu��@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@@�̓��ٿ�cd�G[�@�t#S� 4@�i"�!?�����@�I.wݢٿF2ߍ�l�@5ND�4@����!?~��Q���@�҅d��ٿ�%0����@�%�?T 4@�2%	��!?�bh�6�@�҅d��ٿ�%0����@�%�?T 4@�2%	��!?�bh�6�@�҅d��ٿ�%0����@�%�?T 4@�2%	��!?�bh�6�@�,��ٿ=����@��oa� 4@�����!?(�@�L���ٿ�:����@Ǆg�R�3@�1#ך�!?��3\o3�@�L���ٿ�:����@Ǆg�R�3@�1#ך�!?��3\o3�@�L���ٿ�:����@Ǆg�R�3@�1#ך�!?��3\o3�@�L���ٿ�:����@Ǆg�R�3@�1#ך�!?��3\o3�@�L���ٿ�:����@Ǆg�R�3@�1#ך�!?��3\o3�@���ٿz�)�`u�@�^ysf 4@�/�|��!?ڋ�>\D�@���ٿz�)�`u�@�^ysf 4@�/�|��!?ڋ�>\D�@�� ���ٿZsu�@�:`�/4@~�w���!?�W�g3��@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@T-��`�ٿ�M����@iR�E�3@�����!?-�����@X�r��ٿ��%=�@�ギ4@���&i�!?)^����@X�r��ٿ��%=�@�ギ4@���&i�!?)^����@X�r��ٿ��%=�@�ギ4@���&i�!?)^����@X�r��ٿ��%=�@�ギ4@���&i�!?)^����@X�r��ٿ��%=�@�ギ4@���&i�!?)^����@�M圖�ٿ^�Dww��@�+ �� 4@+&�d�!?N�"W���@�M圖�ٿ^�Dww��@�+ �� 4@+&�d�!?N�"W���@�M圖�ٿ^�Dww��@�+ �� 4@+&�d�!?N�"W���@|	�O�ٿ��;��E�@]�%���3@PDƷ��!?����y�@|	�O�ٿ��;��E�@]�%���3@PDƷ��!?����y�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@�0��;�ٿ�����@eOd� 4@�[�3��!?��e:�K�@��6G�ٿ���w?��@�~]�4@�NNa��!?5_˫��@��6G�ٿ���w?��@�~]�4@�NNa��!?5_˫��@G�O���ٿ]�V��C�@<�܉4@O� ���!?������@G�O���ٿ]�V��C�@<�܉4@O� ���!?������@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@����K�ٿ�sV�G�@e�@r�4@�J�!?Y��d4V�@T��I��ٿ����q-�@Bx�,� 4@�`�A�!?�=��,�@T��I��ٿ����q-�@Bx�,� 4@�`�A�!?�=��,�@T��I��ٿ����q-�@Bx�,� 4@�`�A�!?�=��,�@Q�G���ٿbh_���@(M����3@�xđ0�!?�b>��@Q�G���ٿbh_���@(M����3@�xđ0�!?�b>��@q��l�ٿ�Ǘc��@޷ʑ��3@v��
�!?����IL�@q��l�ٿ�Ǘc��@޷ʑ��3@v��
�!?����IL�@q��l�ٿ�Ǘc��@޷ʑ��3@v��
�!?����IL�@A�'�ٿI� �\P�@[��'=�3@���Տ!?���B�@)b�B�ٿ��, ��@v�`,4@��'\i�!?l�F��7�@�v�PY�ٿ��^	z��@���L�4@ŵ=��!?@o�oB��@�v�PY�ٿ��^	z��@���L�4@ŵ=��!?@o�oB��@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@� "�ٿE�J���@H�1b� 4@��F٤�!?4��g���@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@��c�ٿ�@G���@�B�x� 4@��0Ï!?'`P��@[f�"=�ٿ_�_���@g3�� 4@��r�Ǐ!?�f��@U�Lt�ٿ+IǘT��@B�+��3@�4m
�!?��ԠM��@U�Lt�ٿ+IǘT��@B�+��3@�4m
�!?��ԠM��@U�Lt�ٿ+IǘT��@B�+��3@�4m
�!?��ԠM��@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@$G]��ٿ���{Ъ�@�BFq� 4@}{}�Տ!?�ƞ�8	�@/�JSV�ٿ+ܢ m�@��4%� 4@.�}��!?B�C����@�z�C�ٿ���<��@�_s���3@a��藏!?�se����@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�P��J�ٿ^	�t�@���W 4@嫰�!?������@�ZX�ٿ՛@%��@��V� 4@�Go��!?�E�,��@�ZX�ٿ՛@%��@��V� 4@�Go��!?�E�,��@�ZX�ٿ՛@%��@��V� 4@�Go��!?�E�,��@�ZX�ٿ՛@%��@��V� 4@�Go��!?�E�,��@�ZX�ٿ՛@%��@��V� 4@�Go��!?�E�,��@���糩ٿ��s:G��@&3:"14@o����!?�V���B�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@���V�ٿ��/=;�@1�7u4@^D���!?�r��D�@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@N�Q{�ٿ�y���@�wB� 4@�m����!?�P3�l��@�b��ٿ>	#����@���4@�����!?e[�m��@%�H�0�ٿ@_��Ս�@����� 4@{�?ڏ!?�H��o�@%�H�0�ٿ@_��Ս�@����� 4@{�?ڏ!?�H��o�@%�H�0�ٿ@_��Ս�@����� 4@{�?ڏ!?�H��o�@%�H�0�ٿ@_��Ս�@����� 4@{�?ڏ!?�H��o�@m@[ʲ�ٿy�v�zH�@B&�+��3@p��Տ!?��*e��@m@[ʲ�ٿy�v�zH�@B&�+��3@p��Տ!?��*e��@�<6��ٿ��Ԛ��@{?�t��3@k�t��!?�����U�@���١ٿ�f�*��@ȋ8�3@����$�!?+h�*�i�@���١ٿ�f�*��@ȋ8�3@����$�!?+h�*�i�@���١ٿ�f�*��@ȋ8�3@����$�!?+h�*�i�@���١ٿ�f�*��@ȋ8�3@����$�!?+h�*�i�@���١ٿ�f�*��@ȋ8�3@����$�!?+h�*�i�@7�Ջ�ٿTl�����@�̛�3@�p�ӏ!?Uꪲ"?�@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�'Q�ɫٿdO<-V=�@9�8�$�3@�0����!?r[Qe��@�wA���ٿ��|'�s�@C���` 4@�b��B�!?3�ZE6�@�wA���ٿ��|'�s�@C���` 4@�b��B�!?3�ZE6�@ې��ٿ��F���@p���� 4@:��L�!?<R�s�@Ǫٯ�ٿ���x �@+�\�3@�"b�!?�.��?��@Ǫٯ�ٿ���x �@+�\�3@�"b�!?�.��?��@Ǫٯ�ٿ���x �@+�\�3@�"b�!?�.��?��@Ǫٯ�ٿ���x �@+�\�3@�"b�!?�.��?��@����~�ٿi�@{��~]�3@0�d�!?��7���@����~�ٿi�@{��~]�3@0�d�!?��7���@�8�Ag�ٿ������@����3@l�V�ŏ!?
�U�>h�@�8�Ag�ٿ������@����3@l�V�ŏ!?
�U�>h�@�8�Ag�ٿ������@����3@l�V�ŏ!?
�U�>h�@3�ډ�ٿ F���@�����3@Z ���!?3G�)��@3�ډ�ٿ F���@�����3@Z ���!?3G�)��@K���f�ٿ���v��@��� 4@�����!?I?�����@K���f�ٿ���v��@��� 4@�����!?I?�����@��65w�ٿ3.��5��@=A�54@�?�X�!?����@��65w�ٿ3.��5��@=A�54@�?�X�!?����@��65w�ٿ3.��5��@=A�54@�?�X�!?����@��65w�ٿ3.��5��@=A�54@�?�X�!?����@.��'��ٿ�F�-j�@���`�4@(�
�S�!?�;f�9�@.��'��ٿ�F�-j�@���`�4@(�
�S�!?�;f�9�@�����ٿ�����t�@)��t 4@�'�}�!?`*u(�-�@�O�ٿ��o��@X�]���3@���"��!?d���� �@�O�ٿ��o��@X�]���3@���"��!?d���� �@�O�ٿ��o��@X�]���3@���"��!?d���� �@�O�ٿ��o��@X�]���3@���"��!?d���� �@�O�ٿ��o��@X�]���3@���"��!?d���� �@'?����ٿbه�{��@{����3@b�d���!?�w�u{�@'?����ٿbه�{��@{����3@b�d���!?�w�u{�@'?����ٿbه�{��@{����3@b�d���!?�w�u{�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@6���T�ٿЦ��i�@���m�3@/�Rn��!?>�MQ5g�@\���ٿ;��L$��@��h,� 4@v�e/o�!?�E��?�@\���ٿ;��L$��@��h,� 4@v�e/o�!?�E��?�@\���ٿ;��L$��@��h,� 4@v�e/o�!?�E��?�@\���ٿ;��L$��@��h,� 4@v�e/o�!?�E��?�@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@���L#�ٿ��f%[�@Ʈ]V1 4@<獦��!?�V�����@�[����ٿ���p�V�@�-!>�3@R�W'��!?��3S��@�[����ٿ���p�V�@�-!>�3@R�W'��!?��3S��@˕�F+�ٿ��la'��@|�ą 4@��l�!?��֋�l�@�	*+�ٿ�n�<P&�@��B]4@��m��!?��f���@�	*+�ٿ�n�<P&�@��B]4@��m��!?��f���@�	*+�ٿ�n�<P&�@��B]4@��m��!?��f���@�	*+�ٿ�n�<P&�@��B]4@��m��!?��f���@�	*+�ٿ�n�<P&�@��B]4@��m��!?��f���@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@��|��ٿ�GH��@�Tod'4@�R#W�!?R ���6�@ڄ��ٿ/Ny�-��@?^v�4@q,¶�!?Y��>��@ڄ��ٿ/Ny�-��@?^v�4@q,¶�!?Y��>��@ڄ��ٿ/Ny�-��@?^v�4@q,¶�!?Y��>��@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�2�}�ٿ�@u��@g��)M 4@���f�!?�f T�@�]u\F�ٿ}iP\z*�@/dx�E4@K���l�!?Lgڇ�C�@�]u\F�ٿ}iP\z*�@/dx�E4@K���l�!?Lgڇ�C�@�]u\F�ٿ}iP\z*�@/dx�E4@K���l�!?Lgڇ�C�@�]u\F�ٿ}iP\z*�@/dx�E4@K���l�!?Lgڇ�C�@�]u\F�ٿ}iP\z*�@/dx�E4@K���l�!?Lgڇ�C�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@����z�ٿ՜�9��@6��w��3@	��ܕ�!?��0$�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@�{�Ţ�ٿ)�٫U��@�ܰ�{�3@K�Π�!?�c�G5�@)}�Z�ٿ Bz� �@�	�&~�3@���̏!?�G����@)}�Z�ٿ Bz� �@�	�&~�3@���̏!?�G����@���'ԬٿӠ$J"��@���[�4@�JNo�!?;����@�hQk�ٿ���H��@ ���)4@���
�!?���w�X�@�hQk�ٿ���H��@ ���)4@���
�!?���w�X�@�hQk�ٿ���H��@ ���)4@���
�!?���w�X�@�hQk�ٿ���H��@ ���)4@���
�!?���w�X�@�R>��ٿ��Lf`�@GҢ}��3@���v�!?�W�s���@�E�d�ٿ������@�j�o 4@QY�H�!?Hgy�Gc�@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@a��̥ٿ�
uV���@K�q� 4@j~0@�!?���&��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@�6|�ٿ<	.IE�@a��v�3@wc,�!?G�,��@隫���ٿ!�H��@��S~�3@ےU���!?F��D�@隫���ٿ!�H��@��S~�3@ےU���!?F��D�@����ٿ�3��@'�d��3@8�L���!?>�/!!�@#�z^�ٿ�B#c��@j�{4@��mx��!?�ơp��@#�z^�ٿ�B#c��@j�{4@��mx��!?�ơp��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@��;ʨٿ�����@)-����3@ߖ��!?�=5;��@7��:��ٿ�X�J%��@�����3@ŉpw�!?���Q�@7��:��ٿ�X�J%��@�����3@ŉpw�!?���Q�@��K8�ٿj�=��@��3��3@�¥+��!?��ɴp�@��K8�ٿj�=��@��3��3@�¥+��!?��ɴp�@��K)�ٿ�ubTA�@	�h�4@��@�!?zI4���@��K)�ٿ�ubTA�@	�h�4@��@�!?zI4���@��K)�ٿ�ubTA�@	�h�4@��@�!?zI4���@��K)�ٿ�ubTA�@	�h�4@��@�!?zI4���@��K)�ٿ�ubTA�@	�h�4@��@�!?zI4���@�N��ٿ�B+$2�@R�<�4@�A����!?��x]\�@�N��ٿ�B+$2�@R�<�4@�A����!?��x]\�@�N��ٿ�B+$2�@R�<�4@�A����!?��x]\�@U*�ٿ�Wƶ��@&0��k 4@4`���!?�|z�}�@��(D,�ٿ(�D�Ѹ�@o|8���3@fR̏!?9܃�V�@��(D,�ٿ(�D�Ѹ�@o|8���3@fR̏!?9܃�V�@��(D,�ٿ(�D�Ѹ�@o|8���3@fR̏!?9܃�V�@��(D,�ٿ(�D�Ѹ�@o|8���3@fR̏!?9܃�V�@������ٿ�5� �U�@s�7\�3@�r��!?_!$���@������ٿ�5� �U�@s�7\�3@�r��!?_!$���@������ٿ�5� �U�@s�7\�3@�r��!?_!$���@������ٿ�5� �U�@s�7\�3@�r��!?_!$���@OYG;�ٿ�[� ��@n���D 4@l��ҏ!?�/�~�@���4�ٿ>7���@@	��� 4@�U$G�!?���$�Z�@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@S��r�ٿ�HJ3�:�@��n4@�|,���!?+�~����@�;;:͞ٿ%�Ĕ�	�@'//DH4@٤���!?���F�@�;;:͞ٿ%�Ĕ�	�@'//DH4@٤���!?���F�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@H���>�ٿ�3�! �@�}3E� 4@��[�r�!?����gR�@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@�h�uc�ٿ�		�Ԫ�@���{��3@"m�H�!?+���@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@��U<ӫٿ�E����@+�Ԏ� 4@qG��{�!?�?��?��@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@�H��Q�ٿf�WN��@����4@��L�Z�!?g�b����@���C�ٿf���i�@��|}��3@ͧ����!?���\�@���C�ٿf���i�@��|}��3@ͧ����!?���\�@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@ ��ٿ϶ ����@��И 4@�Y|�!?2��K}��@�Π��ٿz�]����@`NM��3@��f�!?�"|#���@�Π��ٿz�]����@`NM��3@��f�!?�"|#���@�Π��ٿz�]����@`NM��3@��f�!?�"|#���@�Π��ٿz�]����@`NM��3@��f�!?�"|#���@�Π��ٿz�]����@`NM��3@��f�!?�"|#���@��šٿ�Yh�=�@H?�g 4@@\&q�!?���r�@����ٿ�ƌ�E�@W{I�4@��|i��!?�}FL���@����ٿ�ƌ�E�@W{I�4@��|i��!?�}FL���@����ٿ�ƌ�E�@W{I�4@��|i��!?�}FL���@#	G�ٿ�K�t�'�@�s��Z4@,il���!?0�6��@#	G�ٿ�K�t�'�@�s��Z4@,il���!?0�6��@��!���ٿ�X�K��@�	����3@��^��!?�A&�)�@��!���ٿ�X�K��@�	����3@��^��!?�A&�)�@��!���ٿ�X�K��@�	����3@��^��!?�A&�)�@��!���ٿ�X�K��@�	����3@��^��!?�A&�)�@d�A�ϕٿ�Z��9��@�y���3@�?z��!?�X��@d�A�ϕٿ�Z��9��@�y���3@�?z��!?�X��@2��b��ٿ�FBgС�@�ږ*��3@tֻvr�!?|4A��K�@2��b��ٿ�FBgС�@�ږ*��3@tֻvr�!?|4A��K�@2��b��ٿ�FBgС�@�ږ*��3@tֻvr�!?|4A��K�@2��b��ٿ�FBgС�@�ږ*��3@tֻvr�!?|4A��K�@��n�ߙٿ�+3��@ou��>�3@ӌ�v�!?��C�$�@��n�ߙٿ�+3��@ou��>�3@ӌ�v�!?��C�$�@��n�ߙٿ�+3��@ou��>�3@ӌ�v�!?��C�$�@��n�ߙٿ�+3��@ou��>�3@ӌ�v�!?��C�$�@&��Ğٿ����w��@����3@M��J��!?���vM�@�Xb��ٿ�z#����@𦗭��3@!��U�!?NΎq�:�@az�jC�ٿn��3`�@�XΨ��3@�u�ҙ�!?D�?�@az�jC�ٿn��3`�@�XΨ��3@�u�ҙ�!?D�?�@�T�}ٞٿ���7���@��T1% 4@R�?饏!?#$���@�T�}ٞٿ���7���@��T1% 4@R�?饏!?#$���@�T�}ٞٿ���7���@��T1% 4@R�?饏!?#$���@�T�}ٞٿ���7���@��T1% 4@R�?饏!?#$���@�T�}ٞٿ���7���@��T1% 4@R�?饏!?#$���@_�,ީٿt?����@��Q�y4@�"���!?���d��@��ٿX% ��p�@r�: 4@���fȏ!?	�d�C�@��ٿX% ��p�@r�: 4@���fȏ!?	�d�C�@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@oJQs�ٿ���� o�@�]��4@xRWs�!?E_a����@���/�ٿ�d���!�@	�%�4@渑�]�!?EHw����@޵ͩ9�ٿ9O�$J��@RV�
4@��զˏ!?�HO���@޵ͩ9�ٿ9O�$J��@RV�
4@��զˏ!?�HO���@޵ͩ9�ٿ9O�$J��@RV�
4@��զˏ!?�HO���@޵ͩ9�ٿ9O�$J��@RV�
4@��զˏ!?�HO���@޵ͩ9�ٿ9O�$J��@RV�
4@��զˏ!?�HO���@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@�QKO�ٿ����<�@�aY+4@�i���!?~^�Wb��@���#��ٿZ��\���@U�P�\ 4@iDn!?��3I�U�@���#��ٿZ��\���@U�P�\ 4@iDn!?��3I�U�@�e�F]�ٿ8��15#�@����4@��ˏ!?�x$��@xQA�ٿʓ��Q�@�5�(@�3@Z�B�
�!?�%� ��@xQA�ٿʓ��Q�@�5�(@�3@Z�B�
�!?�%� ��@xQA�ٿʓ��Q�@�5�(@�3@Z�B�
�!?�%� ��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@?���W�ٿ���3|��@ČI���3@��*R�!?�`<�!��@�&�b�ٿ��C+�@����34@Ε�٭�!?�������@�&�b�ٿ��C+�@����34@Ε�٭�!?�������@�&�b�ٿ��C+�@����34@Ε�٭�!?�������@:'��,�ٿ\��vJ�@��_a��3@X�l}Џ!?_F��@:'��,�ٿ\��vJ�@��_a��3@X�l}Џ!?_F��@:'��,�ٿ\��vJ�@��_a��3@X�l}Џ!?_F��@:'��,�ٿ\��vJ�@��_a��3@X�l}Џ!?_F��@:'��,�ٿ\��vJ�@��_a��3@X�l}Џ!?_F��@CaX���ٿ�~�#���@f����4@�Q~��!?I<�`�'�@CaX���ٿ�~�#���@f����4@�Q~��!?I<�`�'�@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@�p3*�ٿ���,P�@K2�� 4@�6P��!?��!}��@��㬚ٿ��T��@�B�YK�3@;�v��!?A��(x��@��㬚ٿ��T��@�B�YK�3@;�v��!?A��(x��@��㬚ٿ��T��@�B�YK�3@;�v��!?A��(x��@u�O���ٿ�� Z��@0=3ʎ 4@��R��!?3�_���@u�O���ٿ�� Z��@0=3ʎ 4@��R��!?3�_���@u�O���ٿ�� Z��@0=3ʎ 4@��R��!?3�_���@u�O���ٿ�� Z��@0=3ʎ 4@��R��!?3�_���@�$�~�ٿE�ч�<�@�%Z� 4@� m��!?����N�@�$�~�ٿE�ч�<�@�%Z� 4@� m��!?����N�@�$�~�ٿE�ч�<�@�%Z� 4@� m��!?����N�@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@A";${�ٿ,φ?	�@�*n� 4@Jr�q�!?Y�>���@2H���ٿoY*����@�k�� 4@�{W��!?KbJb�@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@��"��ٿy�h#*��@7h�, 4@q�mY��!?�ܠ1i��@�����ٿ�Õa��@:c]N� 4@Jely�!?4�c��b�@�����ٿ�Õa��@:c]N� 4@Jely�!?4�c��b�@�����ٿ�Õa��@:c]N� 4@Jely�!?4�c��b�@JFF4ءٿ�=�q�@�YX��4@��v�3�!?���.G�@JFF4ءٿ�=�q�@�YX��4@��v�3�!?���.G�@�v8�}�ٿ*���@����4@���tA�!?�kG�� �@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@?�O5�ٿ��A���@��o�k4@1�Z�!?��)^��@��D!N�ٿD����@�&�hS4@S
f�!?ڌ�����@��D!N�ٿD����@�&�hS4@S
f�!?ڌ�����@��D!N�ٿD����@�&�hS4@S
f�!?ڌ�����@��D!N�ٿD����@�&�hS4@S
f�!?ڌ�����@��D!N�ٿD����@�&�hS4@S
f�!?ڌ�����@ϡm�O�ٿD��]e�@]�0�� 4@>����!?� 96°�@�/��ٿS-F�VD�@��<l�3@�!�Ǐ!?�_�?]Y�@ }�k�ٿ#���N��@����! 4@X9�dm�!?�P���}�@ }�k�ٿ#���N��@����! 4@X9�dm�!?�P���}�@ }�k�ٿ#���N��@����! 4@X9�dm�!?�P���}�@ }�k�ٿ#���N��@����! 4@X9�dm�!?�P���}�@ }�k�ٿ#���N��@����! 4@X9�dm�!?�P���}�@u���ٿzj����@��7[t 4@�Ҝ��!?�Y�(�@u���ٿzj����@��7[t 4@�Ҝ��!?�Y�(�@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@|Q�խٿ1B+��@krt�{4@n���!?5�(uT��@���+-�ٿv����@��q�� 4@3=��ۏ!?��1>���@���+-�ٿv����@��q�� 4@3=��ۏ!?��1>���@���+-�ٿv����@��q�� 4@3=��ۏ!?��1>���@���?�ٿ�(���@���& 4@�u%�Ǐ!?�9�D�@���?�ٿ�(���@���& 4@�u%�Ǐ!?�9�D�@���?�ٿ�(���@���& 4@�u%�Ǐ!?�9�D�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@nB���ٿ�'���@��Ǫ� 4@���5Ϗ!?�y[�q�@Ϻ��ٿXn޸��@�9x�� 4@�ݰ8��!?��4eF�@Ϻ��ٿXn޸��@�9x�� 4@�ݰ8��!?��4eF�@Ϻ��ٿXn޸��@�9x�� 4@�ݰ8��!?��4eF�@Ϻ��ٿXn޸��@�9x�� 4@�ݰ8��!?��4eF�@Ϻ��ٿXn޸��@�9x�� 4@�ݰ8��!?��4eF�@[��s�ٿZ���H �@Nb 4@j��w	�!?NV�U;�@[��s�ٿZ���H �@Nb 4@j��w	�!?NV�U;�@��A괜ٿ�{2G��@-'h4@)R�!?́k��m�@��A괜ٿ�{2G��@-'h4@)R�!?́k��m�@��A괜ٿ�{2G��@-'h4@)R�!?́k��m�@�{�Y��ٿ�2�a��@���Z 4@�m�!��!?���?C�@�2�@��ٿ�"��/�@��[Q�4@��,��!?��7{�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@���ٿ;��bl�@v6�44@��w}��!?��i1�@d��!��ٿ���꜒�@�]��$4@�_��!?����R
�@d��!��ٿ���꜒�@�]��$4@�_��!?����R
�@d��!��ٿ���꜒�@�]��$4@�_��!?����R
�@d��!��ٿ���꜒�@�]��$4@�_��!?����R
�@d��!��ٿ���꜒�@�]��$4@�_��!?����R
�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@�:���ٿb��.O��@�*��4@~�#ŏ!?�0ث3�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@'�}L�ٿ�9��~��@�u\�x 4@� �ŏ!?X�/	C�@���I�ٿ+p�
5��@
�j�� 4@j%ŕ��!?��
�@���I�ٿ+p�
5��@
�j�� 4@j%ŕ��!?��
�@���I�ٿ+p�
5��@
�j�� 4@j%ŕ��!?��
�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@;WS��ٿ�ŴW���@�G�O4@`��&��!?�[�@�@��0���ٿg���:k�@����B4@�����!?��R;M!�@��;��ٿ����@K�Y-4@sPr���!?�**��@��;��ٿ����@K�Y-4@sPr���!?�**��@��;��ٿ����@K�Y-4@sPr���!?�**��@��;��ٿ����@K�Y-4@sPr���!?�**��@��;��ٿ����@K�Y-4@sPr���!?�**��@����ݭٿA�!X���@ ӊB��3@��)��!?f^�Ch/�@����ݭٿA�!X���@ ӊB��3@��)��!?f^�Ch/�@��L��ٿ�I,��@zQ�<O 4@'�����!?��͜y��@��L��ٿ�I,��@zQ�<O 4@'�����!?��͜y��@��L��ٿ�I,��@zQ�<O 4@'�����!?��͜y��@+�3lV�ٿ��Im���@��X�4@L�_��!?���h}�@¤交ٿ��h����@x�'*�4@W:\��!?�M�m�@¤交ٿ��h����@x�'*�4@W:\��!?�M�m�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@��
|�ٿ���g��@��@y�4@IG�ɏ!?��ߐ!�@+�$��ٿ#5�.��@bM !�4@��IRu�!?�K����@+�$��ٿ#5�.��@bM !�4@��IRu�!?�K����@���R�ٿ
Δ���@����4@JE���!?p��Iw��@���R�ٿ
Δ���@����4@JE���!?p��Iw��@���R�ٿ
Δ���@����4@JE���!?p��Iw��@���R�ٿ
Δ���@����4@JE���!?p��Iw��@���R�ٿ
Δ���@����4@JE���!?p��Iw��@���R�ٿ
Δ���@����4@JE���!?p��Iw��@�S[߯ٿx�Ud8C�@��N
4@�s�׏!?�/�T��@�?�=��ٿL�w����@3�����3@��%TЏ!?���7��@���W/�ٿh���{y�@�k���3@����!?�n�@��@���W/�ٿh���{y�@�k���3@����!?�n�@��@���W/�ٿh���{y�@�k���3@����!?�n�@��@�a�fl�ٿnߦ%���@ր/� 4@D3�{�!?���8��@�a�fl�ٿnߦ%���@ր/� 4@D3�{�!?���8��@�a�fl�ٿnߦ%���@ր/� 4@D3�{�!?���8��@�a�fl�ٿnߦ%���@ր/� 4@D3�{�!?���8��@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@����ٿ$S��@|���u�3@V�Q�g�!?��'�p�@�J�5�ٿA�ѭ��@�r�e 4@�&3B,�!?�N�w�@5�k��ٿ�p�|���@zZ� 4@��f#�!?@����@3x�	\�ٿ��K�Z�@~�u�_4@ӯI~E�!?N��M<�@[��z�ٿ�O�|�@@ª4@��F��!?ͶT���@[��z�ٿ�O�|�@@ª4@��F��!?ͶT���@[��z�ٿ�O�|�@@ª4@��F��!?ͶT���@Ў�{Q�ٿr��q��@A��p4@g�IV��!?�R?�R��@Ў�{Q�ٿr��q��@A��p4@g�IV��!?�R?�R��@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@c�t-�ٿ{�O�9��@�#W��4@�&�͏!?�B�U+�@�T�6�ٿ�g��b�@��(�C 4@l�,U�!?��t���@�Ȫ⇗ٿ�����<�@�j4@H/�x��!?�Oy��@�Ȫ⇗ٿ�����<�@�j4@H/�x��!?�Oy��@�Ȫ⇗ٿ�����<�@�j4@H/�x��!?�Oy��@�Ȫ⇗ٿ�����<�@�j4@H/�x��!?�Oy��@�Ȫ⇗ٿ�����<�@�j4@H/�x��!?�Oy��@ ўٿ�W��7/�@kr��-4@��ґ�!?5��+��@ ўٿ�W��7/�@kr��-4@��ґ�!?5��+��@ ўٿ�W��7/�@kr��-4@��ґ�!?5��+��@5�yۛٿ��=���@ N�zv4@5�ُ!?�O��H��@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@i�h]��ٿ�첎FT�@}�y\� 4@���ݏ!?n"�'�@R��J�ٿ�^qw�@��j�v 4@�E�9Џ!?iO;�6�@R��J�ٿ�^qw�@��j�v 4@�E�9Џ!?iO;�6�@R��J�ٿ�^qw�@��j�v 4@�E�9Џ!?iO;�6�@R��J�ٿ�^qw�@��j�v 4@�E�9Џ!?iO;�6�@R��J�ٿ�^qw�@��j�v 4@�E�9Џ!?iO;�6�@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@�*��1�ٿ��	�$�@Y�]a 4@ԃHK!?�-��@W�ٿ�S#P�@B�7���3@o܀Wo�!?g��~X�@W�ٿ�S#P�@B�7���3@o܀Wo�!?g��~X�@�9����ٿ�|��@]�@!�3j�3@�]�k�!?h�u��1�@�9����ٿ�|��@]�@!�3j�3@�]�k�!?h�u��1�@�Y�㡤ٿ�V�L~��@����3@v*(|��!?|�֦���@�Y�㡤ٿ�V�L~��@����3@v*(|��!?|�֦���@�;{��ٿן~���@����� 4@��%֫�!?���z�@�;{��ٿן~���@����� 4@��%֫�!?���z�@�;{��ٿן~���@����� 4@��%֫�!?���z�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@��`��ٿ�j�f���@�,f�4@�6���!?`U�CI�@PvT��ٿD�(�#�@A@�?� 4@���D��!?�A�o��@PvT��ٿD�(�#�@A@�?� 4@���D��!?�A�o��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@L�f	[�ٿ�uq��@���� 4@�Ɔo�!?��[v��@���Z�ٿa"{�ְ�@j���$�3@Ωj�f�!?7��4��@���Z�ٿa"{�ְ�@j���$�3@Ωj�f�!?7��4��@���Z�ٿa"{�ְ�@j���$�3@Ωj�f�!?7��4��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@tu|بٿ<y�"��@c����3@�@��ҏ!?\qVaP��@��.���ٿ
���	1�@�f���3@�7���!?^�x89��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@��ױ�ٿOy��L�@�w|�k�3@;�Vfɏ!?�x��g��@�I��ٿn��a���@D�4@��C��!?L�x�C�@��5�[�ٿ�����@��>�q 4@5D�H��!?^MS'��@�3�q�ٿ˨r�{�@�m����3@(�+D��!?�w��x�@�3�q�ٿ˨r�{�@�m����3@(�+D��!?�w��x�@�3�q�ٿ˨r�{�@�m����3@(�+D��!?�w��x�@�Z��)�ٿp�V���@ל�� 4@v���!?�p}o��@�Z��)�ٿp�V���@ל�� 4@v���!?�p}o��@%�,��ٿP��@���@�↹ �3@E*�+Џ!?_�2�k��@%�,��ٿP��@���@�↹ �3@E*�+Џ!?_�2�k��@%�,��ٿP��@���@�↹ �3@E*�+Џ!?_�2�k��@%�,��ٿP��@���@�↹ �3@E*�+Џ!?_�2�k��@%�,��ٿP��@���@�↹ �3@E*�+Џ!?_�2�k��@[�*�*�ٿ8� ~S��@�c���3@&1�͏!?�B�b�@[�*�*�ٿ8� ~S��@�c���3@&1�͏!?�B�b�@[�*�*�ٿ8� ~S��@�c���3@&1�͏!?�B�b�@Rmn��ٿR�ذ��@ܵmI4@Ԥq�؏!?��v��.�@Rmn��ٿR�ذ��@ܵmI4@Ԥq�؏!?��v��.�@Rmn��ٿR�ذ��@ܵmI4@Ԥq�؏!?��v��.�@Rmn��ٿR�ذ��@ܵmI4@Ԥq�؏!?��v��.�@�]�v�ٿ�`�'���@�j���3@��z��!?�+|����@�]�v�ٿ�`�'���@�j���3@��z��!?�+|����@�]�v�ٿ�`�'���@�j���3@��z��!?�+|����@�]�v�ٿ�`�'���@�j���3@��z��!?�+|����@�]�v�ٿ�`�'���@�j���3@��z��!?�+|����@�4���ٿ��7�@8���\4@�9��]�!?��΂�>�@0O�%�ٿ%eZ)E�@ �o�4@��D���!?6��.F�@0O�%�ٿ%eZ)E�@ �o�4@��D���!?6��.F�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@ox���ٿ&O衐��@/�AN4@�v!�Ǐ!?^M<�A�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@r8!c�ٿ�ԚU`��@]U�4�3@8�G�܏!?��e	!�@T�
�[�ٿ](�3Ҋ�@��Պ��3@�"O���!?*�&*�@T�
�[�ٿ](�3Ҋ�@��Պ��3@�"O���!?*�&*�@T�
�[�ٿ](�3Ҋ�@��Պ��3@�"O���!?*�&*�@T�
�[�ٿ](�3Ҋ�@��Պ��3@�"O���!?*�&*�@T�
�[�ٿ](�3Ҋ�@��Պ��3@�"O���!?*�&*�@��i�ٿ�*��y�@Z�m. 4@��U��!?���+'�@��i�ٿ�*��y�@Z�m. 4@��U��!?���+'�@��i�ٿ�*��y�@Z�m. 4@��U��!?���+'�@��_"�ٿq�����@�gJ�� 4@��R`̏!?7W�s��@��_"�ٿq�����@�gJ�� 4@��R`̏!?7W�s��@��_"�ٿq�����@�gJ�� 4@��R`̏!?7W�s��@��_"�ٿq�����@�gJ�� 4@��R`̏!?7W�s��@�r1�ҥٿR�<gA�@���]4@sB�ﳏ!?����R�@���ih�ٿ�������@����4@~�+n��!?��tc~�@���ih�ٿ�������@����4@~�+n��!?��tc~�@���$�ٿ�a�z2��@=�{J�4@|�ʜ��!?�>���@Xd���ٿ�m��Q�@�Y4@+�&ej�!?+^�r�@�S6�ٿ]nC��@�$��4@����!??/��@�S6�ٿ]nC��@�$��4@����!??/��@�S6�ٿ]nC��@�$��4@����!??/��@�S6�ٿ]nC��@�$��4@����!??/��@�-��ٿ#5��r�@%�Kh��3@�V"`��!?�x�Y�:�@�-��ٿ#5��r�@%�Kh��3@�V"`��!?�x�Y�:�@�-��ٿ#5��r�@%�Kh��3@�V"`��!?�x�Y�:�@�-��ٿ#5��r�@%�Kh��3@�V"`��!?�x�Y�:�@j5R��ٿ�C?ZX�@ǳ*��3@��	�!?����(&�@j5R��ٿ�C?ZX�@ǳ*��3@��	�!?����(&�@j5R��ٿ�C?ZX�@ǳ*��3@��	�!?����(&�@�i��ٿ\&�e�g�@40�04@�	}���!?M/6VX�@�#ZK�ٿ����N{�@V��� 4@Kŗ0�!?���_�@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@��L�ٿ�|�ز��@��:-{4@Yg�1/�!?m��L��@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@cXÛ�ٿ��n���@�m�i 4@�f$n��!?�O�M�%�@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�`���ٿ֐^]y��@ �E��3@_��я!?
�� ��@�5r�+�ٿe�D��@���� 4@��Y;܏!?c�`�K�@�5r�+�ٿe�D��@���� 4@��Y;܏!?c�`�K�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@X���ٿ�;�d���@p 1��3@�	{�ȏ!?~���}�@m7�ٿD9ↅ��@4���| 4@5��H�!?ЃI����@m7�ٿD9ↅ��@4���| 4@5��H�!?ЃI����@m7�ٿD9ↅ��@4���| 4@5��H�!?ЃI����@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@��*��ٿ�V�����@Um�ǳ�3@j���!?w�(�[��@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@(�ֱǛٿ�p�%�@?�Mo4@\}K쿏!?5���@'2
+�ٿp�pB��@��P 4@?s��ڏ!?�ݞ#9�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@M�ߙٿ�K<k���@�R0��4@��y��!?���V�M�@�c�7��ٿn�/���@8�<D4@
�A�!?
!hi�@�c�7��ٿn�/���@8�<D4@
�A�!?
!hi�@�c�7��ٿn�/���@8�<D4@
�A�!?
!hi�@�c�7��ٿn�/���@8�<D4@
�A�!?
!hi�@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@S!���ٿǟ�oF��@��^j��3@�yz.�!?�ůo��@}r�@ �ٿU�*����@1A�J4@��C�Ώ!?�Vo֚k�@}r�@ �ٿU�*����@1A�J4@��C�Ώ!?�Vo֚k�@z�U�E�ٿX�����@��X�4@ُ!?|~�d�@�F�ٿ�TC߅��@r'$ 4@�Z���!?�C��]�@�F�ٿ�TC߅��@r'$ 4@�Z���!?�C��]�@�F�ٿ�TC߅��@r'$ 4@�Z���!?�C��]�@�F�ٿ�TC߅��@r'$ 4@�Z���!?�C��]�@�F�ٿ�TC߅��@r'$ 4@�Z���!?�C��]�@}OҬ�ٿ���1�I�@ɇ��4@0x�̯�!?���ɬ�@}OҬ�ٿ���1�I�@ɇ��4@0x�̯�!?���ɬ�@}OҬ�ٿ���1�I�@ɇ��4@0x�̯�!?���ɬ�@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@��4��ٿ��_�A��@��y�d4@+A����!?LYn>��@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@���e�ٿq篧�d�@����4@t4��!?K>cQ)�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@ЊCP�ٿkP��su�@���p8 4@-�����!?�3>e?�@Y���حٿ:���jP�@���en�3@�n���!?F�����@Y���حٿ:���jP�@���en�3@�n���!?F�����@J&��*�ٿ��4آ��@Dߢ�� 4@i��d�!?
|��k9�@J&��*�ٿ��4آ��@Dߢ�� 4@i��d�!?
|��k9�@J&��*�ٿ��4آ��@Dߢ�� 4@i��d�!?
|��k9�@J&��*�ٿ��4آ��@Dߢ�� 4@i��d�!?
|��k9�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�\�K�ٿ5Sÿ2��@E��d4@.�r1^�!?���v�@�	丢ٿxXIT�y�@Mf՜�4@z����!?E`๨�@�	丢ٿxXIT�y�@Mf՜�4@z����!?E`๨�@�{7��ٿ��[n���@�B�e 4@0w$��!?�Y��@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@�-����ٿ
f9��:�@ý� 4@ʼ�r�!?����@gM���ٿp���Gl�@���	4@gɊ���!?6�����@P����ٿ�����c�@��5� 4@n)8��!??�����@P����ٿ�����c�@��5� 4@n)8��!??�����@P����ٿ�����c�@��5� 4@n)8��!??�����@*,NR��ٿP�q�A�@�=C�4@��g�[�!?�/�i���@*,NR��ٿP�q�A�@�=C�4@��g�[�!?�/�i���@>\~��ٿ�+��5�@A}� � 4@�
�C��!?َJ=<s�@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���[�ٿ�����o�@�ٝ� 4@}f�nӏ!?u4�F��@���U��ٿ8ƝZq�@vע���3@�@�檏!?l4P\��@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@؞��ʠٿ�����@쩇� 4@���W��!?�c9����@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@���"�ٿ��(�q��@�A��3@�ꎞ�!?V62g�"�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@Ą B�ٿne�/�.�@�Du%��3@��_��!?�ك"6�@��9�ٿ�r#�<�@�"k!h4@F�K�b�!?6��Q��@��9�ٿ�r#�<�@�"k!h4@F�K�b�!?6��Q��@�夬ٿ0��]!/�@��R4@����!?l�/F5�@_\��ٿb��[6U�@O�P�� 4@,���!?�K~(*��@��mκ�ٿ����y��@Tgk�3@���̏!?��(���@��mκ�ٿ����y��@Tgk�3@���̏!?��(���@SJ�i�ٿ�����@��� 4@�����!?@���.��@X����ٿKOf�@�AXe� 4@��Mo��!?�Pq�O�@X����ٿKOf�@�AXe� 4@��Mo��!?�Pq�O�@X����ٿKOf�@�AXe� 4@��Mo��!?�Pq�O�@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@M�?3�ٿ|0B���@�yh[��3@�-��!?�HZ��@̷5��ٿ$�q�@�J����3@OȨFŏ!?�ޘ]i��@̷5��ٿ$�q�@�J����3@OȨFŏ!?�ޘ]i��@̷5��ٿ$�q�@�J����3@OȨFŏ!?�ޘ]i��@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��߳�ٿ��T���@���l\ 4@�Y�ݏ!?D�N���@��?��ٿ`�LB��@�?Z���3@eFX���!?�ӺH��@��shr�ٿ�"]f�@�7��, 4@�[|�p�!?�Z�ߏ��@��shr�ٿ�"]f�@�7��, 4@�[|�p�!?�Z�ߏ��@��2���ٿ�Ϲ��@�L�O� 4@��Jz��!?C�im���@��2���ٿ�Ϲ��@�L�O� 4@��Jz��!?C�im���@��2���ٿ�Ϲ��@�L�O� 4@��Jz��!?C�im���@��2���ٿ�Ϲ��@�L�O� 4@��Jz��!?C�im���@a
���ٿى�%���@����4@
�����!?$�-���@a
���ٿى�%���@����4@
�����!?$�-���@�ZqW�ٿW>LR��@!�O� 4@0�}��!?pٍNt�@�ZqW�ٿW>LR��@!�O� 4@0�}��!?pٍNt�@�ZqW�ٿW>LR��@!�O� 4@0�}��!?pٍNt�@%ᓋ�ٿ����[�@�U,� 4@S�!��!?������@���ܔٿW�j}=��@���x��3@��a\��!?-\<J;�@���ܔٿW�j}=��@���x��3@��a\��!?-\<J;�@��؟�ٿ�� ��=�@(��r�3@��Yx��!?���Ǳ��@��؟�ٿ�� ��=�@(��r�3@��Yx��!?���Ǳ��@��؟�ٿ�� ��=�@(��r�3@��Yx��!?���Ǳ��@��؟�ٿ�� ��=�@(��r�3@��Yx��!?���Ǳ��@��؟�ٿ�� ��=�@(��r�3@��Yx��!?���Ǳ��@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@7D7�ٿ�0m:zM�@2�Z�3@�0�̏!?wb�
h�@׼4��ٿ nÆ�S�@�����3@r/9U��!?�"GU�@�(�F+�ٿ�þ�! �@���C��3@N���!?�@�����@�(�F+�ٿ�þ�! �@���C��3@N���!?�@�����@�(�F+�ٿ�þ�! �@���C��3@N���!?�@�����@�Ak���ٿ�q����@��H��3@�WvЏ!?���L��@}�i0��ٿ�R�����@�)�S�3@D0Ú�!?�T>m�@}�i0��ٿ�R�����@�)�S�3@D0Ú�!?�T>m�@}�i0��ٿ�R�����@�)�S�3@D0Ú�!?�T>m�@�yr�2�ٿr��j���@G��.��3@Sܒ���!?<��s��@�yr�2�ٿr��j���@G��.��3@Sܒ���!?<��s��@�yr�2�ٿr��j���@G��.��3@Sܒ���!?<��s��@��ߟ�ٿF�D+��@����3@*jK���!?ͯ��@��ߟ�ٿF�D+��@����3@*jK���!?ͯ��@l|�v�ٿ%	�4�(�@�[i� 4@�;�3��!?�A6H�x�@l|�v�ٿ%	�4�(�@�[i� 4@�;�3��!?�A6H�x�@l|�v�ٿ%	�4�(�@�[i� 4@�;�3��!?�A6H�x�@J(@0�ٿV,�s�G�@�v"��3@�J�ɏ!?�4�B��@��'~��ٿ����y�@�Խf�3@��̝��!?����2�@����L�ٿ{�\�u�@��8���3@9U>�ݏ!?�@3�E�@����L�ٿ{�\�u�@��8���3@9U>�ݏ!?�@3�E�@����ٿ�R���@6�oMH 4@�?m��!?;�r��F�@����ٿ�R���@6�oMH 4@�?m��!?;�r��F�@����ٿ�R���@6�oMH 4@�?m��!?;�r��F�@����ٿ�R���@6�oMH 4@�?m��!?;�r��F�@�~uڬٿ^���һ�@��*�4@1�����!?�#�V��@�~uڬٿ^���һ�@��*�4@1�����!?�#�V��@�~uڬٿ^���һ�@��*�4@1�����!?�#�V��@�P1@ԫٿO����@A�Fe 4@�����!?�S���E�@�P1@ԫٿO����@A�Fe 4@�����!?�S���E�@N\����ٿ�����@�E�c�4@�����!?������@N\����ٿ�����@�E�c�4@�����!?������@N\����ٿ�����@�E�c�4@�����!?������@N\����ٿ�����@�E�c�4@�����!?������@N\����ٿ�����@�E�c�4@�����!?������@N\����ٿ�����@�E�c�4@�����!?������@�
)q��ٿ����o�@�\ �A 4@�ۏ��!?X��i���@�
)q��ٿ����o�@�\ �A 4@�ۏ��!?X��i���@�
)q��ٿ����o�@�\ �A 4@�ۏ��!?X��i���@�
)q��ٿ����o�@�\ �A 4@�ۏ��!?X��i���@���@�ٿ,lˋ�,�@K-C4@��#я!?�������@���@�ٿ,lˋ�,�@K-C4@��#я!?�������@n�Wޚٿ'ܵ����@�A��`4@�yS��!?8{t�.;�@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@�9�i�ٿ��k�d�@�أ'�4@�$q홏!?�����@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@p  !��ٿ����;l�@����z 4@	��p��!?fk:F��@��n-�ٿ@B4��@q�a� 4@!+�+͏!?!���@��n-�ٿ@B4��@q�a� 4@!+�+͏!?!���@��n-�ٿ@B4��@q�a� 4@!+�+͏!?!���@��n-�ٿ@B4��@q�a� 4@!+�+͏!?!���@��n-�ٿ@B4��@q�a� 4@!+�+͏!?!���@�C�ݾ�ٿT�g���@P��p�4@h�\�!?��jQ��@���h�ٿ��]d���@'K���4@[��AV�!?=T��@���h�ٿ��]d���@'K���4@[��AV�!?=T��@��#`�ٿ�@�6��@�t*�4@K��"��!?Vs.���@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@d!^�ٿ8e�BP/�@�\ �4@�VK��!?7oq�4�@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@��.�s�ٿ�E�X�_�@GY�g�4@�-�Ǐ!?���g��@�O����ٿo(<4���@&P>`4@Q��3��!?�?ZX���@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@������ٿ�n��u�@����4@��"��!?�ܕW��@
�q��ٿ�cKz���@7�7}44@��G��!?��?"��@q3�5�ٿ3:��'g�@���dg4@�RY�v�!?-~�����@�h�#�ٿ,B���I�@i�w�P�3@
g�H.�!?����$�@W����ٿӠ!9��@:�Y[��3@q�^�%�!?)n��Z�@W����ٿӠ!9��@:�Y[��3@q�^�%�!?)n��Z�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@��B�R�ٿ��{��@΂c�O 4@��A�`�!?�oMY�@k�x��ٿ�s���@�ܥ�0�3@ޜ����!?^#k���@k�x��ٿ�s���@�ܥ�0�3@ޜ����!?^#k���@�f����ٿ֕O���@�{÷�3@�r+h�!?n��O�@�f����ٿ֕O���@�{÷�3@�r+h�!?n��O�@�f����ٿ֕O���@�{÷�3@�r+h�!?n��O�@�f����ٿ֕O���@�{÷�3@�r+h�!?n��O�@�f����ٿ֕O���@�{÷�3@�r+h�!?n��O�@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@��q�ٿ������@���5 4@LN�r�!?�0͑���@AQU��ٿ�XFLQ��@k����3@�P��!?��ͅ��@�BC�̮ٿW�)���@NHU�3@����!?�c�Xz�@�BC�̮ٿW�)���@NHU�3@����!?�c�Xz�@�BC�̮ٿW�)���@NHU�3@����!?�c�Xz�@�BC�̮ٿW�)���@NHU�3@����!?�c�Xz�@:���ٿ��U.��@���S 4@��?��!?�q�[���@������ٿ��p�8��@Nױ�1�3@�-����!?x��)V �@������ٿ��p�8��@Nױ�1�3@�-����!?x��)V �@������ٿ��p�8��@Nױ�1�3@�-����!?x��)V �@������ٿ��p�8��@Nױ�1�3@�-����!?x��)V �@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@��D�ٿ6�qd��@�+YL) 4@��ԏ!?�S�G�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@�Ad�ٿ�Bw;���@g!�� 4@^�^��!?[ G��A�@��U�ʟٿ������@.�I�f 4@�S���!?<�#r��@��U�ʟٿ������@.�I�f 4@�S���!?<�#r��@��U�ʟٿ������@.�I�f 4@�S���!?<�#r��@��U�ʟٿ������@.�I�f 4@�S���!?<�#r��@��U�ʟٿ������@.�I�f 4@�S���!?<�#r��@�-�ĝٿ(����@�Jd��3@J۽$�!?�`�$A@�@�-�ĝٿ(����@�Jd��3@J۽$�!?�`�$A@�@�-�ĝٿ(����@�Jd��3@J۽$�!?�`�$A@�@�-�ĝٿ(����@�Jd��3@J۽$�!?�`�$A@�@�-�ĝٿ(����@�Jd��3@J۽$�!?�`�$A@�@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@.��͛ٿO�=��
�@�U�R 4@���!?O��l��@�Jad�ٿ�����@W����3@�]&���!?�g�0��@�Jad�ٿ�����@W����3@�]&���!?�g�0��@�Jad�ٿ�����@W����3@�]&���!?�g�0��@�Jad�ٿ�����@W����3@�]&���!?�g�0��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@{Q_�ٿ��_X���@(~m44@*l[�!?5.�N��@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@��w�;�ٿ�
��>�@���a 4@V�ߏ!?�ܾg�@���ͮٿ?ؚ���@�)�[] 4@0o`|��!?�]���@���ͮٿ?ؚ���@�)�[] 4@0o`|��!?�]���@;�v�ٿl����@Oţ�S4@�8"��!?�V+��@;�v�ٿl����@Oţ�S4@�8"��!?�V+��@��8+��ٿ7�6�1�@��3�~4@u����!?��?!7�@���*��ٿ&݊�P�@����4@���>1�!?-�����@���*��ٿ&݊�P�@����4@���>1�!?-�����@���*��ٿ&݊�P�@����4@���>1�!?-�����@���*��ٿ&݊�P�@����4@���>1�!?-�����@���*��ٿ&݊�P�@����4@���>1�!?-�����@��̴=�ٿG]���@���4@c!��7�!?��EH=�@��̴=�ٿG]���@���4@c!��7�!?��EH=�@��̴=�ٿG]���@���4@c!��7�!?��EH=�@��̴=�ٿG]���@���4@c!��7�!?��EH=�@��̴=�ٿG]���@���4@c!��7�!?��EH=�@.l���ٿN�v���@(�| Z 4@A��"�!?�zw|d�@.l���ٿN�v���@(�| Z 4@A��"�!?�zw|d�@	��£ٿ���G���@�1:e4@���ѝ�!?�ޥ9.a�@	��£ٿ���G���@�1:e4@���ѝ�!?�ޥ9.a�@	��£ٿ���G���@�1:e4@���ѝ�!?�ޥ9.a�@	��£ٿ���G���@�1:e4@���ѝ�!?�ޥ9.a�@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@8�+�ٿ&��ƍ��@:��Z�4@�Ӡ��!?�a����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@H�{�H�ٿy��M�@mB%h4@"gxʏ!?�o`����@J��Ǜٿ'�:E�@p���]4@�<�j��!?���@J��Ǜٿ'�:E�@p���]4@�<�j��!?���@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@Ҳ�Ǎ�ٿ��;=��@Y�)�4@M�z�_�!?I��eW�@�%�ٿ�Qs���@P�+�d4@09��P�!?M�D���@Ac�!�ٿ2_ty��@��d4@X�A֏!?��6��@Ac�!�ٿ2_ty��@��d4@X�A֏!?��6��@Ac�!�ٿ2_ty��@��d4@X�A֏!?��6��@Ac�!�ٿ2_ty��@��d4@X�A֏!?��6��@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@N��Z"�ٿ�B��@5>Y� 4@�@��!?b9�ـ�@��S	ўٿ'�JvS��@���� 4@@ Ǐ!?�|U����@��S	ўٿ'�JvS��@���� 4@@ Ǐ!?�|U����@Ve�]�ٿ��.���@#�����3@P̷�!?�\��>��@Ve�]�ٿ��.���@#�����3@P̷�!?�\��>��@Ae\�ٿ���R���@���v! 4@�~?C�!?f>�T��@Ae\�ٿ���R���@���v! 4@�~?C�!?f>�T��@Ae\�ٿ���R���@���v! 4@�~?C�!?f>�T��@5ຖ-�ٿ2������@�O9w�4@�	h���!?���C��@5ຖ-�ٿ2������@�O9w�4@�	h���!?���C��@5ຖ-�ٿ2������@�O9w�4@�	h���!?���C��@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@�u���ٿ(&K���@+te�4@��'ݹ�!?>g��4�@6�R�z�ٿ��*qE�@T�i�4@������!?��."��@6�R�z�ٿ��*qE�@T�i�4@������!?��."��@6�R�z�ٿ��*qE�@T�i�4@������!?��."��@6�R�z�ٿ��*qE�@T�i�4@������!?��."��@6�R�z�ٿ��*qE�@T�i�4@������!?��."��@ I�ٿRf�k�@�����4@p@DR}�!?+��l�@�2��ٿ4�)���@�y��4@����ҏ!?h/�2��@�2��ٿ4�)���@�y��4@����ҏ!?h/�2��@�2��ٿ4�)���@�y��4@����ҏ!?h/�2��@�2��ٿ4�)���@�y��4@����ҏ!?h/�2��@B����ٿca��@�`ԝS4@߾k�!?��U��L�@B����ٿca��@�`ԝS4@߾k�!?��U��L�@B����ٿca��@�`ԝS4@߾k�!?��U��L�@B����ٿca��@�`ԝS4@߾k�!?��U��L�@�FqӍ�ٿ�T���@��q�� 4@�,O;؏!?v�&X��@�FqӍ�ٿ�T���@��q�� 4@�,O;؏!?v�&X��@�FqӍ�ٿ�T���@��q�� 4@�,O;؏!?v�&X��@�FqӍ�ٿ�T���@��q�� 4@�,O;؏!?v�&X��@�F�]�ٿgS�>�D�@"֑]u4@�����!?mu�����@AEձӱٿ�A�T�@J+� 4@0F��T�!?g��PC�@AEձӱٿ�A�T�@J+� 4@0F��T�!?g��PC�@AEձӱٿ�A�T�@J+� 4@0F��T�!?g��PC�@AEձӱٿ�A�T�@J+� 4@0F��T�!?g��PC�@AEձӱٿ�A�T�@J+� 4@0F��T�!?g��PC�@�&�(��ٿ��Č\�@���4@7��p�!?#����@�&�(��ٿ��Č\�@���4@7��p�!?#����@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@4�D���ٿ���ۛ��@���4@dWRz�!?��1�9�@����
�ٿ�}3��@���B4@~��!��!?��Z��@����
�ٿ�}3��@���B4@~��!��!?��Z��@����
�ٿ�}3��@���B4@~��!��!?��Z��@+��ãٿ�P���@���[4@[#�ߏ!?���`Q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@���'q�ٿ�m��A��@�� 4@�T�w��!?��i�q�@f���3�ٿ���R��@���4@��&��!?G�*ܧ��@f���3�ٿ���R��@���4@��&��!?G�*ܧ��@f���3�ٿ���R��@���4@��&��!?G�*ܧ��@f���3�ٿ���R��@���4@��&��!?G�*ܧ��@�$/䧕ٿa5L<Z��@�9�� 4@g+��R�!?xɘJ�H�@�$/䧕ٿa5L<Z��@�9�� 4@g+��R�!?xɘJ�H�@�$/䧕ٿa5L<Z��@�9�� 4@g+��R�!?xɘJ�H�@�$/䧕ٿa5L<Z��@�9�� 4@g+��R�!?xɘJ�H�@�X��>�ٿ<����@�F�_ 4@�󵪂�!?aS��@�X��>�ٿ<����@�F�_ 4@�󵪂�!?aS��@�X��>�ٿ<����@�F�_ 4@�󵪂�!?aS��@	T��ٿ�h(���@��vg 4@��st��!?"���@	T��ٿ�h(���@��vg 4@��st��!?"���@	T��ٿ�h(���@��vg 4@��st��!?"���@6?�~�ٿ2�
�k��@+_45L 4@�7F�!?���h1�@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��=��ٿ��҄�@�Q(@ 4@â�a��!?��%��@��4�?�ٿ�FN����@�y�,a4@Y��!?�%����@��4�?�ٿ�FN����@�y�,a4@Y��!?�%����@�A[���ٿQV�O�@��!4��3@c@���!?6v,k-�@�A[���ٿQV�O�@��!4��3@c@���!?6v,k-�@�A[���ٿQV�O�@��!4��3@c@���!?6v,k-�@�A[���ٿQV�O�@��!4��3@c@���!?6v,k-�@�A[���ٿQV�O�@��!4��3@c@���!?6v,k-�@��/��ٿ����0�@SZ���3@�r��w�!?U����V�@
_V�ٿ9�pv��@�޴�a 4@���k�!?�E�Ս��@Ӓ�1�ٿ������@����3@zsb\�!?l7�`�@Ӓ�1�ٿ������@����3@zsb\�!?l7�`�@�Ov��ٿ��^H}��@P��\��3@��s��!?��ꌄ��@#\V�ٿQ�u�QQ�@���� 4@�$ɇ,�!?n%��4��@#\V�ٿQ�u�QQ�@���� 4@�$ɇ,�!?n%��4��@#\V�ٿQ�u�QQ�@���� 4@�$ɇ,�!?n%��4��@#\V�ٿQ�u�QQ�@���� 4@�$ɇ,�!?n%��4��@#\V�ٿQ�u�QQ�@���� 4@�$ɇ,�!?n%��4��@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@� YW�ٿ(����@y|�� 4@�#:VH�!?�!�����@do��ٿ �&u4��@��t�/�3@uIv���!?��f<�@do��ٿ �&u4��@��t�/�3@uIv���!?��f<�@do��ٿ �&u4��@��t�/�3@uIv���!?��f<�@do��ٿ �&u4��@��t�/�3@uIv���!?��f<�@pu?�P�ٿ��	G��@�c[�7 4@9B.瓏!?�����3�@�lOd,�ٿ��Tp���@�6W]4@LFg�ˏ!?/��{��@�lOd,�ٿ��Tp���@�6W]4@LFg�ˏ!?/��{��@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�ɕ�ٿ�)���@��˲E4@�tT��!?�cʹ���@�Л���ٿ�/��D��@x��J 4@�ERl�!?X"����@��ͨٿ-'Mx���@��hb4@L��Џ!?�31)��@٘��ˤٿ;F�z�@4���4@M4�ɏ!?��J���@���y�ٿ���O(�@���� 4@�h@�$�!?��pםX�@���y�ٿ���O(�@���� 4@�h@�$�!?��pםX�@���y�ٿ���O(�@���� 4@�h@�$�!?��pםX�@���y�ٿ���O(�@���� 4@�h@�$�!?��pםX�@��n.�ٿT�F6���@��1�4@Q�\ �!?���9�@��n.�ٿT�F6���@��1�4@Q�\ �!?���9�@��n.�ٿT�F6���@��1�4@Q�\ �!?���9�@��n.�ٿT�F6���@��1�4@Q�\ �!?���9�@��n.�ٿT�F6���@��1�4@Q�\ �!?���9�@��ٿ_�����@
�}}4@���Ǐ!?.~�	Q��@��ٿ_�����@
�}}4@���Ǐ!?.~�	Q��@��ٿ_�����@
�}}4@���Ǐ!?.~�	Q��@�w5[��ٿ�.v7�o�@�Z5J 4@nȮk��!?����&�@�w5[��ٿ�.v7�o�@�Z5J 4@nȮk��!?����&�@�`�H-�ٿ�3EJ��@}r�% 4@`��"~�!?f����@�`�H-�ٿ�3EJ��@}r�% 4@`��"~�!?f����@���r��ٿ(1��ԯ�@�ߕ�l 4@�[tj�!?	� ���@���r��ٿ(1��ԯ�@�ߕ�l 4@�[tj�!?	� ���@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@�Z7���ٿ�V
#��@@@Q8=4@��8��!?$0
s��@��J��ٿS�W_�@׉�%4@p�%:�!?��T�n�@���љ�ٿ��bK�@=�1@4@��<ʏ!?�agҁ��@���љ�ٿ��bK�@=�1@4@��<ʏ!?�agҁ��@���љ�ٿ��bK�@=�1@4@��<ʏ!?�agҁ��@���љ�ٿ��bK�@=�1@4@��<ʏ!?�agҁ��@���љ�ٿ��bK�@=�1@4@��<ʏ!?�agҁ��@A_���ٿ��\%6�@�|)���3@+�OLҏ!?�l�7˳�@A_���ٿ��\%6�@�|)���3@+�OLҏ!?�l�7˳�@A_���ٿ��\%6�@�|)���3@+�OLҏ!?�l�7˳�@A_���ٿ��\%6�@�|)���3@+�OLҏ!?�l�7˳�@<rLf�ٿV��0��@���i�4@jV���!?j������@<rLf�ٿV��0��@���i�4@jV���!?j������@<rLf�ٿV��0��@���i�4@jV���!?j������@A�L��ٿǫ��{��@A�[��3@�C�Y��!?�����@A�L��ٿǫ��{��@A�[��3@�C�Y��!?�����@A�L��ٿǫ��{��@A�[��3@�C�Y��!?�����@A�L��ٿǫ��{��@A�[��3@�C�Y��!?�����@��:�0�ٿ�ߚ���@���� 4@Q	�q�!?8�>���@��:�0�ٿ�ߚ���@���� 4@Q	�q�!?8�>���@��:�0�ٿ�ߚ���@���� 4@Q	�q�!?8�>���@,��ٿ�F���<�@���H�4@p.���!?���I�d�@,��ٿ�F���<�@���H�4@p.���!?���I�d�@,��ٿ�F���<�@���H�4@p.���!?���I�d�@,��ٿ�F���<�@���H�4@p.���!?���I�d�@,��ٿ�F���<�@���H�4@p.���!?���I�d�@�6��ٿ��s���@��6�w4@�/Di��!?�|��E��@�6��ٿ��s���@��6�w4@�/Di��!?�|��E��@�6��ٿ��s���@��6�w4@�/Di��!?�|��E��@�6��ٿ��s���@��6�w4@�/Di��!?�|��E��@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@��"��ٿ֫o�e��@�(>�|4@�֬Ҡ�!?y�����@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@t�W|P�ٿH�/́f�@�x{�8�3@�ܲy��!?���@��@�w�W�ٿp�ɽ���@��n�@�3@��2�u�!?9�ʨ��@�w�W�ٿp�ɽ���@��n�@�3@��2�u�!?9�ʨ��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��k;��ٿZ~�xf�@}<�4@�t�H��!?t ']��@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@��S�}�ٿ�.��@�� 4@��Q
̏!?3c�d�@���.r�ٿ��4���@��x1� 4@@ ��ԏ!?�;�UƓ�@���.r�ٿ��4���@��x1� 4@@ ��ԏ!?�;�UƓ�@���.r�ٿ��4���@��x1� 4@@ ��ԏ!?�;�UƓ�@���.r�ٿ��4���@��x1� 4@@ ��ԏ!?�;�UƓ�@���.r�ٿ��4���@��x1� 4@@ ��ԏ!?�;�UƓ�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@j>�#�ٿs�/q���@�u���3@�B�"��!?�'��;H�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@��y��ٿ��`�B�@�gX!4@��^#p�!?6�Ñ�D�@���*��ٿ�X��kv�@w��W 4@�	gڔ�!?e�@����@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Z��ٿ�1�q���@Ҥt"�4@_��^֏!?C���)��@��Ҩi�ٿ����@2�� 4@�n��!?,�&L�@��Ҩi�ٿ����@2�� 4@�n��!?,�&L�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@KK�`f�ٿ�Yn����@4��~<�3@5��U��!?q;r�<�@�#��_�ٿ/��DG�@����3@8��?��!?�b9�A�@��Ñ�ٿ�]NV���@X��;s 4@�J[���!?��+M��@��Ñ�ٿ�]NV���@X��;s 4@�J[���!?��+M��@��Ñ�ٿ�]NV���@X��;s 4@�J[���!?��+M��@��Ñ�ٿ�]NV���@X��;s 4@�J[���!?��+M��@��R��ٿe
IN��@˵��
4@u�D8��!?t�3o��@��R��ٿe
IN��@˵��
4@u�D8��!?t�3o��@��R��ٿe
IN��@˵��
4@u�D8��!?t�3o��@��R��ٿe
IN��@˵��
4@u�D8��!?t�3o��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@���Üٿ�g�w��@���n�3@��1���!?��/( ��@<2���ٿ"�;@�@��tL� 4@����Q�!?��QF��@<2���ٿ"�;@�@��tL� 4@����Q�!?��QF��@<2���ٿ"�;@�@��tL� 4@����Q�!?��QF��@��6���ٿZJT|��@R�h.4@NtxJ�!?�V����@��6���ٿZJT|��@R�h.4@NtxJ�!?�V����@�����ٿ�[RR{��@|b�R�3@)-��P�!?��+�C��@����_�ٿ�g��j��@7�-c�3@5[�ξ�!?H(����@����_�ٿ�g��j��@7�-c�3@5[�ξ�!?H(����@����_�ٿ�g��j��@7�-c�3@5[�ξ�!?H(����@����_�ٿ�g��j��@7�-c�3@5[�ξ�!?H(����@L�D�G�ٿkP�:��@��U��3@�V8�!?��m(��@L�D�G�ٿkP�:��@��U��3@�V8�!?��m(��@L�D�G�ٿkP�:��@��U��3@�V8�!?��m(��@-�BQ;�ٿ<������@��:�4@�#t�!?����C��@�Fg�ܦٿ7���l�@F��4@�=7�d�!?���E�@�Fg�ܦٿ7���l�@F��4@�=7�d�!?���E�@�Fg�ܦٿ7���l�@F��4@�=7�d�!?���E�@h��]�ٿ���kK9�@O�)q`�3@����!?�d��@h��]�ٿ���kK9�@O�)q`�3@����!?�d��@h��]�ٿ���kK9�@O�)q`�3@����!?�d��@����|�ٿD�����@lЍ.�3@�$��X�!?��Z`��@����|�ٿD�����@lЍ.�3@�$��X�!?��Z`��@c�)6�ٿz3.�`�@ef���3@�����!?�؂Վb�@�'���ٿTz�8��@�����3@M#G\o�!?{<j
0�@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@�I$��ٿ?�W��w�@����� 4@-�穏!?c�����@��mcM�ٿ��ԁ\�@�6�ZZ4@�C:x�!?��=���@*3�z�ٿ���E)�@����9 4@�FtP��!?�ř�C�@*3�z�ٿ���E)�@����9 4@�FtP��!?�ř�C�@�U56ܢٿ�|�A�o�@d�h���3@�Ǫ�!?�~�fI��@�U56ܢٿ�|�A�o�@d�h���3@�Ǫ�!?�~�fI��@�U56ܢٿ�|�A�o�@d�h���3@�Ǫ�!?�~�fI��@�U56ܢٿ�|�A�o�@d�h���3@�Ǫ�!?�~�fI��@�U56ܢٿ�|�A�o�@d�h���3@�Ǫ�!?�~�fI��@GI>��ٿ��E_-��@w ��4@=F3:��!?�AVƶ�@GI>��ٿ��E_-��@w ��4@=F3:��!?�AVƶ�@�2I���ٿ�;1�D��@l�)��3@�MhPُ!?��Ȋ%�@�2I���ٿ�;1�D��@l�)��3@�MhPُ!?��Ȋ%�@�2I���ٿ�;1�D��@l�)��3@�MhPُ!?��Ȋ%�@�2I���ٿ�;1�D��@l�)��3@�MhPُ!?��Ȋ%�@Q;�=Şٿ�J�g8�@o��� 4@�%��!?�Y�U�3�@Q;�=Şٿ�J�g8�@o��� 4@�%��!?�Y�U�3�@M� �^�ٿjdY)���@�&����3@2/�L��!?0R���|�@M� �^�ٿjdY)���@�&����3@2/�L��!?0R���|�@M� �^�ٿjdY)���@�&����3@2/�L��!?0R���|�@M� �^�ٿjdY)���@�&����3@2/�L��!?0R���|�@֕�[�ٿZoO����@l_;��4@^�!��!?|�����@֕�[�ٿZoO����@l_;��4@^�!��!?|�����@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@B,���ٿ�H�,ĸ�@���g4@��Õ~�!?�)S'A��@-!��H�ٿR�Zx��@�^��4@�h�Տ!?"O%M��@-!��H�ٿR�Zx��@�^��4@�h�Տ!?"O%M��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@C���`�ٿ1)̈M�@�h؏4@�u-Ï!?M�<DC��@_D�ٿ[-Ÿ�@�/~��3@ms�'w�!?X����@_D�ٿ[-Ÿ�@�/~��3@ms�'w�!?X����@_D�ٿ[-Ÿ�@�/~��3@ms�'w�!?X����@�'?���ٿD���P�@�!�g4@H�S�+�!?�4�`��@#��1�ٿ�K+E*��@
�~��4@d8H�!?0��))�@#��1�ٿ�K+E*��@
�~��4@d8H�!?0��))�@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@q��'�ٿBx���@�A7B 4@�%��w�!?w�ҳK��@8���V�ٿ���:.��@IS��3@�sIf��!?U��ߦ�@8���V�ٿ���:.��@IS��3@�sIf��!?U��ߦ�@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@7��[֛ٿ�$55���@3L���4@�P~稏!?1B1 ��@�>�[��ٿ�wp���@�)�L[4@
$\���!?7�x�<�@i�67v�ٿ����@�ɼ@d4@�Íÿ�!?-�3T.M�@K�ZI�ٿ�G�m�S�@2П�� 4@"����!?�z��ڛ�@K�ZI�ٿ�G�m�S�@2П�� 4@"����!?�z��ڛ�@	��C��ٿz�Q�.��@1��uf4@������!?J����@	��C��ٿz�Q�.��@1��uf4@������!?J����@	��C��ٿz�Q�.��@1��uf4@������!?J����@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�� �G�ٿ`ᡦ��@�+	c4@�3��!?��G{�@�pk���ٿ������@���~4@\�r���!?@�pԔ�@�pk���ٿ������@���~4@\�r���!?@�pԔ�@�pk���ٿ������@���~4@\�r���!?@�pԔ�@�pk���ٿ������@���~4@\�r���!?@�pԔ�@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�ܜa�ٿZ�?�&'�@$1�4@� ���!?� MY��@�>��ٿ��W�@R�ɑ�4@�\)�!?�3�q���@�.o-�ٿ؎����@��.�4@@d�&��!?���l:��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@�Tj�ٿ�nd���@]��4@�:�Կ�!?�v~œ��@����ٿˊ�F�@�m*�4@���£�!?�؝�@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�l�ٿX3 � ��@f�M�4@��7��!?Oբ���@�r��x�ٿɥr��H�@u y�(4@�+��ߏ!?�>�����@�r��x�ٿɥr��H�@u y�(4@�+��ߏ!?�>�����@�r��x�ٿɥr��H�@u y�(4@�+��ߏ!?�>�����@T<��ٿ���_��@P2q4@r�(J��!?̼<����@,w����ٿ���@1 ��,�3@nЅϏ!?�p���R�@,w����ٿ���@1 ��,�3@nЅϏ!?�p���R�@,w����ٿ���@1 ��,�3@nЅϏ!?�p���R�@,w����ٿ���@1 ��,�3@nЅϏ!?�p���R�@���s��ٿ��0���@�.��� 4@���~��!?�����D�@���s��ٿ��0���@�.��� 4@���~��!?�����D�@7��"ڤٿ�oB��7�@.#
u4@ye-&��!?�^��&�@7��"ڤٿ�oB��7�@.#
u4@ye-&��!?�^��&�@7��"ڤٿ�oB��7�@.#
u4@ye-&��!?�^��&�@7��"ڤٿ�oB��7�@.#
u4@ye-&��!?�^��&�@�����ٿ<]ŧ#��@2!���4@F�a�!?��L@��@�����ٿ<]ŧ#��@2!���4@F�a�!?��L@��@�����ٿ<]ŧ#��@2!���4@F�a�!?��L@��@b��}�ٿ/4ռ	{�@�M�L	4@�yN��!?��̒0�@b��}�ٿ/4ռ	{�@�M�L	4@�yN��!?��̒0�@��c}�ٿc�F�\�@�F*�!4@�!rC��!?	��~AU�@K��<�ٿ�ѥ��@���4@Z�,��!??�Vs��@�'�6�ٿ�)��7�@>"֓� 4@�����!?��i\�@"7	��ٿ�n���m�@�0(4@�Ż~��!?�������@"7	��ٿ�n���m�@�0(4@�Ż~��!?�������@"7	��ٿ�n���m�@�0(4@�Ż~��!?�������@;�W���ٿ�^��h�@Vۣ� 4@ ����!?�7FY�@;�W���ٿ�^��h�@Vۣ� 4@ ����!?�7FY�@LA�8��ٿ��*?�I�@<�\Ѯ 4@H��6��!?�O�H���@���ٿ�0W[p?�@v@�P 4@b��p��!?ɪ��^�@���ٿ�0W[p?�@v@�P 4@b��p��!?ɪ��^�@���ٿ�0W[p?�@v@�P 4@b��p��!?ɪ��^�@���ٿ�0W[p?�@v@�P 4@b��p��!?ɪ��^�@���ٿ�0W[p?�@v@�P 4@b��p��!?ɪ��^�@���5D�ٿ ��i�@�.��| 4@s��!?��R� �@���5D�ٿ ��i�@�.��| 4@s��!?��R� �@���5D�ٿ ��i�@�.��| 4@s��!?��R� �@���5D�ٿ ��i�@�.��| 4@s��!?��R� �@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@W��(W�ٿ��*�D�@���?4@�^�t�!?�}�R�@��LZ�ٿ��#�@�ڱ$ 4@L�B ��!?jrA�8u�@��2�ٿw������@H�Vݹ 4@�JW�!?���a��@��2�ٿw������@H�Vݹ 4@�JW�!?���a��@��2�ٿw������@H�Vݹ 4@�JW�!?���a��@�0�ٿn2���@��Oo�3@��~�!?��S}�e�@�0�ٿn2���@��Oo�3@��~�!?��S}�e�@�0�ٿn2���@��Oo�3@��~�!?��S}�e�@�0�ٿn2���@��Oo�3@��~�!?��S}�e�@Wav	�ٿ�����6�@�̃�� 4@�=��!?�P��w�@Wav	�ٿ�����6�@�̃�� 4@�=��!?�P��w�@Wav	�ٿ�����6�@�̃�� 4@�=��!?�P��w�@Wav	�ٿ�����6�@�̃�� 4@�=��!?�P��w�@Wav	�ٿ�����6�@�̃�� 4@�=��!?�P��w�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@�ԐU4�ٿ�k��@8�4@(����!?M�t��4�@������ٿ�S�O���@�:�+4@4�S�ߏ!?+��W��@������ٿ�S�O���@�:�+4@4�S�ߏ!?+��W��@������ٿ�S�O���@�:�+4@4�S�ߏ!?+��W��@������ٿ�S�O���@�:�+4@4�S�ߏ!?+��W��@������ٿ�S�O���@�:�+4@4�S�ߏ!?+��W��@��ͼP�ٿ��J��@��c�Y 4@.~�[��!?���0D�@��ͼP�ٿ��J��@��c�Y 4@.~�[��!?���0D�@�&Ov��ٿ���g�+�@T>ל�4@�����!?�Ό'��@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@C8u���ٿf�	;4��@,R/� 4@�KF���!?R�mq�@�ryݵٿ������@7v�� 4@�s{���!?0zc3�N�@����X�ٿ��G����@�5\M��3@��{�Ώ!?	�B�G��@����X�ٿ��G����@�5\M��3@��{�Ώ!?	�B�G��@����X�ٿ��G����@�5\M��3@��{�Ώ!?	�B�G��@����X�ٿ��G����@�5\M��3@��{�Ώ!?	�B�G��@����X�ٿ��G����@�5\M��3@��{�Ώ!?	�B�G��@�n�j-�ٿ�L���k�@.>� 4@�%����!?N�oΟ��@�n�j-�ٿ�L���k�@.>� 4@�%����!?N�oΟ��@�n�j-�ٿ�L���k�@.>� 4@�%����!?N�oΟ��@�n�j-�ٿ�L���k�@.>� 4@�%����!?N�oΟ��@���2�ٿ��j7��@$���f�3@2��j�!?���x"��@���2�ٿ��j7��@$���f�3@2��j�!?���x"��@�]p�̦ٿh��H��@�,h� 4@�.5�8�!?�m��j��@�]p�̦ٿh��H��@�,h� 4@�.5�8�!?�m��j��@�]p�̦ٿh��H��@�,h� 4@�.5�8�!?�m��j��@�]p�̦ٿh��H��@�,h� 4@�.5�8�!?�m��j��@�]p�̦ٿh��H��@�,h� 4@�.5�8�!?�m��j��@�#Eh�ٿ���\��@���h��3@8�;��!?��8G��@�#Eh�ٿ���\��@���h��3@8�;��!?��8G��@�#Eh�ٿ���\��@���h��3@8�;��!?��8G��@Í�X�ٿ[�TW�1�@wu�q��3@h�E���!?\E��U��@Í�X�ٿ[�TW�1�@wu�q��3@h�E���!?\E��U��@Í�X�ٿ[�TW�1�@wu�q��3@h�E���!?\E��U��@�1ʜٿ�*껪��@]�0Ҿ�3@��q��!?���O_�@�1ʜٿ�*껪��@]�0Ҿ�3@��q��!?���O_�@�,O�W�ٿ�<�U��@��gO� 4@F��׏!?��[���@�,O�W�ٿ�<�U��@��gO� 4@F��׏!?��[���@�,O�W�ٿ�<�U��@��gO� 4@F��׏!?��[���@��^�ٿۚ���Y�@]��p��3@	n@׏!?�[�&���@��^�ٿۚ���Y�@]��p��3@	n@׏!?�[�&���@��^�ٿۚ���Y�@]��p��3@	n@׏!?�[�&���@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@^r{���ٿ�)�����@25�� 4@���j͏!?Q��@t�nC�ٿ�l����@iU���4@��m���!?�������@t�nC�ٿ�l����@iU���4@��m���!?�������@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@{I��ߞٿ�r����@�=Eg 4@X���!?x��L�@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@Y.f�ٿ�� ���@������3@ۓ୏!?��K���@�M/]�ٿ9�X�\�@I���4@K����!?
�q�RL�@�M/]�ٿ9�X�\�@I���4@K����!?
�q�RL�@�M/]�ٿ9�X�\�@I���4@K����!?
�q�RL�@6�ܝٿ�s�~�@6�X[�4@�x�B��!?�CZ���@}�W'��ٿ����f�@%Co}�4@�K�Џ!?1&�x�8�@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@�:;2Q�ٿҥ�2�@���� 4@�%�b��!?9/�@+��@����ٿՠ � �@����4@� �˳�!?m���@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@��_j�ٿ��ZDѭ�@-���w�3@�5湱�!?���y�f�@�Z{p[�ٿ!��B=�@��|�4@�#l���!?�`��)�@�Z{p[�ٿ!��B=�@��|�4@�#l���!?�`��)�@�Z{p[�ٿ!��B=�@��|�4@�#l���!?�`��)�@�Z{p[�ٿ!��B=�@��|�4@�#l���!?�`��)�@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@`O+S��ٿ�fD,6��@%�@�"�3@�_*x��!?`���B��@i�Lc�ٿ�!��r�@c��o 4@�X��t�!?!�FIC�@i�Lc�ٿ�!��r�@c��o 4@�X��t�!?!�FIC�@i�Lc�ٿ�!��r�@c��o 4@�X��t�!?!�FIC�@���ٿ��c���@,G%74@�|�y�!?J3@�I��@���ٿ��c���@,G%74@�|�y�!?J3@�I��@���ٿ��c���@,G%74@�|�y�!?J3@�I��@���ٿ��c���@,G%74@�|�y�!?J3@�I��@K�	[�ٿ`L����@�F�>1 4@�xЀ�!?�^O���@K�	[�ٿ`L����@�F�>1 4@�xЀ�!?�^O���@����ٿcX��<��@>ۣ|Y 4@��%ɏ!?׀�n�@����ٿcX��<��@>ۣ|Y 4@��%ɏ!?׀�n�@����ٿcX��<��@>ۣ|Y 4@��%ɏ!?׀�n�@����ٿcX��<��@>ۣ|Y 4@��%ɏ!?׀�n�@����ٿcX��<��@>ۣ|Y 4@��%ɏ!?׀�n�@�ڀ�1�ٿ�9*d�@Ǫy|,4@���߻�!?�@�1P�@�ڀ�1�ٿ�9*d�@Ǫy|,4@���߻�!?�@�1P�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@qඨ3�ٿ�ֿb��@̺��y�3@[����!?�ޮ�G�@�*����ٿ�޷���@o$� 4@iw)���!?���ԡ�@�*����ٿ�޷���@o$� 4@iw)���!?���ԡ�@R(���ٿ>��g�@W����3@��⹏!?3�Av)+�@R(���ٿ>��g�@W����3@��⹏!?3�Av)+�@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@\��5S�ٿ���3i��@|E[�#�3@��O̏!?���72��@�Fy��ٿSt����@K���L4@��οɏ!?��?�$��@Ƴ�oܙٿ|�����@yi��4@ �U�!?1��<��@�|�j�ٿ���S��@��p�.4@V����!?��_X��@�|�j�ٿ���S��@��p�.4@V����!?��_X��@�|�j�ٿ���S��@��p�.4@V����!?��_X��@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@secp(�ٿ�L����@��Z 4@c$���!?J��p�@Y�/,�ٿ�Czv�;�@s�<�"�3@"�ը�!?�Dc�"]�@Y�/,�ٿ�Czv�;�@s�<�"�3@"�ը�!?�Dc�"]�@��{�\�ٿ���� /�@�Wt 4@wI �!?�ȳR�@��{�\�ٿ���� /�@�Wt 4@wI �!?�ȳR�@��{�\�ٿ���� /�@�Wt 4@wI �!?�ȳR�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@��Kݢٿt��&�@�
zp@ 4@=S�{�!?(@+z�y�@G�コ�ٿ'�!"6�@����3@�	�q�!?��k��@G�コ�ٿ'�!"6�@����3@�	�q�!?��k��@G�コ�ٿ'�!"6�@����3@�	�q�!?��k��@G�コ�ٿ'�!"6�@����3@�	�q�!?��k��@G�コ�ٿ'�!"6�@����3@�	�q�!?��k��@ET��M�ٿ��T��@���f4@V��{��!?t�5���@	y�\ڢٿ.��A��@�Yq�|4@x���!?o`��~��@E]7��ٿ�w]��@J�G�4@G	�J��!?P�*� ��@E]7��ٿ�w]��@J�G�4@G	�J��!?P�*� ��@6�ٿ��\���@�A�%/4@���"�!?c��;�@6�ٿ��\���@�A�%/4@���"�!?c��;�@6�ٿ��\���@�A�%/4@���"�!?c��;�@6�ٿ��\���@�A�%/4@���"�!?c��;�@��C>�ٿ�}�'��@�f/� 4@U�8}�!?{�2�y�@��C>�ٿ�}�'��@�f/� 4@U�8}�!?{�2�y�@��C>�ٿ�}�'��@�f/� 4@U�8}�!?{�2�y�@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@Z^�I|�ٿ��H�0��@[�'z�3@��s�!?;�R���@uLY�ٿ�S1�~��@��MK9�3@����!?]g0ڼ��@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@�X���ٿW�<>�*�@��w�3@n�&̏!?�`țԈ�@4F(�ۨٿ,���k�@|ss�B4@������!??*��@4F(�ۨٿ,���k�@|ss�B4@������!??*��@^X\�0�ٿzl�T<�@@���1�3@Rڴs��!?�ّ����@^X\�0�ٿzl�T<�@@���1�3@Rڴs��!?�ّ����@^X\�0�ٿzl�T<�@@���1�3@Rڴs��!?�ّ����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@y� ��ٿqH�l�@�^��4@Lq`���!?_����@L�(�ٿ�wf��?�@A7�c�3@ߊ�聏!?� �mG�@j�ydc�ٿg�x܄��@����b4@^5dT�!?�qG�a�@j�ydc�ٿg�x܄��@����b4@^5dT�!?�qG�a�@��?m�ٿ#�"$���@?�� 4@ȸ]3��!?�f*	���@��?m�ٿ#�"$���@?�� 4@ȸ]3��!?�f*	���@��?m�ٿ#�"$���@?�� 4@ȸ]3��!?�f*	���@��?m�ٿ#�"$���@?�� 4@ȸ]3��!?�f*	���@��]�ٿ	�ċ��@��u��3@5p1kq�!?�}���@��]�ٿ	�ċ��@��u��3@5p1kq�!?�}���@[-x,��ٿ~�����@�9"�� 4@��ć�!?��{�C~�@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@����ٿF�h~��@�	�� 4@#�F��!?�"r��@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@.X���ٿ����@��^.��3@���:|�!?M���@�����ٿN��1���@6�����3@��gYڏ!? F��]:�@���Y�ٿ�1Z��s�@<6�ζ�3@d�<�I�!?�i:K�@���Y�ٿ�1Z��s�@<6�ζ�3@d�<�I�!?�i:K�@���Y�ٿ�1Z��s�@<6�ζ�3@d�<�I�!?�i:K�@���Y�ٿ�1Z��s�@<6�ζ�3@d�<�I�!?�i:K�@Br��ٿ��EP�@q�f�3@����]�!?-=U�@Br��ٿ��EP�@q�f�3@����]�!?-=U�@Br��ٿ��EP�@q�f�3@����]�!?-=U�@"����ٿ�E����@���*j�3@<_V6��!?�Rv��@Ԍo �ٿ�y|pA�@�ZѤ�3@sё6u�!?a�/A�_�@���uT�ٿk��6���@O,�` 4@# lc�!?M)�#_�@���uT�ٿk��6���@O,�` 4@# lc�!?M)�#_�@���uT�ٿk��6���@O,�` 4@# lc�!?M)�#_�@���uT�ٿk��6���@O,�` 4@# lc�!?M)�#_�@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@�2w�ٿ�=y�(}�@#�u��4@��&ُ!?�Q���@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@L��A�ٿ1���h��@ل���3@�f��!?I Ȫe�@~�@�?�ٿrJ
��X�@�i*�� 4@�a�ȏ!?�-�7}�@���ٿ]3r{�@D�~'4@��(�!?�?i�t��@���ٿ]3r{�@D�~'4@��(�!?�?i�t��@���ٿ]3r{�@D�~'4@��(�!?�?i�t��@���ٿ]3r{�@D�~'4@��(�!?�?i�t��@ W޸�ٿ�G�Z�@��4@ق��!?�F��H�@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@��e(�ٿ�?�L�h�@�t�� 4@lVAE��!?_y�����@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�[O�8�ٿ(�
"`��@�=R� 4@S���!?a��7}�@�����ٿl��/��@�|����3@22޴�!?�k�ٓ��@�����ٿl��/��@�|����3@22޴�!?�k�ٓ��@�����ٿl��/��@�|����3@22޴�!?�k�ٓ��@��/O��ٿ�s|���@���I��3@|�u��!?%�\u��@��/O��ٿ�s|���@���I��3@|�u��!?%�\u��@��@���ٿ� ` �S�@T�ɫ�3@�`ޏ!?�ܗ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@yI�&��ٿOUt��@
#�2`�3@F��!��!?-�$Ӿ��@�.�x�ٿ�{8�Y��@)�m|R�3@��V��!?��|��O�@�.�x�ٿ�{8�Y��@)�m|R�3@��V��!?��|��O�@�.�x�ٿ�{8�Y��@)�m|R�3@��V��!?��|��O�@	E~�k�ٿaR����@���>�3@[��ߏ!?S��JM�@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��WA�ٿ^�崋��@�T=�3@&qj���!?�a���@��{Xm�ٿ�E�RU�@�X�NW�3@� ��!?|��A�@��{Xm�ٿ�E�RU�@�X�NW�3@� ��!?|��A�@��{Xm�ٿ�E�RU�@�X�NW�3@� ��!?|��A�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@`q�b��ٿ5V�#NW�@m[��^ 4@ʅ:��!?w��9�@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@���+�ٿjUl]c�@����� 4@�hw��!?�>���@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@�1�O�ٿ�w�t���@��y 4@\t��Ǐ!?	܉�O�@V�q�ٿ3����@6�~ 4@��_�׏!?"LCK�'�@V�q�ٿ3����@6�~ 4@��_�׏!?"LCK�'�@V�q�ٿ3����@6�~ 4@��_�׏!?"LCK�'�@Uh��n�ٿ�7�|��@+l�� 4@�daȏ!?Ϛ� ��@Uh��n�ٿ�7�|��@+l�� 4@�daȏ!?Ϛ� ��@Uh��n�ٿ�7�|��@+l�� 4@�daȏ!?Ϛ� ��@�$��(�ٿ�Lg�A��@)w�1[ 4@W���-�!?k���1*�@�$��(�ٿ�Lg�A��@)w�1[ 4@W���-�!?k���1*�@�$��(�ٿ�Lg�A��@)w�1[ 4@W���-�!?k���1*�@�$��(�ٿ�Lg�A��@)w�1[ 4@W���-�!?k���1*�@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@��i�ٿ�!����@*v��B�3@�3M�!?��c��@���랤ٿ�EI7Y��@��%��4@֩O�H�!?s��X�@���~�ٿX	;����@�M��4@V�N���!?x��4S�@��(�M�ٿf֐����@�O��4@��,�ɏ!?G=�@��(�M�ٿf֐����@�O��4@��,�ɏ!?G=�@��(�M�ٿf֐����@�O��4@��,�ɏ!?G=�@��M�^�ٿ��!��m�@�a>��4@\)���!?�Snd�(�@��M�^�ٿ��!��m�@�a>��4@\)���!?�Snd�(�@��M�^�ٿ��!��m�@�a>��4@\)���!?�Snd�(�@��M�^�ٿ��!��m�@�a>��4@\)���!?�Snd�(�@��M�^�ٿ��!��m�@�a>��4@\)���!?�Snd�(�@��iY��ٿ���%BO�@f��~� 4@�j�p�!?V۲�n�@��iY��ٿ���%BO�@f��~� 4@�j�p�!?V۲�n�@��iY��ٿ���%BO�@f��~� 4@�j�p�!?V۲�n�@�VI�Şٿ��:d�@�@��I� 4@���r��!?����<�@�VI�Şٿ��:d�@�@��I� 4@���r��!?����<�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@�B��,�ٿ���(���@I�h4@ :1��!?Ԉ�Wˑ�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@%D�ٿҨ"a���@U��n4@FEI�7�!?�jn~�@�c��l�ٿ0��0��@B��hQ 4@�k�t�!?ԂO�n��@Ag���ٿ/��:��@TP�[d 4@�t��q�!?�p�ç5�@Ag���ٿ/��:��@TP�[d 4@�t��q�!?�p�ç5�@Ag���ٿ/��:��@TP�[d 4@�t��q�!?�p�ç5�@Ag���ٿ/��:��@TP�[d 4@�t��q�!?�p�ç5�@��9�Ȩٿ�;�'\�@���� 4@Ժ��!?1](@��@��9�Ȩٿ�;�'\�@���� 4@Ժ��!?1](@��@��9�Ȩٿ�;�'\�@���� 4@Ժ��!?1](@��@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�X���ٿ�e���@���� 4@��W��!?�K]�,x�@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@�Ff��ٿ���3��@��Y�4@����E�!?�P ���@%j�U�ٿiY%�p�@%���4@�G�q��!?�zh}?�@%j�U�ٿiY%�p�@%���4@�G�q��!?�zh}?�@%j�U�ٿiY%�p�@%���4@�G�q��!?�zh}?�@*wqD1�ٿ#���@�o��3@��[���!?�w�8��@*wqD1�ٿ#���@�o��3@��[���!?�w�8��@D�uA�ٿU��z&�@��x! 4@�DQ��!?��Js��@D�uA�ٿU��z&�@��x! 4@�DQ��!?��Js��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@QY'Oc�ٿ[^��Q9�@��S�� 4@3J��!?����]��@_�>�ʣٿ��;����@��_��3@���w��!?C�#үI�@_�>�ʣٿ��;����@��_��3@���w��!?C�#үI�@_�>�ʣٿ��;����@��_��3@���w��!?C�#үI�@_�>�ʣٿ��;����@��_��3@���w��!?C�#үI�@1򟄤ٿ����۸�@`�� �3@��1Ώ!?)�N���@1򟄤ٿ����۸�@`�� �3@��1Ώ!?)�N���@�t��ٿ�do,M�@#�)��3@��n��!?�5���@�t��ٿ�do,M�@#�)��3@��n��!?�5���@�t��ٿ�do,M�@#�)��3@��n��!?�5���@:d&�$�ٿ��9��3�@2<"���3@�o�͏!?c���Si�@:d&�$�ٿ��9��3�@2<"���3@�o�͏!?c���Si�@:d&�$�ٿ��9��3�@2<"���3@�o�͏!?c���Si�@��o4˪ٿQG�)J�@�է�`�3@J����!?ѥŵ���@)Xl5�ٿ$��>��@����3@Ȅ�S�!?����@�[��ٿP 	�b�@0�h���3@/��<	�!?}L��{�@�[��ٿP 	�b�@0�h���3@/��<	�!?}L��{�@� �F�ٿ���y��@�h��3@����d�!?��\q�&�@��Z<��ٿU������@g����3@FS�䍏!?��ɟX��@��Z<��ٿU������@g����3@FS�䍏!?��ɟX��@��Z<��ٿU������@g����3@FS�䍏!?��ɟX��@<�i���ٿ��R��@�6�u��3@�n�ؘ�!?�ꡬO �@۝4�Ԩٿ��fI�e�@�N	�H�3@v�׳�!?������@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�c�ٿ�CM��i�@ς�� �3@�6V�!?���h�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@�Ѓ�ٿ	�����@<��cq�3@�ί�!?����s�@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@(ˍ⦢ٿ�m�D�)�@���&��3@�iD��!?'~Y���@�V�}�ٿ����;�@te I�3@/;�ԏ!?�Z�P��@�V�}�ٿ����;�@te I�3@/;�ԏ!?�Z�P��@�V�}�ٿ����;�@te I�3@/;�ԏ!?�Z�P��@�V�}�ٿ����;�@te I�3@/;�ԏ!?�Z�P��@��[�ٿ���~���@�7)�J4@����!?f�OyX�@��[�ٿ���~���@�7)�J4@����!?f�OyX�@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@�8Re��ٿ�sfQ=1�@MmΩ4@!�Q3��!?�t�O$��@Rf�!�ٿ����"�@� R4@�4$��!?�(H��@U���ٿ��[��@� �4@�a�>�!?��h����@F}-�E�ٿvy��M�@�a^V�4@�Ń}ԏ!?�C��y�@F}-�E�ٿvy��M�@�a^V�4@�Ń}ԏ!?�C��y�@F}-�E�ٿvy��M�@�a^V�4@�Ń}ԏ!?�C��y�@f_�آٿD��K���@�Q*T�4@a�<�<�!?"�ُ��@f_�آٿD��K���@�Q*T�4@a�<�<�!?"�ُ��@f_�آٿD��K���@�Q*T�4@a�<�<�!?"�ُ��@f_�آٿD��K���@�Q*T�4@a�<�<�!?"�ُ��@f_�آٿD��K���@�Q*T�4@a�<�<�!?"�ُ��@����ٿ� ��A=�@Ϣ]m4@���!?�{&/m��@����ٿ� ��A=�@Ϣ]m4@���!?�{&/m��@����ٿ� ��A=�@Ϣ]m4@���!?�{&/m��@����ٿ� ��A=�@Ϣ]m4@���!?�{&/m��@���N�ٿإ���@q9]j�4@�����!?��Z-�@���N�ٿإ���@q9]j�4@�����!?��Z-�@���N�ٿإ���@q9]j�4@�����!?��Z-�@F�Ј�ٿ}����@GD = 4@�nn��!?�-��h�@F�Ј�ٿ}����@GD = 4@�nn��!?�-��h�@F�Ј�ٿ}����@GD = 4@�nn��!?�-��h�@F�Ј�ٿ}����@GD = 4@�nn��!?�-��h�@F�Ј�ٿ}����@GD = 4@�nn��!?�-��h�@t4���ٿ^�3ʼ��@3���s4@p	4��!?A��} $�@t4���ٿ^�3ʼ��@3���s4@p	4��!?A��} $�@��}���ٿu*��k��@�c`��3@�܏!?2��j�@�"��ٿ��l�l�@N0]_�3@ô�5w�!?!�k��@�"��ٿ��l�l�@N0]_�3@ô�5w�!?!�k��@�"��ٿ��l�l�@N0]_�3@ô�5w�!?!�k��@�"��ٿ��l�l�@N0]_�3@ô�5w�!?!�k��@�"��ٿ��l�l�@N0]_�3@ô�5w�!?!�k��@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@�՛ٿa���̌�@��%<4@�D����!?�|���q�@ɎnR��ٿ@�s��d�@x�P�4@<L�y�!?�N�����@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@6{[+�ٿRv}�@�@�U3o��3@��M���!?i�}��;�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@|��ڞٿ]j-�c�@�5WEO4@���ɏ!?�5�3ۣ�@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@{�ۤٿPNt���@�}$�4@Wɶ�!?�������@�V'蔝ٿ��P6��@��jz�4@k&�a�!?h��@�V'蔝ٿ��P6��@��jz�4@k&�a�!?h��@d�k� �ٿ頼���@ws��4@���w�!?}C��$��@d�k� �ٿ頼���@ws��4@���w�!?}C��$��@d�k� �ٿ頼���@ws��4@���w�!?}C��$��@d�k� �ٿ頼���@ws��4@���w�!?}C��$��@���ٿ��?��@���4@��%=�!?�g��B�@�H�ɼ�ٿ������@X��lx4@�ΰ���!?W%`��@�H�ɼ�ٿ������@X��lx4@�ΰ���!?W%`��@�H�ɼ�ٿ������@X��lx4@�ΰ���!?W%`��@��?�ٿ��n���@���'4@���!?��G��@��?�ٿ��n���@���'4@���!?��G��@���7ơٿZ:��;��@MAܫ4@r;O{2�!?���m�@���7ơٿZ:��;��@MAܫ4@r;O{2�!?���m�@���7ơٿZ:��;��@MAܫ4@r;O{2�!?���m�@���7ơٿZ:��;��@MAܫ4@r;O{2�!?���m�@���7ơٿZ:��;��@MAܫ4@r;O{2�!?���m�@b!V��ٿ��:3��@Sq��4@$�>��!?`�)�'^�@b!V��ٿ��:3��@Sq��4@$�>��!?`�)�'^�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@t4���ٿ=��@�E�� 4@���k�!?ι0�Pp�@u��q�ٿk�M���@ I�1� 4@)B]�!?�⡆uC�@u��q�ٿk�M���@ I�1� 4@)B]�!?�⡆uC�@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@65��%�ٿ��3H�@�P"�_4@��ɏ!?O�w���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@4M�:�ٿ6�-~}�@~a4h 4@j�G�t�!?hX}���@"b�ٿ��G����@/�t�= 4@�=D��!?Τb���@"b�ٿ��G����@/�t�= 4@�=D��!?Τb���@1���X�ٿ������@,��� 4@nd0��!?�0E���@1���X�ٿ������@,��� 4@nd0��!?�0E���@1���X�ٿ������@,��� 4@nd0��!?�0E���@1���X�ٿ������@,��� 4@nd0��!?�0E���@1���X�ٿ������@,��� 4@nd0��!?�0E���@1���X�ٿ������@,��� 4@nd0��!?�0E���@��L�u�ٿ:����@� 4@}�s���!?{�Ad�@��L�u�ٿ:����@� 4@}�s���!?{�Ad�@��L�u�ٿ:����@� 4@}�s���!?{�Ad�@��L�u�ٿ:����@� 4@}�s���!?{�Ad�@��L�u�ٿ:����@� 4@}�s���!?{�Ad�@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@P<�@a�ٿ8�_�Л�@|�n� 4@Wn{�Y�!?s�����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@k��H�ٿ���w��@��V��3@���v�!?�z����@���ٿ��&X�@��zg��3@�V�$�!?�;��n�@���ٿ��&X�@��zg��3@�V�$�!?�;��n�@�J�H�ٿ�>#O��@�z�]�3@yw��C�!?J�@�vM�@�J�H�ٿ�>#O��@�z�]�3@yw��C�!?J�@�vM�@Y:^�$�ٿ��I��@�b�� 4@�n$�i�!?�����@Y:^�$�ٿ��I��@�b�� 4@�n$�i�!?�����@Y:^�$�ٿ��I��@�b�� 4@�n$�i�!?�����@Y:^�$�ٿ��I��@�b�� 4@�n$�i�!?�����@Y:^�$�ٿ��I��@�b�� 4@�n$�i�!?�����@�19|�ٿ���7H�@F����3@��	v��!?G)
���@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@�e��ٿ�ԊPɣ�@	�B�# 4@Q��b�!?�'����@��F��ٿ��e���@���� 4@V��S��!?���L�	�@��F��ٿ��e���@���� 4@V��S��!?���L�	�@��F��ٿ��e���@���� 4@V��S��!?���L�	�@��F��ٿ��e���@���� 4@V��S��!?���L�	�@��0]�ٿ�M���@�a�k[�3@�b���!?�d���@��0]�ٿ�M���@�a�k[�3@�b���!?�d���@��0]�ٿ�M���@�a�k[�3@�b���!?�d���@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@û�6͠ٿ�����@NA:q��3@6��﷏!?0���t��@W�6�ͦٿ6��9�3�@��a!�4@\�v�!?��ɋ��@W�6�ͦٿ6��9�3�@��a!�4@\�v�!?��ɋ��@W�6�ͦٿ6��9�3�@��a!�4@\�v�!?��ɋ��@��!$�ٿHߔ$j�@8�^�3@g���ُ!?�v���@��!$�ٿHߔ$j�@8�^�3@g���ُ!?�v���@��!$�ٿHߔ$j�@8�^�3@g���ُ!?�v���@�ʺ�[�ٿ��1�+�@��4@"=.��!?:}5����@�ʺ�[�ٿ��1�+�@��4@"=.��!?:}5����@�ʺ�[�ٿ��1�+�@��4@"=.��!?:}5����@�ʺ�[�ٿ��1�+�@��4@"=.��!?:}5����@�d�ٿ=�z�@�Dx4@�aif�!?�O�d�(�@�d�ٿ=�z�@�Dx4@�aif�!?�O�d�(�@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@qX��1�ٿv�Z;��@�cZ�64@��P���!?ӇO�9��@ 3e��ٿ|.̂s�@�`LQj4@���!?�5�SK�@ 3e��ٿ|.̂s�@�`LQj4@���!?�5�SK�@ 3e��ٿ|.̂s�@�`LQj4@���!?�5�SK�@ 3e��ٿ|.̂s�@�`LQj4@���!?�5�SK�@ 3e��ٿ|.̂s�@�`LQj4@���!?�5�SK�@!�rﴟٿm��t�@7>��3@{�Z���!?�x�14��@!�rﴟٿm��t�@7>��3@{�Z���!?�x�14��@����ٿ��~���@~;����3@�WR#�!?�F�v���@> <(��ٿ�]�`��@!�"��4@�;�l��!?�c�i���@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@�$T��ٿk'�({��@���*� 4@rM��[�!?�)�6K�@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@-��G�ٿ��:��@"kЯ��3@�/�RZ�!?`$��@w�bf��ٿ��k���@��� 4@��b�m�!?E3-�M��@w�bf��ٿ��k���@��� 4@��b�m�!?E3-�M��@w�bf��ٿ��k���@��� 4@��b�m�!?E3-�M��@³��ٿ�B����@��jh�3@@�kT�!?����m��@³��ٿ�B����@��jh�3@@�kT�!?����m��@³��ٿ�B����@��jh�3@@�kT�!?����m��@³��ٿ�B����@��jh�3@@�kT�!?����m��@�dy%)�ٿ�]ymĚ�@or��3@��N���!?�M6m�@�dy%)�ٿ�]ymĚ�@or��3@��N���!?�M6m�@�dy%)�ٿ�]ymĚ�@or��3@��N���!?�M6m�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@)}P�șٿי���@?,t�S4@S�o���!?�Wv�c�@����ٿ�P�vF�@'�ܔr�3@$I�!?7C�/���@����ٿ�P�vF�@'�ܔr�3@$I�!?7C�/���@�;�뽪ٿ]o���x�@���8��3@�]�P�!?\j�9ȵ�@�;�뽪ٿ]o���x�@���8��3@�]�P�!?\j�9ȵ�@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@����ٿ!-#���@��c 4@�Bgʎ�!?((�J��@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@?���ٿX�*_��@����4@����!?���� i�@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@s��ޟٿ	,�Q��@g֭� 4@�|���!?��0j���@n�N�0�ٿ�ł���@�0Oc�4@Q����!?E\����@n�N�0�ٿ�ł���@�0Oc�4@Q����!?E\����@n�N�0�ٿ�ł���@�0Oc�4@Q����!?E\����@����Ϥٿ��ng�@5�h�
 4@�H=qя!?y�J*t�@����Ϥٿ��ng�@5�h�
 4@�H=qя!?y�J*t�@����Ϥٿ��ng�@5�h�
 4@�H=qя!?y�J*t�@l�k�~�ٿW��v��@�R2W� 4@f��^��!?�B(%��@Uv�PT�ٿǩK_J�@��m�}�3@ѻ�J��!?&G�)�H�@�+Z�ٿh���'�@v�	"� 4@�#vÏ!?٧r�C�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@qݧU)�ٿ_}&��Y�@�@x�� 4@G�}+�!?��.p�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@4�}1�ٿ;�K L)�@
%b� 4@;R��E�!?�� �R�@� <F�ٿMc��,�@�'�e64@�c(�!?۵����@BX@D�ٿ�6_�M�@}�u�| 4@��%��!?wQ<\�@BX@D�ٿ�6_�M�@}�u�| 4@��%��!?wQ<\�@Am�\��ٿM�!*�@"ת���3@�����!?������@���ٿ����>��@�-��m�3@H.�)L�!?0�`�ӯ�@���ٿ����>��@�-��m�3@H.�)L�!?0�`�ӯ�@���ٿ����>��@�-��m�3@H.�)L�!?0�`�ӯ�@���ٿ����>��@�-��m�3@H.�)L�!?0�`�ӯ�@���ٿ����>��@�-��m�3@H.�)L�!?0�`�ӯ�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@/x�1 �ٿMb����@dY����3@�QEg=�!?[���H3�@@�Q$ƙٿ$�L�B��@0I����3@�<���!?J{I��@@�Q$ƙٿ$�L�B��@0I����3@�<���!?J{I��@@�Q$ƙٿ$�L�B��@0I����3@�<���!?J{I��@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@���{�ٿ-�>�a��@5��AS�3@��ŏ!?!Hy��&�@Ol����ٿ@q���@u�f^;�3@��&��!?z�xw��@Ol����ٿ@q���@u�f^;�3@��&��!?z�xw��@Ol����ٿ@q���@u�f^;�3@��&��!?z�xw��@Ol����ٿ@q���@u�f^;�3@��&��!?z�xw��@Ol����ٿ@q���@u�f^;�3@��&��!?z�xw��@�0�C��ٿ�(+����@qT�R��3@3<`>+�!?D�����@8/}jڦٿ�g�[��@}�L 4@�? C�!?�ӟQ�f�@8/}jڦٿ�g�[��@}�L 4@�? C�!?�ӟQ�f�@V�۶�ٿ�3�6�@35�/4@��=��!?���;�y�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@M�B�g�ٿ�<�~��@�b�1C�3@s� f�!?���}�@Y��F �ٿ��'�s�@���'2�3@e���!?y;th�@Y��F �ٿ��'�s�@���'2�3@e���!?y;th�@Y��F �ٿ��'�s�@���'2�3@e���!?y;th�@Y��F �ٿ��'�s�@���'2�3@e���!?y;th�@O��f�ٿ΀��@%av��3@_��=I�!?�S��z�@O��f�ٿ΀��@%av��3@_��=I�!?�S��z�@O��f�ٿ΀��@%av��3@_��=I�!?�S��z�@{�5��ٿX����@M��* 4@ �= 5�!?��{��o�@{�5��ٿX����@M��* 4@ �= 5�!?��{��o�@{�5��ٿX����@M��* 4@ �= 5�!?��{��o�@{�5��ٿX����@M��* 4@ �= 5�!?��{��o�@5���ٿ�R����@:����3@+��=�!?�k�rn!�@5���ٿ�R����@:����3@+��=�!?�k�rn!�@5���ٿ�R����@:����3@+��=�!?�k�rn!�@5���ٿ�R����@:����3@+��=�!?�k�rn!�@��Z�ٿ�Q�`%�@yx����3@�b�21�!?��9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@w�/S��ٿ�JI���@╼Ҫ�3@.C:�@�!?x9���@����5�ٿ�U�yk�@����4@ \���!?��U��@����5�ٿ�U�yk�@����4@ \���!?��U��@����5�ٿ�U�yk�@����4@ \���!?��U��@����5�ٿ�U�yk�@����4@ \���!?��U��@o%4ܕٿ�DJO_w�@�h��4@�wÌ��!?���?�@o%4ܕٿ�DJO_w�@�h��4@�wÌ��!?���?�@o%4ܕٿ�DJO_w�@�h��4@�wÌ��!?���?�@o%4ܕٿ�DJO_w�@�h��4@�wÌ��!?���?�@=�	�ٿ�J!���@`'c��4@����!?����@=�	�ٿ�J!���@`'c��4@����!?����@=�	�ٿ�J!���@`'c��4@����!?����@=�	�ٿ�J!���@`'c��4@����!?����@���^��ٿ3��K)��@@TpW
4@ �s_��!?ҩ�1�4�@���^��ٿ3��K)��@@TpW
4@ �s_��!?ҩ�1�4�@���^��ٿ3��K)��@@TpW
4@ �s_��!?ҩ�1�4�@���^��ٿ3��K)��@@TpW
4@ �s_��!?ҩ�1�4�@���^��ٿ3��K)��@@TpW
4@ �s_��!?ҩ�1�4�@�ú�۔ٿb����@̀K| 4@��XO�!?46����@�ú�۔ٿb����@̀K| 4@��XO�!?46����@�ú�۔ٿb����@̀K| 4@��XO�!?46����@�ú�۔ٿb����@̀K| 4@��XO�!?46����@���q��ٿ��Һ�@�!��3@��.J�!?�����=�@���q��ٿ��Һ�@�!��3@��.J�!?�����=�@���q��ٿ��Һ�@�!��3@��.J�!?�����=�@���q��ٿ��Һ�@�!��3@��.J�!?�����=�@f��~b�ٿ�iϴ��@�@�6� 4@-�4��!?�l{��J�@�Ae1��ٿ�6�I���@BM��3@�>o�t�!?al_�'�@�1���ٿXŲ* �@X����3@��(�!?[}Qq�@�1���ٿXŲ* �@X����3@��(�!?[}Qq�@�1���ٿXŲ* �@X����3@��(�!?[}Qq�@�1���ٿXŲ* �@X����3@��(�!?[}Qq�@�1���ٿXŲ* �@X����3@��(�!?[}Qq�@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@����/�ٿ����t�@6G`���3@u>�ڤ�!?�����@���즙ٿ�t	�LS�@�'�� 4@j3
��!?�r����@���즙ٿ�t	�LS�@�'�� 4@j3
��!?�r����@���즙ٿ�t	�LS�@�'�� 4@j3
��!?�r����@���즙ٿ�t	�LS�@�'�� 4@j3
��!?�r����@����	�ٿ�2��8�@d6JL� 4@���T�!?�E�4�@T�דٿ��a)ͮ�@�Od� 4@�0Mʏ!?nl����@E{�a�ٿ{���@,?��3@K��ӏ!?�S��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@>��/�ٿp���wi�@�&c��3@ ��V*�!?5b�,=��@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@Nd���ٿyJKn���@����%4@���!?-s$W�Q�@���iէٿC�Ut:��@���yP4@e�	�Ǐ!?�κ�::�@|m�+�ٿ��2m��@2P�74@Y�!?@�(��@g��9�ٿF��Yn�@5����3@o�K��!?�F�U��@���c'�ٿMf�L���@P	����3@؇&��!?�l��F�@���c'�ٿMf�L���@P	����3@؇&��!?�l��F�@���c'�ٿMf�L���@P	����3@؇&��!?�l��F�@���c'�ٿMf�L���@P	����3@؇&��!?�l��F�@���c'�ٿMf�L���@P	����3@؇&��!?�l��F�@_Q$�@�ٿYD7�d��@hX�#�4@j�%��!?!z�55�@_Q$�@�ٿYD7�d��@hX�#�4@j�%��!?!z�55�@_Q$�@�ٿYD7�d��@hX�#�4@j�%��!?!z�55�@_Q$�@�ٿYD7�d��@hX�#�4@j�%��!?!z�55�@m&�<��ٿ5� sS�@WW�p� 4@�R�ߏ!?�����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@H�:ۛٿ����@a`E�4@-�����!?F�l����@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@-^�ٿ������@J�=�.4@�����!?3�k@���@%�q��ٿ�l�0t��@?��o4@
����!?('�Q��@%�q��ٿ�l�0t��@?��o4@
����!?('�Q��@%�q��ٿ�l�0t��@?��o4@
����!?('�Q��@��b��ٿ�Jd��@֚�4@�""ن�!?����7�@��b��ٿ�Jd��@֚�4@�""ن�!?����7�@��b��ٿ�Jd��@֚�4@�""ن�!?����7�@��b��ٿ�Jd��@֚�4@�""ن�!?����7�@��b��ٿ�Jd��@֚�4@�""ن�!?����7�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@n
	n�ٿI����@�.Qd`4@h��!?oQ��,�@˼��J�ٿl��*�@G�L�4@S��*��!?��d�A�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@�nd��ٿ�{@���@ʧ��4@b�$|�!?9�9*�@+u��˙ٿcư��@�L�$4@x����!?b��(��@+u��˙ٿcư��@�L�$4@x����!?b��(��@+u��˙ٿcư��@�L�$4@x����!?b��(��@+u��˙ٿcư��@�L�$4@x����!?b��(��@�>��p�ٿ�7!��@�� 4@�O#��!?3�˧{f�@�>��p�ٿ�7!��@�� 4@�O#��!?3�˧{f�@�)H��ٿm�G��K�@҅ԔM 4@��R�!?��-R��@�)H��ٿm�G��K�@҅ԔM 4@��R�!?��-R��@�)H��ٿm�G��K�@҅ԔM 4@��R�!?��-R��@�)H��ٿm�G��K�@҅ԔM 4@��R�!?��-R��@�)H��ٿm�G��K�@҅ԔM 4@��R�!?��-R��@�׺���ٿ&���X�@�g��4@l�|���!?��ާQ�@|���ʥٿI�Pޖ�@1��4@_�4���!?wJ"�G�@|���ʥٿI�Pޖ�@1��4@_�4���!?wJ"�G�@|���ʥٿI�Pޖ�@1��4@_�4���!?wJ"�G�@�� k�ٿ�aW-B�@\@�w4@5��!?v���S�@�� k�ٿ�aW-B�@\@�w4@5��!?v���S�@�� k�ٿ�aW-B�@\@�w4@5��!?v���S�@�� k�ٿ�aW-B�@\@�w4@5��!?v���S�@g�scq�ٿ�R[G���@Ə��4@n��+�!?���w5N�@g�scq�ٿ�R[G���@Ə��4@n��+�!?���w5N�@g�scq�ٿ�R[G���@Ə��4@n��+�!?���w5N�@���ٿ���V��@��H �4@��xI�!?���E�
�@���ٿ���V��@��H �4@��xI�!?���E�
�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@�y��ٿq��n��@T����4@g9�%��!?/炵Y%�@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@#�2m�ٿ��(��@�ڂ4 4@kT׿�!?Q2)�W��@�!����ٿHn'IZ6�@Q3��Z 4@���!?�T�S���@�!����ٿHn'IZ6�@Q3��Z 4@���!?�T�S���@��L�ٿ�0�+[ �@�A�4@d�S��!?b�(�@��@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@C �g�ٿ�F�7{6�@���4@ˢ7��!?ʝ�XNF�@&$B�_�ٿyCO���@ m `�3@@�7O�!? -�f��@&$B�_�ٿyCO���@ m `�3@@�7O�!? -�f��@����J�ٿ:��YW�@<�����3@(���!?,��Դ��@����J�ٿ:��YW�@<�����3@(���!?,��Դ��@����J�ٿ:��YW�@<�����3@(���!?,��Դ��@����J�ٿ:��YW�@<�����3@(���!?,��Դ��@Ի���ٿ�н��*�@O�3"� 4@L;*�!?Mr��@�8��ٿ{�ș��@�.2t4@Q��9�!?��%�~��@�8��ٿ{�ș��@�.2t4@Q��9�!?��%�~��@�8��ٿ{�ș��@�.2t4@Q��9�!?��%�~��@Rk�<J�ٿ4p�}{K�@�N�z?4@a�fb��!?�r	ߤ��@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@9ZZ�z�ٿ�!��6��@�6]�4@�`X�!?�Kq`���@(Nh���ٿa�%�@����Z4@�m�)��!?�y�Q$�@(Nh���ٿa�%�@����Z4@�m�)��!?�y�Q$�@j�9�h�ٿkzl��@Զ��t4@U3n���!?7y��>��@j�9�h�ٿkzl��@Զ��t4@U3n���!?7y��>��@j�9�h�ٿkzl��@Զ��t4@U3n���!?7y��>��@�ϽJ��ٿ�4KI2�@sG��4@狀��!?6~�v1�@�ϽJ��ٿ�4KI2�@sG��4@狀��!?6~�v1�@�ϽJ��ٿ�4KI2�@sG��4@狀��!?6~�v1�@�ϽJ��ٿ�4KI2�@sG��4@狀��!?6~�v1�@�ϽJ��ٿ�4KI2�@sG��4@狀��!?6~�v1�@J���ٿ|���X�@�rk4@i����!?7wL�4�@�P���ٿe����@�cj�4@@q�J�!?�A溠�@�P���ٿe����@�cj�4@@q�J�!?�A溠�@�_���ٿhm�-}�@�	� 4@��G�!?�=���0�@)�ytw�ٿ-�.�e�@B�y� �3@.��W�!?*�=�C��@�	���ٿ�3���@E�$�3@�X�j�!?�!�f�@�	���ٿ�3���@E�$�3@�X�j�!?�!�f�@E ���ٿ�F�O��@?�����3@z�Q�!?@X�ɖ�@E ���ٿ�F�O��@?�����3@z�Q�!?@X�ɖ�@E ���ٿ�F�O��@?�����3@z�Q�!?@X�ɖ�@E ���ٿ�F�O��@?�����3@z�Q�!?@X�ɖ�@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@Ɛ�1�ٿy�&_�@�k� 4@�c��h�!? t���@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@p�.%�ٿe� H#��@�Υ�4@H��ai�!?@��M�@��o�!�ٿzR��rS�@"�	�� 4@�>��!? h"�Vi�@��o�!�ٿzR��rS�@"�	�� 4@�>��!? h"�Vi�@��o�!�ٿzR��rS�@"�	�� 4@�>��!? h"�Vi�@��o�!�ٿzR��rS�@"�	�� 4@�>��!? h"�Vi�@��sS�ٿI�l����@f4mQN4@b�!?�6�)k�@��sS�ٿI�l����@f4mQN4@b�!?�6�)k�@��sS�ٿI�l����@f4mQN4@b�!?�6�)k�@�'d��ٿנ5J4e�@-'}��3@�0�-Ǐ!?KӎY��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@ON{şٿ�|)�ǌ�@�F�	 4@c�;��!?�@�.<��@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@;Y^���ٿTT�`��@���b 4@P�jH��!?�xi��G�@U��ٿ��x���@K���m 4@|�wዏ!?�Ζ���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@t?\�ۦٿ�0Tl��@�U���3@����!?�&���@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@����n�ٿ[��~�@���9�3@�*�x�!?����@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q�5���ٿg1B/�f�@����;�3@T�L�ˏ!?��t��@Q� o7�ٿ]n�F���@��WW��3@p�V��!?=�F:�@Q� o7�ٿ]n�F���@��WW��3@p�V��!?=�F:�@Q� o7�ٿ]n�F���@��WW��3@p�V��!?=�F:�@Q� o7�ٿ]n�F���@��WW��3@p�V��!?=�F:�@�t�ٿ�gj����@WH ~B�3@8�5K�!?��L�0�@�t�ٿ�gj����@WH ~B�3@8�5K�!?��L�0�@�t�ٿ�gj����@WH ~B�3@8�5K�!?��L�0�@ �^��ٿ:L� ��@�/�m4@Ty��z�!?u[C@���@ �^��ٿ:L� ��@�/�m4@Ty��z�!?u[C@���@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@Y���ٿt�T0��@�1�� 4@�&�o�!?���Fys�@�	x�y�ٿ^g����@�M�X 4@����h�!?�Y�u*�@Fc	N�ٿx� ��@W��+j4@������!?-���B�@Fc	N�ٿx� ��@W��+j4@������!?-���B�@v�ٿT��q��@"dD+� 4@��h6��!?:v4�s~�@v�ٿT��q��@"dD+� 4@��h6��!?:v4�s~�@v�ٿT��q��@"dD+� 4@��h6��!?:v4�s~�@v�ٿT��q��@"dD+� 4@��h6��!?:v4�s~�@v�ٿT��q��@"dD+� 4@��h6��!?:v4�s~�@\�!##�ٿ�a����@��J� 4@R��߿�!?�`�c���@\�!##�ٿ�a����@��J� 4@R��߿�!?�`�c���@\�!##�ٿ�a����@��J� 4@R��߿�!?�`�c���@��5ғ�ٿ(�����@VJPz4@�}eY��!?X�g_��@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@"���զٿ�@)�$`�@jR&S4@��c\��!?��>��%�@���ٿ��ɣ�r�@���4@$���`�!?�Nr�@��@���ٿ��ɣ�r�@���4@$���`�!?�Nr�@��@���ٿ��ɣ�r�@���4@$���`�!?�Nr�@��@���ٿ��ɣ�r�@���4@$���`�!?�Nr�@��@���ٿ��ɣ�r�@���4@$���`�!?�Nr�@��@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@�ՔR��ٿ<*�����@�T��4@�����!?�]#B�
�@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@4S����ٿ��h�M�@�J�4@Y�Hŗ�!?�[nav��@s��ٿV!��b�@�~��4@3����!?�^A����@ϖ�ѪٿIx�~>�@�kj;t4@�u܏!?�����@ϖ�ѪٿIx�~>�@�kj;t4@�u܏!?�����@ϖ�ѪٿIx�~>�@�kj;t4@�u܏!?�����@WjrѪٿ�� ��@�K�R4@\�s��!?rז�D��@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�l�j��ٿ�e�I:��@�y��04@�p���!?9�a�̫�@�d@Шٿ|��`��@:��b�4@�=�ϙ�!?}����y�@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@���z�ٿ`cݾ��@H�T�4@�	���!?A�'�.��@�v��ٿ��n%c��@��&4@ՆϏ!?�r�(�M�@�vc[l�ٿ�p�6�S�@b~rV� 4@�/c�a�!?[�)���@�vc[l�ٿ�p�6�S�@b~rV� 4@�/c�a�!?[�)���@�`r�I�ٿ��tl�@�GzD�4@c��0��!?ʔ����@�`r�I�ٿ��tl�@�GzD�4@c��0��!?ʔ����@�`r�I�ٿ��tl�@�GzD�4@c��0��!?ʔ����@�`r�I�ٿ��tl�@�GzD�4@c��0��!?ʔ����@��f�ٿ��sg�j�@���4@�2�b�!?�n~X���@Ô�`�ٿ��?4c��@��
1�4@����!?����T��@Ô�`�ٿ��?4c��@��
1�4@����!?����T��@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@	Qʤ/�ٿnI��1�@X��w�4@T��`�!?�l���@vS2���ٿt3�X���@�]Ǯ14@7�w�!?�w'Y�@vS2���ٿt3�X���@�]Ǯ14@7�w�!?�w'Y�@vS2���ٿt3�X���@�]Ǯ14@7�w�!?�w'Y�@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@0�Фٿ�{��Ƶ�@e%���3@�΋M\�!?�-+� �@�s�|�ٿ<�,R��@C�;� 4@z�Ȧ�!?zd��e�@�p���ٿ3�(�@~(b�r4@Z�����!?飲���@�p���ٿ3�(�@~(b�r4@Z�����!?飲���@�p���ٿ3�(�@~(b�r4@Z�����!?飲���@�J*V�ٿDh9����@�ٚ� 4@��R��!?\���`I�@�J*V�ٿDh9����@�ٚ� 4@��R��!?\���`I�@�J*V�ٿDh9����@�ٚ� 4@��R��!?\���`I�@H��|�ٿ �8��@�Wu�� 4@ϐF1Ϗ!?���ou�@H��|�ٿ �8��@�Wu�� 4@ϐF1Ϗ!?���ou�@�$7p�ٿ/�[v3�@ߑk{ 4@��!?rP��d�@�$7p�ٿ/�[v3�@ߑk{ 4@��!?rP��d�@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@d�쌙ٿ��:�W�@<lwF�3@c.k��!?�H��.��@бxٺ�ٿ� �T�@��d���3@:a�܇�!?�3t���@бxٺ�ٿ� �T�@��d���3@:a�܇�!?�3t���@бxٺ�ٿ� �T�@��d���3@:a�܇�!?�3t���@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@�]j]s�ٿ�d�"��@p�1=4@M.�O�!?�^~�@cJ����ٿH�=�"��@
��4@�~.�>�!?����H�@cJ����ٿH�=�"��@
��4@�~.�>�!?����H�@?�V�ٮٿΩ�t��@R@�4@��×L�!?N�����@?�V�ٮٿΩ�t��@R@�4@��×L�!?N�����@?�V�ٮٿΩ�t��@R@�4@��×L�!?N�����@?�V�ٮٿΩ�t��@R@�4@��×L�!?N�����@?�V�ٮٿΩ�t��@R@�4@��×L�!?N�����@��+-��ٿ��E��
�@���4@޾;)ŏ!?MAܽ��@��+-��ٿ��E��
�@���4@޾;)ŏ!?MAܽ��@�y`��ٿ��.CB�@����4@�����!?�k�@�y`��ٿ��.CB�@����4@�����!?�k�@<��"��ٿ:XX����@)�L74@��V@�!?�m��@��Ԟٿ޵J��4�@TP}�4@!�9L?�!?*oG����@��Ԟٿ޵J��4�@TP}�4@!�9L?�!?*oG����@��Ԟٿ޵J��4�@TP}�4@!�9L?�!?*oG����@4�R���ٿ@=�zZ�@N��FA4@|�Q^�!?^Kq�@4�R���ٿ@=�zZ�@N��FA4@|�Q^�!?^Kq�@4�R���ٿ@=�zZ�@N��FA4@|�Q^�!?^Kq�@Ay���ٿ�lZ�#�@�\1�4@t�E��!??LК���@Ay���ٿ�lZ�#�@�\1�4@t�E��!??LК���@Ay���ٿ�lZ�#�@�\1�4@t�E��!??LК���@�p	���ٿD,�� ��@G�;� 4@uÙ��!?�_*���@�p	���ٿD,�� ��@G�;� 4@uÙ��!?�_*���@�p	���ٿD,�� ��@G�;� 4@uÙ��!?�_*���@�;
�k�ٿ(c�L��@ �`��4@W�D&��!?R��L��@�;
�k�ٿ(c�L��@ �`��4@W�D&��!?R��L��@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@'�0��ٿj�d����@�E��4@���S��!?ꚗBEN�@���)�ٿ� �t��@<n�
E 4@6���!?�8���@�:m��ٿ �5vu��@��0�}4@�p���!?�S�����@�:m��ٿ �5vu��@��0�}4@�p���!?�S�����@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@��ߤ�ٿ�`ߏ�@��l���3@����ޏ!?Ŏ�L�j�@���q��ٿ���.>�@%�Oc 4@�G�C�!?
�xq<�@���q��ٿ���.>�@%�Oc 4@�G�C�!?
�xq<�@� �!��ٿhr�ʠ	�@���3@5�]�	�!?,_K�8}�@� �!��ٿhr�ʠ	�@���3@5�]�	�!?,_K�8}�@� �!��ٿhr�ʠ	�@���3@5�]�	�!?,_K�8}�@|��Bo�ٿ�{0�Bk�@ު�( 4@p��#��!?���:c��@|��Bo�ٿ�{0�Bk�@ު�( 4@p��#��!?���:c��@�ݸH}�ٿĐ��U��@�uB��3@ g��f�!?��]����@�����ٿ����@ D��3@�^���!?&��셹�@�����ٿ����@ D��3@�^���!?&��셹�@�����ٿ����@ D��3@�^���!?&��셹�@�����ٿ����@ D��3@�^���!?&��셹�@�����ٿ����@ D��3@�^���!?&��셹�@�b�}ƣٿ
����@	�n~6�3@� �Wt�!?���F�A�@�b�}ƣٿ
����@	�n~6�3@� �Wt�!?���F�A�@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@�8��ٿ��
�5��@{��i 4@���t}�!?BNm�?��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@��IΜ�ٿ�1`2�j�@�f� 4@�ɽ+~�!?�<ut��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@j޼B_�ٿ�-���@���H��3@h�7�i�!?9�{&}��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@��! F�ٿ{��k��@\F��t�3@}����!?���YZ��@�����ٿ�0�M�8�@f�u
� 4@�3�Y��!?�%7�[�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�����ٿ`�_>�@��q 4@]��=�!?K	�	�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@�y �ٿ��5����@S���j�3@a�=-l�!?�ҧ�h)�@q^J߿�ٿ`���:��@��=i�3@�J���!?`���P��@q^J߿�ٿ`���:��@��=i�3@�J���!?`���P��@ￂ_�ٿ��Z��@���b�3@�����!?!��� |�@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@Z��u�ٿF�v�@��2�^4@��}媏!?r�b��@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@�1����ٿM"���v�@$�`��4@�8 ���!?Y�<Ѝ�@`��ȩٿg��<��@C/ K�4@G�BY�!?YCm���@��kʨٿ��J֏��@��4@B_����!?�[�j)�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@FԤ��ٿk\ ��d�@{φ�H4@?09"��!?��˞t>�@��J���ٿr縫l��@�j�4@#'���!?4���z�@��J���ٿr縫l��@�j�4@#'���!?4���z�@��J���ٿr縫l��@�j�4@#'���!?4���z�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@~\NVҫٿN��x��@�g��4@����؏!?�Z�|-�@D���I�ٿҶ\�@+"�+�4@�����!?6Ï&8j�@D���I�ٿҶ\�@+"�+�4@�����!?6Ï&8j�@D���I�ٿҶ\�@+"�+�4@�����!?6Ï&8j�@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@$�F�{�ٿz
d�e��@��=�q4@�$E�Ώ!?�F���@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@Y��Ƈ�ٿ`�_d/��@�� 4@�w{ɱ�!?�H�,��@u&N��ٿU���om�@�I(�p4@g�Ƀ�!?<vs~̩�@u&N��ٿU���om�@�I(�p4@g�Ƀ�!?<vs~̩�@u&N��ٿU���om�@�I(�p4@g�Ƀ�!?<vs~̩�@��Q��ٿ&QL�Z��@�`-	P4@� l�!?�]����@��Q��ٿ&QL�Z��@�`-	P4@� l�!?�]����@��Q��ٿ&QL�Z��@�`-	P4@� l�!?�]����@��Q��ٿ&QL�Z��@�`-	P4@� l�!?�]����@���X�ٿA�L����@Mj�w4@�d����!?�?��4��@���X�ٿA�L����@Mj�w4@�d����!?�?��4��@���X�ٿA�L����@Mj�w4@�d����!?�?��4��@���M��ٿX�e���@B<� 4@i���!?�9_��@���M��ٿX�e���@B<� 4@i���!?�9_��@���M��ٿX�e���@B<� 4@i���!?�9_��@���M��ٿX�e���@B<� 4@i���!?�9_��@���M��ٿX�e���@B<� 4@i���!?�9_��@���M��ٿX�e���@B<� 4@i���!?�9_��@�X3^�ٿ�E�����@�P�V8 4@cu�Q�!?3R��"�@�X3^�ٿ�E�����@�P�V8 4@cu�Q�!?3R��"�@N�{M�ٿ.�4\y*�@��=��4@�B6��!?(O�@��_�ٿ��	����@vĥN@4@oy7�!?|��oR�@A����ٿ+^*�i��@���k4@�
�J�!?�'�7;��@A����ٿ+^*�i��@���k4@�
�J�!?�'�7;��@\��ϗٿ세�h�@"(`&4@]��qg�!?�������@��)�k�ٿB�:���@<��@z 4@�h;nA�!?§��@��)�k�ٿB�:���@<��@z 4@�h;nA�!?§��@��)�k�ٿB�:���@<��@z 4@�h;nA�!?§��@��)�k�ٿB�:���@<��@z 4@�h;nA�!?§��@pTk{E�ٿ��Ħ�@NNJ4@��=��!?b�f�@pTk{E�ٿ��Ħ�@NNJ4@��=��!?b�f�@pTk{E�ٿ��Ħ�@NNJ4@��=��!?b�f�@pTk{E�ٿ��Ħ�@NNJ4@��=��!?b�f�@pTk{E�ٿ��Ħ�@NNJ4@��=��!?b�f�@���䂣ٿ��d��(�@���4@�53���!?d���!��@���䂣ٿ��d��(�@���4@�53���!?d���!��@sh�ٿZ0#~�@z�A�4@�0>��!?�yT��@sh�ٿZ0#~�@z�A�4@�0>��!?�yT��@sh�ٿZ0#~�@z�A�4@�0>��!?�yT��@sh�ٿZ0#~�@z�A�4@�0>��!?�yT��@sh�ٿZ0#~�@z�A�4@�0>��!?�yT��@M}]x�ٿ)��L���@b6�@��3@K��"v�!?e�I�C�@M}]x�ٿ)��L���@b6�@��3@K��"v�!?e�I�C�@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@J<��ٿ�\� �@��c��3@��?f�!?��[����@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@�#Yv�ٿ9�.���@�'[@= 4@M=;�k�!?�(���@��Ӵ>�ٿ��W�r�@�1���4@�u\�r�!?�(�'o+�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@M�D5�ٿ�v�����@7���(4@H���A�!?�2��}^�@Z+��ٿ��A-�@��{a4@K[�)�!?�]�d��@1��@�ٿMik	҈�@�<V�#�3@i1qy�!?�]�����@t>H�ٿiY؎9S�@�}���3@��J�!?�<��1K�@t>H�ٿiY؎9S�@�}���3@��J�!?�<��1K�@t>H�ٿiY؎9S�@�}���3@��J�!?�<��1K�@t>H�ٿiY؎9S�@�}���3@��J�!?�<��1K�@t>H�ٿiY؎9S�@�}���3@��J�!?�<��1K�@p���ٿ����@.~����3@EF�x�!?/�Q��@p���ٿ����@.~����3@EF�x�!?/�Q��@p���ٿ����@.~����3@EF�x�!?/�Q��@�
��ٿ+U��B��@&
�=��3@_�b���!?3���e�@�
��ٿ+U��B��@&
�=��3@_�b���!?3���e�@����6�ٿ�aF��@�_"�5�3@����!?M�m�׷�@�Fg��ٿh��iF��@V�ܲ�3@�C]��!?�����@�Fg��ٿh��iF��@V�ܲ�3@�C]��!?�����@���Y�ٿ���� �@9�y� �3@(�@X�!?�;� @S�@���Y�ٿ���� �@9�y� �3@(�@X�!?�;� @S�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@b9Kr�ٿ��oDzt�@_��S4@���o�!?^�\�>�@���*�ٿ��pK��@s0�Q(4@&�B�!?X�`�	~�@���*�ٿ��pK��@s0�Q(4@&�B�!?X�`�	~�@���*�ٿ��pK��@s0�Q(4@&�B�!?X�`�	~�@���*�ٿ��pK��@s0�Q(4@&�B�!?X�`�	~�@��H��ٿ�������@_u$$A4@I�_-�!?�q��'T�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��_尳ٿc��0��@'ޖ�� 4@	_����!?:L5�3�@��2G�ٿ�jg=z�@�^�]�4@����Ϗ!?�j_���@��2G�ٿ�jg=z�@�^�]�4@����Ϗ!?�j_���@��2G�ٿ�jg=z�@�^�]�4@����Ϗ!?�j_���@��2G�ٿ�jg=z�@�^�]�4@����Ϗ!?�j_���@�^M�E�ٿ�FS���@�TK� 4@�f�;D�!?Ԫ����@�^M�E�ٿ�FS���@�TK� 4@�f�;D�!?Ԫ����@�^M�E�ٿ�FS���@�TK� 4@�f�;D�!?Ԫ����@�^M�E�ٿ�FS���@�TK� 4@�f�;D�!?Ԫ����@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@@ҢY٫ٿ��㗛8�@!�1Q��3@�0���!?���@�Hԫٿ��Y�є�@���	��3@�{M�!?ʎ��0]�@�:9�U�ٿ������@��`W4@Eڳ�ۏ!?�ݳz}�@�:9�U�ٿ������@��`W4@Eڳ�ۏ!?�ݳz}�@�:9�U�ٿ������@��`W4@Eڳ�ۏ!?�ݳz}�@�:9�U�ٿ������@��`W4@Eڳ�ۏ!?�ݳz}�@���!A�ٿ���o�J�@�@��m4@!s�ď!?]\Cn��@���!A�ٿ���o�J�@�@��m4@!s�ď!?]\Cn��@yL����ٿ�=F_�@x�r�, 4@*&�`Ǐ!?t�l�L��@yL����ٿ�=F_�@x�r�, 4@*&�`Ǐ!?t�l�L��@yL����ٿ�=F_�@x�r�, 4@*&�`Ǐ!?t�l�L��@�]�ٿ=f��L��@����R 4@�7�#̏!?�:k�B��@�]�ٿ=f��L��@����R 4@�7�#̏!?�:k�B��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@H��>�ٿw���Ƅ�@����� 4@������!?��Cs\��@_��t�ٿΛ�S^��@G���4@�b鞏!?������@_��t�ٿΛ�S^��@G���4@�b鞏!?������@_��t�ٿΛ�S^��@G���4@�b鞏!?������@_��t�ٿΛ�S^��@G���4@�b鞏!?������@_��t�ٿΛ�S^��@G���4@�b鞏!?������@_��t�ٿΛ�S^��@G���4@�b鞏!?������@þ��ٿ��Ic;�@��ǅg4@�V?���!?f-��@þ��ٿ��Ic;�@��ǅg4@�V?���!?f-��@þ��ٿ��Ic;�@��ǅg4@�V?���!?f-��@þ��ٿ��Ic;�@��ǅg4@�V?���!?f-��@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@��Ɯٿ��wy�@���i 4@�����!?:��=�@�VĂ��ٿ����{�@ ����4@%]�1��!?7!��L��@�VĂ��ٿ����{�@ ����4@%]�1��!?7!��L��@��P�ٿ�%qʼ^�@q�\.t4@W�$r�!?�1��@��P�ٿ�%qʼ^�@q�\.t4@W�$r�!?�1��@��P�ٿ�%qʼ^�@q�\.t4@W�$r�!?�1��@��P�ٿ�%qʼ^�@q�\.t4@W�$r�!?�1��@��P�ٿ�%qʼ^�@q�\.t4@W�$r�!?�1��@dBǳ��ٿ�]��d�@b+�� 4@`�G���!?@Y/P��@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@��'��ٿgB�i%3�@����)4@q,�~�!?������@~]�F��ٿz#�Q���@���:4@�-)���!?v��Ŕ��@~]�F��ٿz#�Q���@���:4@�-)���!?v��Ŕ��@~]�F��ٿz#�Q���@���:4@�-)���!?v��Ŕ��@~]�F��ٿz#�Q���@���:4@�-)���!?v��Ŕ��@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@_W�=�ٿqyZ$�Q�@@[�(�3@?��|�!?5[s����@?QA��ٿu9�+�@��0��3@)s���!?�{2���@?QA��ٿu9�+�@��0��3@)s���!?�{2���@�G?ԝٿm����(�@�E�3@���l��!?L���h��@j�Yj�ٿ0)�<<4�@�LA��3@G.�ѳ�!?��ܡ�g�@j�Yj�ٿ0)�<<4�@�LA��3@G.�ѳ�!?��ܡ�g�@j�Yj�ٿ0)�<<4�@�LA��3@G.�ѳ�!?��ܡ�g�@j�Yj�ٿ0)�<<4�@�LA��3@G.�ѳ�!?��ܡ�g�@j�v���ٿ�z�x�@�����3@xj��!?���WH��@b�����ٿ�n��@G�xR4@$��!?U©S%�@b�����ٿ�n��@G�xR4@$��!?U©S%�@b�����ٿ�n��@G�xR4@$��!?U©S%�@b�����ٿ�n��@G�xR4@$��!?U©S%�@b�����ٿ�n��@G�xR4@$��!?U©S%�@b�����ٿ�n��@G�xR4@$��!?U©S%�@�C�M��ٿ��1�>��@0����3@F��ӏ!?q�����@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�����ٿ/�����@<�s���3@` ����!?�`eM��@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@�&cx��ٿ�؏�A�@ɉ�� 4@Q�o���!?NR�U���@o(����ٿ�E)<�"�@�];3��3@�C���!?sB�m1?�@o(����ٿ�E)<�"�@�];3��3@�C���!?sB�m1?�@o(����ٿ�E)<�"�@�];3��3@�C���!?sB�m1?�@o(����ٿ�E)<�"�@�];3��3@�C���!?sB�m1?�@o(����ٿ�E)<�"�@�];3��3@�C���!?sB�m1?�@��ܨL�ٿ��o��@�+�b�4@N0L���!?\�$���@��ܨL�ٿ��o��@�+�b�4@N0L���!?\�$���@��ܨL�ٿ��o��@�+�b�4@N0L���!?\�$���@��ܨL�ٿ��o��@�+�b�4@N0L���!?\�$���@=�d���ٿT/�T�@���b� 4@�پIM�!?�o&�Y��@=�d���ٿT/�T�@���b� 4@�پIM�!?�o&�Y��@=�d���ٿT/�T�@���b� 4@�پIM�!?�o&�Y��@=�d���ٿT/�T�@���b� 4@�پIM�!?�o&�Y��@=�d���ٿT/�T�@���b� 4@�پIM�!?�o&�Y��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@�w����ٿ�������@)��,� 4@��w��!?�(;��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@*Q�5b�ٿ"0ڑ��@���4@�+���!?���.I��@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@n��h>�ٿĥ��˖�@��
�� 4@mh8���!?q|�nf�@yٳy�ٿ]�J����@;kp� 4@"�ED��!?��U��@yٳy�ٿ]�J����@;kp� 4@"�ED��!?��U��@yٳy�ٿ]�J����@;kp� 4@"�ED��!?��U��@yٳy�ٿ]�J����@;kp� 4@"�ED��!?��U��@yٳy�ٿ]�J����@;kp� 4@"�ED��!?��U��@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@S�,i�ٿm1ްm�@����3@m�쾥�!?��9�Z�@H�0H�ٿh�ۂ��@���� 4@s��a��!?6FN�X��@H�0H�ٿh�ۂ��@���� 4@s��a��!?6FN�X��@ �J4��ٿ��a'z��@��ݛ 4@3搾N�!?[0�ԛ��@:}Z��ٿ~�=�s�@���D�4@R�R[�!?����@�K���ٿB������@��
%+4@B �/��!?�=�α��@�K���ٿB������@��
%+4@B �/��!?�=�α��@�K���ٿB������@��
%+4@B �/��!?�=�α��@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@fi�^��ٿ#��8\��@���� 4@�0QF�!?�Yv�}�@?i�Ú�ٿEy��n|�@#Nu�� 4@7̉Kk�!?"r4�@?i�Ú�ٿEy��n|�@#Nu�� 4@7̉Kk�!?"r4�@?i�Ú�ٿEy��n|�@#Nu�� 4@7̉Kk�!?"r4�@?i�Ú�ٿEy��n|�@#Nu�� 4@7̉Kk�!?"r4�@���Ƹ�ٿ�����@Xd�7 4@9�h8��!?�Q#�M�@���Ƹ�ٿ�����@Xd�7 4@9�h8��!?�Q#�M�@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@���Ok�ٿ6+-X:��@?�+ 4@��?��!?J���`��@-�� ��ٿ@Տ���@���]4@�X�6��!?���*
��@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@��,`�ٿ��7bt��@���4@�f�ԏ!?�c��A�@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@6��܃�ٿ�x�SB7�@]���4@Z�Cُ!?��'�K��@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@?�L�q�ٿͧEŤ�@��A�4@�����!?��|�m�@����ןٿi�c�N	�@đ�t 4@y��׏!?N�h��3�@����ןٿi�c�N	�@đ�t 4@y��׏!?N�h��3�@����ןٿi�c�N	�@đ�t 4@y��׏!?N�h��3�@����ןٿi�c�N	�@đ�t 4@y��׏!?N�h��3�@j�W��ٿB�8Kq��@:�L4@�4���!?{��aT�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@Z<R*�ٿ�e;��@;@��54@�ɊH��!?���/�@�$�Kנٿ^N�kMP�@'70��4@t�ޚ�!?�B�FL��@�$�Kנٿ^N�kMP�@'70��4@t�ޚ�!?�B�FL��@�$�Kנٿ^N�kMP�@'70��4@t�ޚ�!?�B�FL��@٦5�3�ٿv���]�@UoP
 4@%
��ӏ!?
l��|�@��|���ٿ��*o.�@��=�( 4@�M�ត!?��_���@��ɜٿ��k@��@�Tks4@a& ��!?��0�\��@��ɜٿ��k@��@�Tks4@a& ��!?��0�\��@��ɜٿ��k@��@�Tks4@a& ��!?��0�\��@��ɜٿ��k@��@�Tks4@a& ��!?��0�\��@�v=@�ٿ�L�����@���:4@������!?]20�Q��@�v=@�ٿ�L�����@���:4@������!?]20�Q��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�	��a�ٿ� ���@���t� 4@T����!?)��m��@�v�ٿ]��O��@[����3@,�����!?j�Z���@�v�ٿ]��O��@[����3@,�����!?j�Z���@�6����ٿGϐcĉ�@ׯG;m�3@D!����!?`�q2u��@k��:��ٿ���k��@V�,���3@o%mُ!?Q������@k��:��ٿ���k��@V�,���3@o%mُ!?Q������@k��:��ٿ���k��@V�,���3@o%mُ!?Q������@k��:��ٿ���k��@V�,���3@o%mُ!?Q������@k��:��ٿ���k��@V�,���3@o%mُ!?Q������@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@0���ٿJoӁq��@�({�& 4@C�
Թ�!?��+���@�D(�X�ٿ�K���@�b�6�3@v��
Ϗ!?-1i��@�D(�X�ٿ�K���@�b�6�3@v��
Ϗ!?-1i��@�D(�X�ٿ�K���@�b�6�3@v��
Ϗ!?-1i��@�D(�X�ٿ�K���@�b�6�3@v��
Ϗ!?-1i��@���R1�ٿ�k �/��@*�����3@&����!?�ڰ�k�@���R1�ٿ�k �/��@*�����3@&����!?�ڰ�k�@���R1�ٿ�k �/��@*�����3@&����!?�ڰ�k�@���R1�ٿ�k �/��@*�����3@&����!?�ڰ�k�@��ٿ'�Cj�@Rђ2G�3@������!?./�O��@�;���ٿձc���@�kD�O�3@PW���!?Ų�#|�@�;���ٿձc���@�kD�O�3@PW���!?Ų�#|�@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��r�ٿ��b��X�@�s%?c4@�re͟�!?e�����@��u���ٿg�G�_��@�υ�4@��w��!?�̔�@��u���ٿg�G�_��@�υ�4@��w��!?�̔�@��u���ٿg�G�_��@�υ�4@��w��!?�̔�@��u���ٿg�G�_��@�υ�4@��w��!?�̔�@��u���ٿg�G�_��@�υ�4@��w��!?�̔�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@n��`ìٿ�\�p���@a�w�O�3@:i�j��!?7a��F�@��>���ٿeJ�ԙ�@�Fn���3@	|彏!?̤��g�@��>���ٿeJ�ԙ�@�Fn���3@	|彏!?̤��g�@�L|�ٿ�l�&5��@bK�g��3@|0�5��!?J%����@�L|�ٿ�l�&5��@bK�g��3@|0�5��!?J%����@�L|�ٿ�l�&5��@bK�g��3@|0�5��!?J%����@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@=���H�ٿwƦ&��@���O�3@����!?=�Adi_�@<䫯�ٿ��y
��@�� 4@���[��!?������@<䫯�ٿ��y
��@�� 4@���[��!?������@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@8�4˯ٿi䭑��@�Ԛ��3@����!?
�*5��@���ٿ��j5���@8��y��3@�Nҙ��!?O��X��@���ٿ��j5���@8��y��3@�Nҙ��!?O��X��@���ٿ��j5���@8��y��3@�Nҙ��!?O��X��@C]m���ٿ��t$��@t��u0 4@�&��!?��S �@C]m���ٿ��t$��@t��u0 4@�&��!?��S �@�]��ٿ��QQ��@W��� 4@��(a��!?�a��*?�@�]��ٿ��QQ��@W��� 4@��(a��!?�a��*?�@Ћp�p�ٿ�B"���@K��!4@��*��!?�X@���@Ћp�p�ٿ�B"���@K��!4@��*��!?�X@���@Ћp�p�ٿ�B"���@K��!4@��*��!?�X@���@Ћp�p�ٿ�B"���@K��!4@��*��!?�X@���@Ћp�p�ٿ�B"���@K��!4@��*��!?�X@���@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@� +��ٿ��>ιX�@���`�3@�´��!?���ς�@/Qը�ٿ��[�L[�@Y�� 4@�M]"n�!?��>�g�@�RR�ٿno "=�@D�I;�4@U�eAt�!?".J#O��@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@��5V�ٿ���+�u�@#,�U4@t7e뺏!?`��r���@v�xS�ٿ+���lp�@%õ-)4@�6Q
�!?J�f���@v�xS�ٿ+���lp�@%õ-)4@�6Q
�!?J�f���@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@n��� �ٿ��&�.�@Mw�j� 4@t�=���!?���d�@��A�[�ٿ2������@�-�\�4@�,ꝝ�!?6����@��A�[�ٿ2������@�-�\�4@�,ꝝ�!?6����@��A�[�ٿ2������@�-�\�4@�,ꝝ�!?6����@��A�[�ٿ2������@�-�\�4@�,ꝝ�!?6����@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@:�k��ٿ`� S��@�bV�I4@�Ea�!?{|}��(�@9`_W�ٿ!m�:�@�0NJ�4@,�N��!?`i����@9`_W�ٿ!m�:�@�0NJ�4@,�N��!?`i����@�q��}�ٿ���G�@OےK4@�kT��!?���\��@�q��}�ٿ���G�@OےK4@�kT��!?���\��@�����ٿ��:��@�w"D&4@�p����!?�:��&��@��A��ٿ�E�$�@����4@��G~�!?v� i��@���Z�ٿ���=��@a-�m4@M�	�!?������@��w�ٿ%�EQ���@����3@���@�!?%ꔁ*�@��w�ٿ%�EQ���@����3@���@�!?%ꔁ*�@�Q땬ٿ]�~?��@i��� 4@��ӏ!?�J�
K��@�Q땬ٿ]�~?��@i��� 4@��ӏ!?�J�
K��@�Q땬ٿ]�~?��@i��� 4@��ӏ!?�J�
K��@�Q땬ٿ]�~?��@i��� 4@��ӏ!?�J�
K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�mBi��ٿ������@d�F 4@R��n�!?�d��K��@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@�(���ٿ�qǻ�D�@���>4@>�L��!?Ֆe�ĺ�@��E�ٿ���L�'�@e>�ؿ�3@8%o��!?�\��S��@��E�ٿ���L�'�@e>�ؿ�3@8%o��!?�\��S��@��E�ٿ���L�'�@e>�ؿ�3@8%o��!?�\��S��@��E�ٿ���L�'�@e>�ؿ�3@8%o��!?�\��S��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@*~ϥa�ٿ�~m��7�@ӗ58 4@��縷�!?��\i��@��&��ٿ%��v�*�@@
V[4@����!?PuOE���@��&��ٿ%��v�*�@@
V[4@����!?PuOE���@��&��ٿ%��v�*�@@
V[4@����!?PuOE���@������ٿS��V/�@��v.�4@�^K:r�!?����w�@0\�:Z�ٿ'�X-1�@�3�d: 4@y�2C^�!?�c�xU��@0\�:Z�ٿ'�X-1�@�3�d: 4@y�2C^�!?�c�xU��@0\�:Z�ٿ'�X-1�@�3�d: 4@y�2C^�!?�c�xU��@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@"�xKU�ٿ��:�+��@{�r4@6�5y|�!?�~ ���@uQ_]Мٿ�~Y���@�+NJ�4@��dX�!?�멅���@uQ_]Мٿ�~Y���@�+NJ�4@��dX�!?�멅���@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@�ľc[�ٿ�k��e��@�Z[�24@P��벏!?�L����@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���h�ٿ���a&�@�cŊ 4@S\�bΏ!?�
��m�@���=�ٿ�)��@�hDȓ�3@�]D=�!?[N���L�@���=�ٿ�)��@�hDȓ�3@�]D=�!?[N���L�@��M�~�ٿw@.�7��@�q)���3@c1�uҏ!?��|h�D�@��M�~�ٿw@.�7��@�q)���3@c1�uҏ!?��|h�D�@��M�~�ٿw@.�7��@�q)���3@c1�uҏ!?��|h�D�@8e��j�ٿ}��T0F�@�'O 4@j���!?����0��@8e��j�ٿ}��T0F�@�'O 4@j���!?����0��@8e��j�ٿ}��T0F�@�'O 4@j���!?����0��@8e��j�ٿ}��T0F�@�'O 4@j���!?����0��@	�k��ٿد4��K�@�K���4@s]�W�!?s7G�d�@���t�ٿ}��vb!�@��z��3@����k�!?
H���@���t�ٿ}��vb!�@��z��3@����k�!?
H���@���t�ٿ}��vb!�@��z��3@����k�!?
H���@���t�ٿ}��vb!�@��z��3@����k�!?
H���@�볘ٿT ��{��@'w���3@P1�;��!?"
�Ƚ�@�볘ٿT ��{��@'w���3@P1�;��!?"
�Ƚ�@��!\6�ٿ=��ԛd�@|�0;`�3@�fR׽�!?EAq��@��!\6�ٿ=��ԛd�@|�0;`�3@�fR׽�!?EAq��@��!\6�ٿ=��ԛd�@|�0;`�3@�fR׽�!?EAq��@��!\6�ٿ=��ԛd�@|�0;`�3@�fR׽�!?EAq��@`d�R
�ٿ'p��@�tT�4@}8|Ϣ�!?H�=��<�@C���Цٿg��ʗ�@�*��� 4@����J�!?ɣ�}���@C���Цٿg��ʗ�@�*��� 4@����J�!?ɣ�}���@C���Цٿg��ʗ�@�*��� 4@����J�!?ɣ�}���@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@J�#���ٿ�u�ޱ�@�$���4@��vy�!?��8q)��@){��z�ٿ�Ò��@��� 4@z��[�!?L�f'���@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@�>���ٿtԍ��S�@D�=�� 4@e�2̜�!?��F��@����ٿN1֯`�@��+ 4@M�ɷ�!?���1�k�@����ٿN1֯`�@��+ 4@M�ɷ�!?���1�k�@����ٿN1֯`�@��+ 4@M�ɷ�!?���1�k�@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@�gŧٿG�D�9�@r�����3@X�����!?	������@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@0n�+e�ٿ�1�s��@'8|� 4@Bx\H^�!?o����@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@TS�Co�ٿ�b����@�Il4@g� |�!?Y�n���@f�n��ٿ�����@�տ4@1���~�!?+����I�@f�n��ٿ�����@�տ4@1���~�!?+����I�@f�n��ٿ�����@�տ4@1���~�!?+����I�@f�n��ٿ�����@�տ4@1���~�!?+����I�@o�6ԭٿ�mx��@E�O� 4@�\4���!?�Ȕfe�@o�6ԭٿ�mx��@E�O� 4@�\4���!?�Ȕfe�@o�6ԭٿ�mx��@E�O� 4@�\4���!?�Ȕfe�@���I�ٿ�����f�@��[\9 4@�V<Mޏ!?D@v"�@���I�ٿ�����f�@��[\9 4@�V<Mޏ!?D@v"�@���I�ٿ�����f�@��[\9 4@�V<Mޏ!?D@v"�@���I�ٿ�����f�@��[\9 4@�V<Mޏ!?D@v"�@���I�ٿ�����f�@��[\9 4@�V<Mޏ!?D@v"�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�6�;ĥٿi�L*(��@8oc1* 4@V� �!?�p���,�@�@>b�ٿ}���c~�@$7	�3@�<�ߏ!?dc�`z�@�@>b�ٿ}���c~�@$7	�3@�<�ߏ!?dc�`z�@U�z�Οٿ�*���e�@�gԚ4@�.��!?=R����@U�z�Οٿ�*���e�@�gԚ4@�.��!?=R����@U�z�Οٿ�*���e�@�gԚ4@�.��!?=R����@�tYa�ٿSEX�@PA-�4@��k���!??��"I��@�tYa�ٿSEX�@PA-�4@��k���!??��"I��@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@<Y��؞ٿ�2�Z��@�ŗQ�3@o>�H��!?}��|���@1%��	�ٿ��a�A��@��94@b�^�!?���r�@1%��	�ٿ��a�A��@��94@b�^�!?���r�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@?�֥�ٿZYc��@�.`4@�ǝ���!?
��\�@ޖ�ߛ�ٿM7���i�@�S�C(4@�^�ڛ�!?%1hG&[�@ޖ�ߛ�ٿM7���i�@�S�C(4@�^�ڛ�!?%1hG&[�@ޖ�ߛ�ٿM7���i�@�S�C(4@�^�ڛ�!?%1hG&[�@ũ4B�ٿ��̆��@��a�e 4@(|��!?X��u�J�@ũ4B�ٿ��̆��@��a�e 4@(|��!?X��u�J�@x��쑥ٿC; &5S�@?���� 4@�au��!?�Kh�f��@x��쑥ٿC; &5S�@?���� 4@�au��!?�Kh�f��@�_l�e�ٿCi�y{�@/���4@^2��!?�ȍ՝�@
����ٿ�
h�#��@QBipZ 4@(�����!?�Z3�T�@
����ٿ�
h�#��@QBipZ 4@(�����!?�Z3�T�@
����ٿ�
h�#��@QBipZ 4@(�����!?�Z3�T�@��/��ٿ�-J�gX�@�u}�}4@Y!/@�!?e����@��/��ٿ�-J�gX�@�u}�}4@Y!/@�!?e����@��/��ٿ�-J�gX�@�u}�}4@Y!/@�!?e����@��/��ٿ�-J�gX�@�u}�}4@Y!/@�!?e����@Gr�û�ٿP���`�@��s/�4@σϏ!??v��lf�@Gr�û�ٿP���`�@��s/�4@σϏ!??v��lf�@Gr�û�ٿP���`�@��s/�4@σϏ!??v��lf�@Gr�û�ٿP���`�@��s/�4@σϏ!??v��lf�@��3�ٿ���-j��@�{�@4@�G)��!?��١��@��3�ٿ���-j��@�{�@4@�G)��!?��١��@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@?��'�ٿ�K��)�@�xдH 4@Au����!?^�O{J�@m�GN�ٿC�a��z�@�i��}�3@y�����!?���	R��@m�GN�ٿC�a��z�@�i��}�3@y�����!?���	R��@m�GN�ٿC�a��z�@�i��}�3@y�����!?���	R��@m�GN�ٿC�a��z�@�i��}�3@y�����!?���	R��@�$M��ٿ�Q�@Ɖ�@��?��3@�J�ʌ�!?�l���@�$M��ٿ�Q�@Ɖ�@��?��3@�J�ʌ�!?�l���@:7 ΅�ٿ�x���@�m���3@��H��!?޲����@:7 ΅�ٿ�x���@�m���3@��H��!?޲����@�5��֖ٿ�3����@'�����3@�� 0�!?rC�>�-�@�5��֖ٿ�3����@'�����3@�� 0�!?rC�>�-�@�5��֖ٿ�3����@'�����3@�� 0�!?rC�>�-�@�5��֖ٿ�3����@'�����3@�� 0�!?rC�>�-�@�0.�ٿ¢�J=7�@��dZ 4@��m���!?v�#T��@�0.�ٿ¢�J=7�@��dZ 4@��m���!?v�#T��@�+@�ٿY\�����@od�t�4@��Z%w�!?q_n���@�+@�ٿY\�����@od�t�4@��Z%w�!?q_n���@�+@�ٿY\�����@od�t�4@��Z%w�!?q_n���@�+@�ٿY\�����@od�t�4@��Z%w�!?q_n���@sM/�ٿu�h��@���e 4@Aʝe��!?�)�X��@sM/�ٿu�h��@���e 4@Aʝe��!?�)�X��@9�.�x�ٿƭ����@?e��4@
����!?s�[ߥ�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@,�q��ٿ�[\ę��@��4@�l�Ъ�!?Ʌ^�_�@�<t;�ٿ�`�V���@0�J� 4@��ݝݏ!?C�̿�C�@�<t;�ٿ�`�V���@0�J� 4@��ݝݏ!?C�̿�C�@�<t;�ٿ�`�V���@0�J� 4@��ݝݏ!?C�̿�C�@�<t;�ٿ�`�V���@0�J� 4@��ݝݏ!?C�̿�C�@�<t;�ٿ�`�V���@0�J� 4@��ݝݏ!?C�̿�C�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@�C���ٿ�-�Ť�@�L�[�3@��,���!?��c��j�@ȓ��ٿy `�@/	k���3@����!?1gi���@ȓ��ٿy `�@/	k���3@����!?1gi���@ȓ��ٿy `�@/	k���3@����!?1gi���@ȓ��ٿy `�@/	k���3@����!?1gi���@ȓ��ٿy `�@/	k���3@����!?1gi���@u�ԮI�ٿ�����@S����3@bK����!?�ڿ���@u�ԮI�ٿ�����@S����3@bK����!?�ڿ���@u�ԮI�ٿ�����@S����3@bK����!?�ڿ���@u�ԮI�ٿ�����@S����3@bK����!?�ڿ���@/[r��ٿ���D��@Ñ��M4@@oL:��!?�4!`��@/[r��ٿ���D��@Ñ��M4@@oL:��!?�4!`��@/[r��ٿ���D��@Ñ��M4@@oL:��!?�4!`��@/[r��ٿ���D��@Ñ��M4@@oL:��!?�4!`��@/[r��ٿ���D��@Ñ��M4@@oL:��!?�4!`��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@���(��ٿv��(���@Q�O�4@3�3K��!?����_��@~��9�ٿ����_'�@�B�14@�]|�!?���A�K�@~��9�ٿ����_'�@�B�14@�]|�!?���A�K�@~��9�ٿ����_'�@�B�14@�]|�!?���A�K�@~��9�ٿ����_'�@�B�14@�]|�!?���A�K�@~��9�ٿ����_'�@�B�14@�]|�!?���A�K�@կ����ٿ;.�O��@�6JK4@��T�!?պu�S��@կ����ٿ;.�O��@�6JK4@��T�!?պu�S��@կ����ٿ;.�O��@�6JK4@��T�!?պu�S��@��a\��ٿN�(��@���� 4@�$M���!?a������@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@���Q#�ٿ�
ѹ�^�@P>y��4@�-.#ď!?G�h�@	�q9��ٿ�57���@��ܳ�4@����!?�ЬP���@�ӫ�v�ٿ�"��o��@�
H��4@�3�ď!?�7���@�ӫ�v�ٿ�"��o��@�
H��4@�3�ď!?�7���@�ӫ�v�ٿ�"��o��@�
H��4@�3�ď!?�7���@")	��ٿgq,K �@�`���4@nc�nǏ!?���Y��@ڍu��ٿr���@���dC 4@�v"3��!?��q�%)�@�(�7�ٿ�@M�ِ�@]W��4@��ɬ�!?�}�K�@�(�7�ٿ�@M�ِ�@]W��4@��ɬ�!?�}�K�@�(�7�ٿ�@M�ِ�@]W��4@��ɬ�!?�}�K�@�(�7�ٿ�@M�ِ�@]W��4@��ɬ�!?�}�K�@��.���ٿ���b�@�C�r4@~wɌz�!?���ִ}�@��.���ٿ���b�@�C�r4@~wɌz�!?���ִ}�@j!?c�ٿ�������@c���<4@��9K�!?���u�E�@j!?c�ٿ�������@c���<4@��9K�!?���u�E�@=���2�ٿ�Y�R��@��ڏ4@B�fMP�!?�Gu0Q�@=���2�ٿ�Y�R��@��ڏ4@B�fMP�!?�Gu0Q�@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@0��x��ٿ�FbUY�@����4@I�Lɢ�!?� ����@�8��Y�ٿY"�T���@nZf�P 4@n^�_ŏ!?�������@0{��!�ٿlc����@tÞ¨4@4ޟ�n�!?G#�m���@0{��!�ٿlc����@tÞ¨4@4ޟ�n�!?G#�m���@0{��!�ٿlc����@tÞ¨4@4ޟ�n�!?G#�m���@0{��!�ٿlc����@tÞ¨4@4ޟ�n�!?G#�m���@0{��!�ٿlc����@tÞ¨4@4ޟ�n�!?G#�m���@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@\D����ٿQ����q�@��¯ 4@�xX�g�!?��8�zy�@x*�ĥٿ�W�z�@mw'� 4@ݸJ�R�!?Ф��;�@x*�ĥٿ�W�z�@mw'� 4@ݸJ�R�!?Ф��;�@x*�ĥٿ�W�z�@mw'� 4@ݸJ�R�!?Ф��;�@x*�ĥٿ�W�z�@mw'� 4@ݸJ�R�!?Ф��;�@w��D�ٿR�ԥT�@�3�D\�3@�rBx�!?���}t�@w��D�ٿR�ԥT�@�3�D\�3@�rBx�!?���}t�@w��D�ٿR�ԥT�@�3�D\�3@�rBx�!?���}t�@w��D�ٿR�ԥT�@�3�D\�3@�rBx�!?���}t�@w��D�ٿR�ԥT�@�3�D\�3@�rBx�!?���}t�@�����ٿ=�i D�@���s* 4@��[��!?��J����@�����ٿ=�i D�@���s* 4@��[��!?��J����@�����ٿ=�i D�@���s* 4@��[��!?��J����@�����ٿ=�i D�@���s* 4@��[��!?��J����@�����ٿ=�i D�@���s* 4@��[��!?��J����@�����ٿ=�i D�@���s* 4@��[��!?��J����@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@;4,�ٿc�{o��@��t���3@�vzt��!?d��l�@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@�����ٿ Ȑ�o��@��e(�3@7sG��!?�%:���@5���ٿ�+�CQ��@��P���3@��U���!?�yC�G�@5���ٿ�+�CQ��@��P���3@��U���!?�yC�G�@5���ٿ�+�CQ��@��P���3@��U���!?�yC�G�@5���ٿ�+�CQ��@��P���3@��U���!?�yC�G�@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@�'�;�ٿ;�=���@��_���3@������!?�̙���@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@���'�ٿf����@��<� 4@^,�A�!?"Hp�?�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@�>��!�ٿ��Hm��@�O�#�4@O%<�y�!?�A��^�@0��,�ٿ=�NP��@;N��� 4@K(��l�!?�Q��r�@���"�ٿuP|t��@����4@���X��!?4(�+;�@���"�ٿuP|t��@����4@���X��!?4(�+;�@���"�ٿuP|t��@����4@���X��!?4(�+;�@���"�ٿuP|t��@����4@���X��!?4(�+;�@�Ш6��ٿ�*R/��@r���4@ۛ�Z��!?R,�<GX�@�Ш6��ٿ�*R/��@r���4@ۛ�Z��!?R,�<GX�@�Ш6��ٿ�*R/��@r���4@ۛ�Z��!?R,�<GX�@�Ш6��ٿ�*R/��@r���4@ۛ�Z��!?R,�<GX�@�Ш6��ٿ�*R/��@r���4@ۛ�Z��!?R,�<GX�@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@Я�!�ٿ�32uS�@F3
�� 4@Y�Nt��!?��j����@�`�ٿ�"��Z��@�p��Q4@ہ�l��!?���@��@�`�ٿ�"��Z��@�p��Q4@ہ�l��!?���@��@��a���ٿ���Z���@w�$$9 4@��d��!?k����@��a���ٿ���Z���@w�$$9 4@��d��!?k����@��a���ٿ���Z���@w�$$9 4@��d��!?k����@�h��ٿ��S����@��=Ƹ4@2�C�Ə!?�~0�@�h��ٿ��S����@��=Ƹ4@2�C�Ə!?�~0�@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@��\n�ٿ������@�K��4@������!?ՠ\n���@e�tm��ٿ�ͷ8���@�!�,44@������!??��l��@e�tm��ٿ�ͷ8���@�!�,44@������!??��l��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@�7�ݟٿ��Iy�@ç��� 4@(bvՏ!?�_�Q��@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@^[��ٿ~���@���0�3@׸���!?�ʝ�Gc�@�� �ٿl�����@ǵd)�3@���Ə!?%V�_�@�� �ٿl�����@ǵd)�3@���Ə!?%V�_�@'+��q�ٿ��:��@�0E�=�3@������!?a�5O��@'+��q�ٿ��:��@�0E�=�3@������!?a�5O��@2�"�C�ٿ�����@�(0���3@�����!? L�	f��@2�"�C�ٿ�����@�(0���3@�����!? L�	f��@hE�c �ٿ�#sP�Y�@�3���3@�A9��!?E���/��@K���c�ٿETJPG%�@.LES� 4@@�ꧏ!?�u�R^"�@K���c�ٿETJPG%�@.LES� 4@@�ꧏ!?�u�R^"�@��`l��ٿ9��9<�@o&\]A4@	���!?.���=�@��`l��ٿ9��9<�@o&\]A4@	���!?.���=�@��`l��ٿ9��9<�@o&\]A4@	���!?.���=�@��`l��ٿ9��9<�@o&\]A4@	���!?.���=�@��`l��ٿ9��9<�@o&\]A4@	���!?.���=�@>iio"�ٿ�G�sz�@]Z���3@�+�_��!?�����@>iio"�ٿ�G�sz�@]Z���3@�+�_��!?�����@>iio"�ٿ�G�sz�@]Z���3@�+�_��!?�����@>iio"�ٿ�G�sz�@]Z���3@�+�_��!?�����@�2߇8�ٿ���-�@�ɀ\��3@*xv���!?��$ɑ�@�2߇8�ٿ���-�@�ɀ\��3@*xv���!?��$ɑ�@�	�z�ٿ��_�@Y��s��3@Z�l�Տ!?������@�	�z�ٿ��_�@Y��s��3@Z�l�Տ!?������@�	�z�ٿ��_�@Y��s��3@Z�l�Տ!?������@�	�z�ٿ��_�@Y��s��3@Z�l�Տ!?������@Hbk���ٿ�j�?3�@��QW�3@I\�~�!?Vl;�"(�@Hbk���ٿ�j�?3�@��QW�3@I\�~�!?Vl;�"(�@Hbk���ٿ�j�?3�@��QW�3@I\�~�!?Vl;�"(�@Hbk���ٿ�j�?3�@��QW�3@I\�~�!?Vl;�"(�@Hbk���ٿ�j�?3�@��QW�3@I\�~�!?Vl;�"(�@R}� ��ٿ�gB��@IU���3@S�Z[��!?ʽ����@���`O�ٿ���V���@�0`��3@C�\Κ�!?�r����@��x<�ٿ&�.=��@�mQ���3@	<���!?�5��|��@��x<�ٿ&�.=��@�mQ���3@	<���!?�5��|��@��x<�ٿ&�.=��@�mQ���3@	<���!?�5��|��@#D���ٿt(�?r�@�/~�Y4@�ɶ��!?�u@P��@#D���ٿt(�?r�@�/~�Y4@�ɶ��!?�u@P��@#D���ٿt(�?r�@�/~�Y4@�ɶ��!?�u@P��@����O�ٿy�-
�h�@D����3@w®A�!?��r���@����O�ٿy�-
�h�@D����3@w®A�!?��r���@� ؘըٿ_���0��@�L[?��3@�2��c�!?�9���@� ؘըٿ_���0��@�L[?��3@�2��c�!?�9���@C,�Z�ٿ���A��@<Q+p��3@3���!?��$o<Q�@C,�Z�ٿ���A��@<Q+p��3@3���!?��$o<Q�@�,�\�ٿ�3�t��@�6��4@b�i6�!?.$^8Q��@�QG�ٿ���q��@���Ά4@�%�:�!?:k��1�@�QG�ٿ���q��@���Ά4@�%�:�!?:k��1�@�QG�ٿ���q��@���Ά4@�%�:�!?:k��1�@���%�ٿ|l�����@X��k4@̏�/s�!? i2��@��'�ٿP}]%U��@��\>4@i��5ُ!?����@��'�ٿP}]%U��@��\>4@i��5ُ!?����@��'�ٿP}]%U��@��\>4@i��5ُ!?����@��'�ٿP}]%U��@��\>4@i��5ُ!?����@��'�ٿP}]%U��@��\>4@i��5ُ!?����@��'�ٿP}]%U��@��\>4@i��5ُ!?����@@x�*~�ٿ��mc[�@��t� 4@�T���!?�&�Ӿ�@@x�*~�ٿ��mc[�@��t� 4@�T���!?�&�Ӿ�@@x�*~�ٿ��mc[�@��t� 4@�T���!?�&�Ӿ�@@x�*~�ٿ��mc[�@��t� 4@�T���!?�&�Ӿ�@u�s��ٿ���J{�@������3@��昏!?$�,��:�@u�s��ٿ���J{�@������3@��昏!?$�,��:�@u�s��ٿ���J{�@������3@��昏!?$�,��:�@u�s��ٿ���J{�@������3@��昏!?$�,��:�@u�s��ٿ���J{�@������3@��昏!?$�,��:�@�o+�ٿ�����A�@#%�4�3@�V��Ï!?��iz���@����_�ٿ�@�U��@�md9�3@����[�!?��,���@����_�ٿ�@�U��@�md9�3@����[�!?��,���@����_�ٿ�@�U��@�md9�3@����[�!?��,���@����ٿ���cF�@1�-� �3@�A�G�!?��"��U�@����ٿ���cF�@1�-� �3@�A�G�!?��"��U�@�
�{�ٿ��7��@����3@
.�~�!?IΗh��@�
�{�ٿ��7��@����3@
.�~�!?IΗh��@�
�{�ٿ��7��@����3@
.�~�!?IΗh��@�
�{�ٿ��7��@����3@
.�~�!?IΗh��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@����ٿU%!�~��@��J�t�3@�ϴB�!?�$�6��@s��z�ٿ����?�@T߇��3@��g�K�!?J h�@dߚV�ٿ��)`��@IP8P4@�[O!?z9 ����@dߚV�ٿ��)`��@IP8P4@�[O!?z9 ����@dߚV�ٿ��)`��@IP8P4@�[O!?z9 ����@dߚV�ٿ��)`��@IP8P4@�[O!?z9 ����@dߚV�ٿ��)`��@IP8P4@�[O!?z9 ����@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@��	�ٿ�Y
��@gv�h�4@]b��b�!?tD��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@O�Ӡٿ=J�\ɧ�@	���� 4@���O�!?����
��@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@1���\�ٿg*{X �@�K�?��3@b�>�`�!?5��E(;�@9qe�o�ٿ�oB���@q  4@��d�؏!?`G���@9qe�o�ٿ�oB���@q  4@��d�؏!?`G���@9qe�o�ٿ�oB���@q  4@��d�؏!?`G���@9qe�o�ٿ�oB���@q  4@��d�؏!?`G���@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@2��ߧٿq#>�1��@��;���3@�}Z��!?�,,��@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@��Q�ٿ�%�g�_�@
*7�	 4@Z���ߏ!?�O�b$J�@�kV̠ٿrT��1�@[DV;� 4@ʕ�`�!?�H燉�@�kV̠ٿrT��1�@[DV;� 4@ʕ�`�!?�H燉�@�kV̠ٿrT��1�@[DV;� 4@ʕ�`�!?�H燉�@+�&��ٿ
e�`C�@�b<�� 4@U�CW�!?��WA���@+�&��ٿ
e�`C�@�b<�� 4@U�CW�!?��WA���@+�&��ٿ
e�`C�@�b<�� 4@U�CW�!?��WA���@+�&��ٿ
e�`C�@�b<�� 4@U�CW�!?��WA���@+�&��ٿ
e�`C�@�b<�� 4@U�CW�!?��WA���@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@�����ٿ��t���@|MJ@7 4@z�ϛ.�!?ۍ��a�@[M����ٿL	���@�@Wr�3@NC^7��!?�-�(��@[M����ٿL	���@�@Wr�3@NC^7��!?�-�(��@?n��ˬٿ=ͺ1��@$�>���3@����!?�&����@?n��ˬٿ=ͺ1��@$�>���3@����!?�&����@�%��ٿ=z����@'�M4@�3^��!?r��Y���@�%��ٿ=z����@'�M4@�3^��!?r��Y���@�%��ٿ=z����@'�M4@�3^��!?r��Y���@�%��ٿ=z����@'�M4@�3^��!?r��Y���@���&��ٿ�6��C�@zA�I�4@7[��!?��¹���@���&��ٿ�6��C�@zA�I�4@7[��!?��¹���@��܍��ٿ��P��z�@�M�- 4@���q�!?Шx���@��܍��ٿ��P��z�@�M�- 4@���q�!?Шx���@��܍��ٿ��P��z�@�M�- 4@���q�!?Шx���@��܍��ٿ��P��z�@�M�- 4@���q�!?Шx���@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@A����ٿT�����@�pē  4@�=0�!?2k3IZ�@�+%���ٿ֚
D�@x��R4@i~�ӏ!?��~t�@�+%���ٿ֚
D�@x��R4@i~�ӏ!?��~t�@'I���ٿ�,����@�a̅4@o=����!?������@�_N��ٿT�,ME3�@� P�4@`���!?؆����@�_N��ٿT�,ME3�@� P�4@`���!?؆����@�_N��ٿT�,ME3�@� P�4@`���!?؆����@�_N��ٿT�,ME3�@� P�4@`���!?؆����@�_N��ٿT�,ME3�@� P�4@`���!?؆����@�_N��ٿT�,ME3�@� P�4@`���!?؆����@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@G��ٿ���Ƅ�@,���4@u+�ŏ!?�z�]���@9�[ʰ�ٿ���~z�@�+Wc4@�ď!?��"y��@9�[ʰ�ٿ���~z�@�+Wc4@�ď!?��"y��@9�[ʰ�ٿ���~z�@�+Wc4@�ď!?��"y��@>�?��ٿ=�I���@�	��4@�;��!?��F��e�@�6P~�ٿ]o���"�@�F�$4@�"��!?���z��@�6P~�ٿ]o���"�@�F�$4@�"��!?���z��@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@q.i,�ٿ�iɋ�	�@{	��4@�k��Z�!?��{�>R�@?U �c�ٿ��� �[�@kZ;ъ�3@� ���!?����@?U �c�ٿ��� �[�@kZ;ъ�3@� ���!?����@p=�R �ٿ��A���@����3@11:��!?��B'�@p=�R �ٿ��A���@����3@11:��!?��B'�@p=�R �ٿ��A���@����3@11:��!?��B'�@p=�R �ٿ��A���@����3@11:��!?��B'�@p=�R �ٿ��A���@����3@11:��!?��B'�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@d_�_�ٿ��U�
�@>Y˛��3@{�h�!?J���׷�@t�ٿ�4��#�@91���3@����!?G?Yƒ��@t�ٿ�4��#�@91���3@����!?G?Yƒ��@t�ٿ�4��#�@91���3@����!?G?Yƒ��@OS3/�ٿٖ�o�C�@ ���4@�M���!?�?!Ӗ�@OS3/�ٿٖ�o�C�@ ���4@�M���!?�?!Ӗ�@OS3/�ٿٖ�o�C�@ ���4@�M���!?�?!Ӗ�@~��y�ٿ؅VדM�@]�� 4@�6�!?q3O���@~��y�ٿ؅VדM�@]�� 4@�6�!?q3O���@~��y�ٿ؅VדM�@]�� 4@�6�!?q3O���@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@�%\�ٿ2&8eM��@�a�{4@`+���!?��?ɪ��@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@I.�ҨٿKC�.��@W!�D 4@2�Az��!?���*�b�@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@>A\�ٿl^�}h��@��%�4@{�f>��!?HK����@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�uުٿ˿�i���@�N:��4@Kw6���!?~FBt)��@�9R��ٿ���!~�@>�L�4@f胏!?Q��	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@�~<̙�ٿh�kg�>�@�N|y�4@�-�9��!?\�	���@,ĵ���ٿ7� �*�@!���U 4@��%:�!?0�-�a�@�ä��ٿ�uG('A�@�Dc�3@��_�!?�ŠY�@�ä��ٿ�uG('A�@�Dc�3@��_�!?�ŠY�@�ä��ٿ�uG('A�@�Dc�3@��_�!?�ŠY�@}�'���ٿ�>� ��@5=|,` 4@8s����!?�?cv`�@}�'���ٿ�>� ��@5=|,` 4@8s����!?�?cv`�@}�'���ٿ�>� ��@5=|,` 4@8s����!?�?cv`�@}�'���ٿ�>� ��@5=|,` 4@8s����!?�?cv`�@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@=D�j��ٿ@�	�:&�@��)���3@]�v��!?9�nO��@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@aVeI~�ٿ�E%��@0Ί� 4@q�1ڞ�!?� ����@�xn��ٿ˧}"��@����4@_?���!?����I��@�xn��ٿ˧}"��@����4@_?���!?����I��@�xn��ٿ˧}"��@����4@_?���!?����I��@�xn��ٿ˧}"��@����4@_?���!?����I��@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@DU��i�ٿ��w͸�@�F��4@�D�[��!?LI:]�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@2�"D�ٿ[ݨ���@������3@��dݏ!?%�t��\�@e�آٿ�+ˮ�1�@�ZT��3@��󡶏!?Y�J�-5�@e�آٿ�+ˮ�1�@�ZT��3@��󡶏!?Y�J�-5�@e�آٿ�+ˮ�1�@�ZT��3@��󡶏!?Y�J�-5�@��S�ٿ�K��4�@�!fɭ 4@����`�!?q�V�@��S�ٿ�K��4�@�!fɭ 4@����`�!?q�V�@��S�ٿ�K��4�@�!fɭ 4@����`�!?q�V�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@�Ͼ��ٿ����f��@T�[�I4@$�B�V�!?2�ڪl�@M9P���ٿ*����@�4�G4@2Ũm-�!?����@M9P���ٿ*����@�4�G4@2Ũm-�!?����@M9P���ٿ*����@�4�G4@2Ũm-�!?����@N�'@�ٿd�=#Ka�@��� 4@���ey�!?o�5��K�@N�'@�ٿd�=#Ka�@��� 4@���ey�!?o�5��K�@N�'@�ٿd�=#Ka�@��� 4@���ey�!?o�5��K�@.���Z�ٿ.#��ե�@�ѕ� 4@@�˷\�!?����@�@.���Z�ٿ.#��ե�@�ѕ� 4@@�˷\�!?����@�@.���Z�ٿ.#��ե�@�ѕ� 4@@�˷\�!?����@�@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��5�A�ٿ�QXP��@�����3@�|�~�!?*�D���@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@��[�L�ٿ�����&�@�#x���3@$z�.��!?��pԹU�@�oS��ٿS~^�x�@ڷ}r��3@��@R�!?:�{�@��l���ٿ-�=�6��@��Ξ� 4@a�;[��!?��"M��@��l���ٿ-�=�6��@��Ξ� 4@a�;[��!?��"M��@aϓ�W�ٿM����@Ng}�Q 4@�8T���!?��YC�@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@̀��.�ٿ�߿@ܥ�@=�04@�Seӽ�!?M��3��@lr�$8�ٿ8����@���S4@������!?gj;#�N�@lr�$8�ٿ8����@���S4@������!?gj;#�N�@lr�$8�ٿ8����@���S4@������!?gj;#�N�@O�f�ëٿevInM�@<c9w�4@Ɏ��!?�¾z���@bQe�ٿ�/ C��@~�4@��G��!?�Q�T�@bQe�ٿ�/ C��@~�4@��G��!?�Q�T�@bQe�ٿ�/ C��@~�4@��G��!?�Q�T�@��gcҧٿG�[H�@�UU� 4@('���!?LKɱpD�@��gcҧٿG�[H�@�UU� 4@('���!?LKɱpD�@��*���ٿx�j����@fi*6�4@�P[�܏!?��]iQ��@f	(B��ٿ�_�I=�@V�nWA4@a�4:��!?���R���@f	(B��ٿ�_�I=�@V�nWA4@a�4:��!?���R���@�fō�ٿ&����@��44@�w$ҏ!?=���}5�@�~���ٿ*�=���@���ɣ4@7fF�!?��~�[�@�~���ٿ*�=���@���ɣ4@7fF�!?��~�[�@X��D�ٿ̡��D�@R?�4@:�󆯏!?<�4�>�@X��D�ٿ̡��D�@R?�4@:�󆯏!?<�4�>�@X��D�ٿ̡��D�@R?�4@:�󆯏!?<�4�>�@X��D�ٿ̡��D�@R?�4@:�󆯏!?<�4�>�@�\���ٿ\o<,���@�1�p�3@#�ɑ�!?Ī:��%�@�\���ٿ\o<,���@�1�p�3@#�ɑ�!?Ī:��%�@�\���ٿ\o<,���@�1�p�3@#�ɑ�!?Ī:��%�@�\���ٿ\o<,���@�1�p�3@#�ɑ�!?Ī:��%�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@�/3�ٿbC�����@��14@n�8�F�!?�S{�@���ٿ`*Č��@n0U�y4@]mn���!?$.��n-�@���ٿ`*Č��@n0U�y4@]mn���!?$.��n-�@���ٿ`*Č��@n0U�y4@]mn���!?$.��n-�@���ٿ`*Č��@n0U�y4@]mn���!?$.��n-�@���ٿ`*Č��@n0U�y4@]mn���!?$.��n-�@\�)I�ٿTMS��@�_�4@�����!?�Z ��@\�)I�ٿTMS��@�_�4@�����!?�Z ��@\�)I�ٿTMS��@�_�4@�����!?�Z ��@\�)I�ٿTMS��@�_�4@�����!?�Z ��@q��)A�ٿX������@eV��� 4@���T��!?����T��@q��)A�ٿX������@eV��� 4@���T��!?����T��@ �s��ٿ��FH���@F<�fX 4@��t�!?�C���@ �s��ٿ��FH���@F<�fX 4@��t�!?�C���@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@.�R�d�ٿ�K�1 ��@�����3@ӛ�!?۴=����@��'��ٿ���!�@x.%t�4@�nis�!?4����@��'��ٿ���!�@x.%t�4@�nis�!?4����@��lϣ�ٿ X�4��@ۊ�
� 4@�m�ӏ!?���i��@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@��V.�ٿ	�*���@���n4@G����!?��>k���@�ӫu�ٿ	��h��@��L�#4@��Q,0�!?��&��@�_v���ٿ�:7�%�@��: - 4@�L)ӏ!?�V69M��@�_v���ٿ�:7�%�@��: - 4@�L)ӏ!?�V69M��@�_v���ٿ�:7�%�@��: - 4@�L)ӏ!?�V69M��@�_v���ٿ�:7�%�@��: - 4@�L)ӏ!?�V69M��@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@{~��[�ٿX�"2��@�����3@G#@
c�!?h<�G[�@��b��ٿ�1�l�t�@��=gq4@���?�!?��:�@��b��ٿ�1�l�t�@��=gq4@���?�!?��:�@vӾ�z�ٿ6�Y?�D�@�N�+�3@�ucn�!?��f2f��@vӾ�z�ٿ6�Y?�D�@�N�+�3@�ucn�!?��f2f��@vӾ�z�ٿ6�Y?�D�@�N�+�3@�ucn�!?��f2f��@vӾ�z�ٿ6�Y?�D�@�N�+�3@�ucn�!?��f2f��@P��ٿGC1�2�@a���� 4@���O��!?&t|���@P��ٿGC1�2�@a���� 4@���O��!?&t|���@P��ٿGC1�2�@a���� 4@���O��!?&t|���@P��ٿGC1�2�@a���� 4@���O��!?&t|���@P��ٿGC1�2�@a���� 4@���O��!?&t|���@P��ٿGC1�2�@a���� 4@���O��!?&t|���@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@�t8�*�ٿ��V��@��D| 4@�T3eR�!?*������@��O��ٿ�=q����@J �4b 4@P���F�!?�71?�6�@��O��ٿ�=q����@J �4b 4@P���F�!?�71?�6�@��O��ٿ�=q����@J �4b 4@P���F�!?�71?�6�@��O��ٿ�=q����@J �4b 4@P���F�!?�71?�6�@�n9k�ٿ���I�@I�h4@�lZ��!?���j�@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@��xՄ�ٿ�k�^<��@���\'4@S�����!?�
߭t��@�4�ٿ�����@Y�~m 4@&��~Џ!?����^E�@�4�ٿ�����@Y�~m 4@&��~Џ!?����^E�@�4�ٿ�����@Y�~m 4@&��~Џ!?����^E�@�4�ٿ�����@Y�~m 4@&��~Џ!?����^E�@�4�ٿ�����@Y�~m 4@&��~Џ!?����^E�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@p��洙ٿQ�Z����@͕�*��3@9|����!?�`R��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@O�yיٿ������@�S���3@0���!?Z��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@$ {ۙٿP:� ��@
c� 4@z ��!?�}��o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@�itgݙٿ |�: ��@���� 4@�SĂ�!?����o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@h�N�ٿ�y�N ��@��B 4@zߴ�!?�2��o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@�����ٿ�ک8 ��@�Q�1 4@t D���!?��"�o�@m�q�ٿ]�g* ��@2Y�� 4@����-�!?��6�o�@m�q�ٿ]�g* ��@2Y�� 4@����-�!?��6�o�@m�q�ٿ]�g* ��@2Y�� 4@����-�!?��6�o�@�����ٿ�ߴ= ��@�d1- 4@��R�j�!?+�]�o�@�����ٿ�ߴ= ��@�d1- 4@��R�j�!?+�]�o�@�����ٿ�ߴ= ��@�d1- 4@��R�j�!?+�]�o�@�����ٿ�ߴ= ��@�d1- 4@��R�j�!?+�]�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�+�}�ٿ��D ��@�Wz> 4@k�V8��!?e�$�o�@�]�Sޙٿ/��7 ��@�z� 4@��k�M�!?<<E!�o�@�]�Sޙٿ/��7 ��@�z� 4@��k�M�!?<<E!�o�@�]�Sޙٿ/��7 ��@�z� 4@��k�M�!?<<E!�o�@�]�Sޙٿ/��7 ��@�z� 4@��k�M�!?<<E!�o�@�]�Sޙٿ/��7 ��@�z� 4@��k�M�!?<<E!�o�@�e��ԙٿ��P1 ��@"I3� 4@�A�!?e�� �o�@�e��ԙٿ��P1 ��@"I3� 4@�A�!?e�� �o�@�e��ԙٿ��P1 ��@"I3� 4@�A�!?e�� �o�@�e��ԙٿ��P1 ��@"I3� 4@�A�!?e�� �o�@�e��ԙٿ��P1 ��@"I3� 4@�A�!?e�� �o�@��ԙٿ��* ��@r{Z� 4@$L\2��!?u�L!�o�@��znיٿ��|$ ��@3��� 4@�ا|=�!?k�o�@��znיٿ��|$ ��@3��� 4@�ا|=�!?k�o�@��ڙٿ�9�  ��@t�X� 4@i`]m�!?�C(�o�@�ٷaٙٿ"�k ��@��, 4@�Wd܏!?&��&�o�@�ٷaٙٿ"�k ��@��, 4@�Wd܏!?&��&�o�@�ٷaٙٿ"�k ��@��, 4@�Wd܏!?&��&�o�@�ÜЙٿ]l ��@^��@ 4@��I��!?W�$�o�@ӳh%͙ٿu�����@��
1 4@��L��!?|��#�o�@kQ�љٿ�vr����@56�  4@�����!?�ߡ �o�@kQ�љٿ�vr����@56�  4@�����!?�ߡ �o�@`l#ʙٿ��1 ��@�mmi  4@K��4��!?[ۖ�o�@�Im̙ٿe ��@9�Cp  4@3uڏ!?3|q!�o�@g��Йٿ]۔ ��@�@�  4@y�~�%�!?�>m"�o�@�L�P֙ٿ�5 ��@�
  4@7���E�!?��8 �o�@!�֙ٿØ[ ��@�m{���3@|e�S�!?N��o�@�hW�әٿ�= ��@��  4@_`
d�!?��^�o�@I���Ιٿ��� ��@;��  4@�S@f�!?�|H�o�@)��ƙٿ�^ ��@d�f��3@���y��!?j`,�o�@��R��ٿ.������@�����3@�Xh)��!?�ש�o�@*����ٿAbM����@��b���3@��w���!?y���o�@Olz�ٿ�Z�����@	�����3@?�)�Ï!?V>��o�@Olz�ٿ�Z�����@	�����3@?�)�Ï!?V>��o�@Olz�ٿ�Z�����@	�����3@?�)�Ï!?V>��o�@N=��ٿȴ�����@�:&���3@�����!?B)��o�@N=��ٿȴ�����@�:&���3@�����!?B)��o�@�Ր��ٿ�NA����@:(�d��3@�C�!?��o�o�@�ʙٿ�C����@j�����3@1G6 <�!?�g~�o�@�ʙٿ�C����@j�����3@1G6 <�!?�g~�o�@�ʙٿ�C����@j�����3@1G6 <�!?�g~�o�@\�ȥΙٿH�s����@��(���3@��vI��!?����o�@\�ȥΙٿH�s����@��(���3@��vI��!?����o�@\�ȥΙٿH�s����@��(���3@��vI��!?����o�@�D�֙ٿ/z�  ��@���- 4@��a"ۏ!?Q���o�@e%1�֙ٿvC� ��@vw.L 4@�-�/͏!?���o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@�יٿ Q ��@q'�B 4@;�]�T�!?��o�o�@Ȕ|�ۙٿ��
 ��@�s�2 4@`���!?*g��o�@H�(ؙٿT�� ��@WK� 4@��6�!?�p��o�@�Ff�ٙٿɋ� ��@��S� 4@��[�!?�l��o�@Ъ&�֙ٿdOx ��@^W�T 4@E�z�Z�!?���o�@Zi_ۙٿ@�7& ��@( 4@�@A�!?�� �o�@sZ)�ٿO�3 ��@��r� 4@���@�!?�a%�o�@sZ)�ٿO�3 ��@��r� 4@���@�!?�a%�o�@sZ)�ٿO�3 ��@��r� 4@���@�!?�a%�o�@sZ)�ٿO�3 ��@��r� 4@���@�!?�a%�o�@-5�ޙٿ��) ��@���� 4@d�_^ �!?FP&�o�@-5�ޙٿ��) ��@���� 4@d�_^ �!?FP&�o�@-5�ޙٿ��) ��@���� 4@d�_^ �!?FP&�o�@�h�ۙٿm��% ��@[�b# 4@k9���!?& �%�o�@��Ǐڙٿ�2 ��@�im` 4@�l�s��!?�PY%�o�@��Ǐڙٿ�2 ��@�im` 4@�l�s��!?�PY%�o�@�O�ٙٿ�dI ��@��� 4@��p��!?8�!�o�@}y
oܙٿr ��@�vɤ 4@s�'��!?�M�!�o�@}y
oܙٿr ��@�vɤ 4@s�'��!?�M�!�o�@}y
oܙٿr ��@�vɤ 4@s�'��!?�M�!�o�@}y
oܙٿr ��@�vɤ 4@s�'��!?�M�!�o�@��59ޙٿ��5 ��@L�^[ 4@������!?�'�o�@�o����ٿ9�� ��@9�+ 4@�Ϲ}��!?S���o�@�o����ٿ9�� ��@9�+ 4@�Ϲ}��!?S���o�@�o����ٿ9�� ��@9�+ 4@�Ϲ}��!?S���o�@��}��ٿ�A ��@�=�� 4@\v�!?���o�@��J�ߙٿ��� ��@�O�� 4@�@�!?����o�@?/�ߙٿ�ֿ
 ��@6O* 4@���f[�!?��o�@�V���ٿ"&� ��@|4I 4@�"�Xm�!?����o�@�pT��ٿ�EF ��@7�j� 4@�uK�!?�Ѐ�o�@�pT��ٿ�EF ��@7�j� 4@�uK�!?�Ѐ�o�@�pT��ٿ�EF ��@7�j� 4@�uK�!?�Ѐ�o�@g]%��ٿ�-% ��@` 4@����!?��1�o�@��<��ٿ��$ ��@9�'p 4@�j�	+�!?.)�o�@��<��ٿ��$ ��@9�'p 4@�j�	+�!?.)�o�@���)�ٿ>pX$ ��@�:�h 4@����!?*��o�@z9�ܙٿ��. ��@�Xc 4@\ȓ���!?.12�o�@z9�ܙٿ��. ��@�Xc 4@\ȓ���!?.12�o�@l�(ޙٿ|�2 ��@�Չ� 4@���Nm�!?d� �o�@B���ݙٿ-�6> ��@�7? 4@�C���!?5?*#�o�@����ޙٿ@��9 ��@�/`- 4@U��^!?�!!�o�@Gӡ��ٿ
��< ��@i��o 4@y��6��!?R�)!�o�@Gӡ��ٿ
��< ��@i��o 4@y��6��!?R�)!�o�@Gӡ��ٿ
��< ��@i��o 4@y��6��!?R�)!�o�@Gӡ��ٿ
��< ��@i��o 4@y��6��!?R�)!�o�@'�Qݙٿ/v"D ��@�� 4@|&
V��!?Mrx#�o�@���Gיٿ��> ��@m�� 4@ߐI��!?X'�#�o�@JBIoԙٿ�y�@ ��@�* 4@&m</j�!?1l�!�o�@�r[�әٿE'0B ��@�ZW 4@�*ӏH�!?�@�!�o�@��]gΙٿn�A ��@��ƻ 4@�����!?<7�!�o�@��̪Йٿ�B ��@Oyr 4@a�����!?l.�!�o�@|�c�әٿM��P ��@�� 4@?�<���!?N|,&�o�@�_�sԙٿR�tO ��@�� 4@����!?d.�%�o�@d#�љٿ��
Z ��@�W� 4@��MZ�!?��J'�o�@d#�љٿ��
Z ��@�W� 4@��MZ�!?��J'�o�@�F;ҙٿ��\ ��@�� 4@�ͬ Z�!?y��)�o�@�I:;ԙٿQ��Z ��@I:�� 4@��\]�!?�@�)�o�@��&Ιٿy�sX ��@�T� 4@/L��c�!?�v(�o�@�BGԙٿA
b ��@��	 4@�A�P��!?sa�(�o�@�BGԙٿA
b ��@��	 4@�A�P��!?sa�(�o�@��2}ԙٿɎT[ ��@�~�� 4@9�ق��!?��'�o�@��2}ԙٿɎT[ ��@�~�� 4@9�ق��!?��'�o�@��2}ԙٿɎT[ ��@�~�� 4@9�ق��!?��'�o�@��2}ԙٿɎT[ ��@�~�� 4@9�ق��!?��'�o�@�Q�Йٿ<��k ��@t�>�
 4@�m���!?��Q*�o�@�<ՙٿ�qe ��@%E��
 4@gd[���!?�(+�o�@�<ՙٿ�qe ��@%E��
 4@gd[���!?�(+�o�@�<ՙٿ�qe ��@%E��
 4@gd[���!?�(+�o�@�<ՙٿ�qe ��@%E��
 4@gd[���!?�(+�o�@�<ՙٿ�qe ��@%E��
 4@gd[���!?�(+�o�@wb0vҙٿ��e ��@��A;
 4@���(�!?0,�o�@���әٿ� �_ ��@��q:	 4@v���!?�!-�o�@$�ԙٿGM&T ��@�].� 4@����!?�B�,�o�@벶Tϙٿ��\c ��@1�	 4@
ӵ�
�!?� p/�o�@��t�ϙٿ��lP ��@�%] 4@a�Dя!?Z��(�o�@��t�ϙٿ��lP ��@�%] 4@a�Dя!?Z��(�o�@�F\Xʙٿj�ko ��@��=�	 4@$�l��!?�~7/�o�@�F\Xʙٿj�ko ��@��=�	 4@$�l��!?�~7/�o�@�F\Xʙٿj�ko ��@��=�	 4@$�l��!?�~7/�o�@���ęٿ�f� ��@�{� 4@`�F��!?.��5�o�@���ęٿ�f� ��@�{� 4@`�F��!?.��5�o�@�b�Ùٿ,��� ��@�F�	 4@�Y&e��!?�}5�o�@.[�ٿ�Ӏ� ��@���< 4@��#��!?'�,;�o�@	*��ٿ	n&� ��@�H� 4@�}j��!?���:�o�@��<rșٿ��\� ��@C�Pl 4@%����!?��T7�o�@�~iǙٿ�Fe� ��@жl� 4@2�(/��!?\��;�o�@�7^Tϙٿe(�� ��@�G�� 4@ӵM;��!?$g�3�o�@Gْ�͙ٿ'�� ��@���� 4@���Ę�!?tYZ<�o�@:M��șٿ��&� ��@��� 4@��͏!?�aB@�o�@U��fřٿT��� ��@�݈� 4@�w���!?�}=�o�@5q<�ęٿH�Z� ��@�v�� 4@�4�*��!?�RP?�o�@5q<�ęٿH�Z� ��@�v�� 4@�4�*��!?�RP?�o�@�&��ٿD'�� ��@i+D 4@Q�
�!?� A�o�@Y���ٿ�KA� ��@"�$K 4@��\�!?I~Y<�o�@�@|�ƙٿ�7�� ��@�ľP 4@���&��!?���4�o�@��U���ٿ0X�� ��@��^C 4@٤2�*�!?�$�?�o�@[��řٿ"}�� ��@�LR 4@��B3�!?�m=�o�@��ęٿ�:3� ��@b�� 4@K~��	�!?��v<�o�@��ęٿ�:3� ��@b�� 4@K~��	�!?��v<�o�@�/-շ�ٿFu�� ��@^�f� 4@U+*��!?]B�H�o�@w�v��ٿ�]N��@���� 4@���*�!?Q��P�o�@w�v��ٿ�]N��@���� 4@���*�!?Q��P�o�@w�v��ٿ�]N��@���� 4@���*�!?Q��P�o�@ҕ訙ٿn��%��@_��J 4@|c�<�!?�|�W�o�@ҕ訙ٿn��%��@_��J 4@|c�<�!?�|�W�o�@:m+���ٿ����@�+�� 4@F�@-�!?N<$T�o�@:m+���ٿ����@�+�� 4@F�@-�!?N<$T�o�@n�D��ٿ:E+��@̱Y! 4@���K)�!?c6�Y�o�@��k��ٿinc��@CyK� 4@��c��!?L�e�o�@��k��ٿinc��@CyK� 4@��c��!?L�e�o�@x�����ٿ��i���@ ST# 4@�R��D�!?,��x�o�@��=��ٿ����@#u��" 4@=�`��!?5XYw�o�@��=��ٿ����@#u��" 4@=�`��!?5XYw�o�@GSy��ٿ�c�� ��@��V� 4@W�m�ۏ!?a�K�o�@��'��ٿ��� ��@�+ 4@>G��Џ!?d�DH�o�@�N�Ҫ�ٿ=�� ��@5��+ 4@_�9倏!?�/I�o�@���ٿ�i1 ��@�-z� 4@b*���!?�6�I�o�@-��i��ٿQ��� ��@X�� 4@��#}�!?>�AH�o�@��d��ٿ��}� ��@�� 4@��A�!?�]�A�o�@&�|��ٿEm�c��@��� 4@���ܛ�!?QI[�o�@- ����ٿ���T��@��F� 4@�<%���!?��Z�o�@G�i��ٿ�;�k��@p�� 4@�g����!?r\�[�o�@D̙�ٿ2�4u��@�:�N  4@���ԛ�!?s_�]�o�@D̙�ٿ2�4u��@�:�N  4@���ԛ�!?s_�]�o�@D̙�ٿ2�4u��@�:�N  4@���ԛ�!?s_�]�o�@:�K4��ٿ�Ax��@$'S� 4@d��V�!?��8d�o�@:�K4��ٿ�Ax��@$'S� 4@d��V�!?��8d�o�@��Ր�ٿ"�ɰ��@,3��# 4@jap���!?��p�o�@:M=��ٿ/���@*��~# 4@|�X�!?^�uu�o�@�BC�w�ٿf_���@��B, 4@���׏!?D{H��o�@�ֳ�{�ٿ{���@�H�* 4@Lda[ �!?���o�@6� ��ٿ��8���@�5P% 4@��Z^�!?�>p�o�@��Los�ٿ��E��@;}�/ 4@O����!?�߈�o�@�e��f�ٿ�+'���@CFk�6 4@>u���!?�+۞�o�@��of�ٿrO���@�}77 4@۟L��!?E���o�@���%��ٿ����@�40�* 4@�6~��!?�3�{�o�@���%��ٿ����@�40�* 4@�6~��!?�3�{�o�@	�rE��ٿ�L)���@� `! 4@�w���!?�
�e�o�@�u����ٿ%Ww��@�� 4@5�_ɏ!?O+]�o�@�u����ٿ%Ww��@�� 4@5�_ɏ!?O+]�o�@�u����ٿ%Ww��@�� 4@5�_ɏ!?O+]�o�@�u����ٿ%Ww��@�� 4@5�_ɏ!?O+]�o�@��T��ٿ]�Pr��@P�y�  4@;�,���!?Nf9U�o�@�gF���ٿ[%1Q��@�� 4@GN�܏!?��S�o�@#%k��ٿ2�1��@||LR 4@W�:ȏ!?/�=J�o�@�{䥙ٿ�׺C��@E�#� 4@{�{	��!?�A�S�o�@Bm���ٿ�ɶ��@m�� 4@BC����!?[Z�I�o�@;C�ՙٿ�=�> ��@ʍj� 4@�>����!?P��'�o�@�U���ٿ�X>v ��@3�S�	 4@u��0�!?��1�o�@� ���ٿj�e� ��@���" 4@):X0�!?��P<�o�@qL��̙ٿ�~�S ��@��S 4@ʭ�GB�!?�;.�o�@����ęٿ.�	� ��@�g� 4@�S��f�!?���;�o�@Q��ƙٿ�  ��@Y*Q� 4@�0ڏ!?��@�o�@. �7��ٿ��5���@�ٷ�  4@��s��!?w�l�o�@. �7��ٿ��5���@�ٷ�  4@��s��!?w�l�o�@�μ���ٿ��\� ��@�,� 4@�q��y�!?�c,C�o�@:�gv��ٿ�-�� ��@�* 4@��Q��!?��@�o�@�O�M��ٿ���� ��@u�� 4@��U{��!?��[=�o�@�<��ٿ�Ū���@����3@]�]w�!?�d��o�@�����ٿ��$����@�b�^ 4@g�Tz�!?7-�o�@��{ϙٿ5~W ��@`�X	 4@:�Ox�!?ف�&�o�@��{ϙٿ5~W ��@`�X	 4@:�Ox�!?ف�&�o�@�P���ٿ8N�����@�:O��3@l�s�:�!?��o�@�P���ٿ8N�����@�:O��3@l�s�:�!?��o�@���#�ٿ��h����@�Q����3@a��@�!?&��o�@���#�ٿ��h����@�Q����3@a��@�!?&��o�@���#�ٿ��h����@�Q����3@a��@�!?&��o�@���#�ٿ��h����@�Q����3@a��@�!?&��o�@����ęٿ%ę� ��@�e 4@���|�!?��4>�o�@^����ٿd�&��@^gg� 4@��F��!?KK�H�o�@�.l��ٿͼp��@��/ 4@N �]�!?�T_�o�@F�J�j�ٿ>�Q���@�\��; 4@F,͢X�!?j��o�@F�J�j�ٿ>�Q���@�\��; 4@F,͢X�!?j��o�@F�G�ٿ6�ӝ��@��O 4@��9��!?XJ��o�@ve���ٿx9!���@G��!- 4@�!ߨ��!?]kd�o�@ve���ٿx9!���@G��!- 4@�!ߨ��!?]kd�o�@ve���ٿx9!���@G��!- 4@�!ߨ��!?]kd�o�@5�V��ٿY����@	z�=* 4@U��z�!?m�`Y�o�@��ݿ�ٿ�(a� ��@�m- 4@V♺�!?q�8:�o�@�#�ڙٿ5P] ��@ԕ7 4@,��)|�!?�M�o�@�>��Йٿ��� ��@^��G 4@�PF�!?6��%�o�@�>��Йٿ��� ��@^��G 4@�PF�!?6��%�o�@�>��Йٿ��� ��@^��G 4@�PF�!?6��%�o�@M�l>��ٿ�4� ��@�{� 4@�8��!?��3�o�@ڈ*n��ٿ��#��@�� 4@OW>�i�!?;p?3�o�@�w;!��ٿ�iS4��@�<g� 4@3zo'(�!?dA6�o�@�w;!��ٿ�iS4��@�<g� 4@3zo'(�!?dA6�o�@�w;!��ٿ�iS4��@�<g� 4@3zo'(�!?dA6�o�@�w;!��ٿ�iS4��@�<g� 4@3zo'(�!?dA6�o�@�y�}��ٿ}�]��@�Y�7 4@?ާ܋�!?�Q�j�o�@o�/�w�ٿ��c���@��#? 4@�	��n�!?�6���o�@H9���ٿ�����@s��Uh 4@+�T��!?�s@��o�@H9���ٿ�����@s��Uh 4@+�T��!?�s@��o�@H9���ٿ�����@s��Uh 4@+�T��!?�s@��o�@H9���ٿ�����@s��Uh 4@+�T��!?�s@��o�@H9���ٿ�����@s��Uh 4@+�T��!?�s@��o�@F��>�ٿ`b��	��@��*�� 4@_7S��!?=���o�@��O�ٿ�y���@�Ӫ`� 4@�lu���!?�f�o�@��O�ٿ�y���@�Ӫ`� 4@�lu���!?�f�o�@F�|��ٿ$���@�Sk�� 4@�D�w��!?LEx��o�@�b#�w�ٿ<���@�,�%� 4@h{��x�!?���o�@�b#�w�ٿ<���@�,�%� 4@h{��x�!?���o�@\6-��ٿ��^�
��@U��� 4@�3'�ҏ!?�����o�@\6-��ٿ��^�
��@U��� 4@�3'�ҏ!?�����o�@,U6�ژٿ� x.��@���� 4@+�#v̏!?ycg4�o�@,U6�ژٿ� x.��@���� 4@+�#v̏!?ycg4�o�@qJ�>��ٿ��i��@�)� 4@ ��|��!?��k�o�@qJ�>��ٿ��i��@�)� 4@ ��|��!?��k�o�@�@G:�ٿz�[��@�nx\ 4@F*O�!?��w��o�@MڅU�ٿ�")���@�EI���3@K�u���!?H\��o�@�7�-�ٿ�Y�[���@�6Ha�3@ �YBZ�!?�*ë�o�@�7�-�ٿ�Y�[���@�6Ha�3@ �YBZ�!?�*ë�o�@�J��ܚٿ|"JF���@��Ŋ�3@�O?�g�!?&��o�@�� �ٿ���9���@�Y���3@P����!?�����o�@�� �ٿ���9���@�Y���3@P����!?�����o�@ϾU0d�ٿ�0^����@�����3@�k���!?F��u�o�@9�-���ٿ.r���@�d�m>�3@&3ŏ!?��6�o�@9�-���ٿ.r���@�d�m>�3@&3ŏ!?��6�o�@l�w��ٿMxR���@$�9&�3@V��k�!?O� �o�@l�w��ٿMxR���@$�9&�3@V��k�!?O� �o�@l�w��ٿMxR���@$�9&�3@V��k�!?O� �o�@�K�@�ٿ�1M����@�%��_�3@�Zp �!?��n�o�@�%J��ٿ[�����@��S��3@s�A��!?�2�o�@�zmՆ�ٿ
�Z���@�T�ż�3@&�q�!?B�Q�o�@�zmՆ�ٿ
�Z���@�T�ż�3@&�q�!?B�Q�o�@L�D88�ٿ]�����@*��w�3@+��4��!?�E�k�o�@L�D88�ٿ]�����@*��w�3@+��4��!?�E�k�o�@L�D88�ٿ]�����@*��w�3@+��4��!?�E�k�o�@L�D88�ٿ]�����@*��w�3@+��4��!?�E�k�o�@���/�ٿ�e9���@}�n8��3@�dt{w�!?A2���o�@���/�ٿ�e9���@}�n8��3@�dt{w�!?A2���o�@ qk$��ٿwE�t��@̓m5H 4@�>"uŏ!?Z&�o�@��a���ٿ���{��@�2!2 4@�,�5��!?���o�@�:��ٿ�jJ���@�٢ˊ 4@$��wl�!?z����o�@q�ĸf�ٿ�;�=��@�hq}T 4@E#|��!?��8e�o�@а��u�ٿ9s����@��A�M 4@� y|�!?~2�L�o�@� ���ٿ֓?���@�e��4@�622��!?�	���o�@��\�ٿvq����@��5�o 4@�v����!?�u�$�o�@6����ٿ�X����@��pp 4@���}ȏ!?"�Pd�o�@��.P�ٿ�&%>���@}��7��3@m�17��!?�^1�o�@��a�ٿJ������@ѵ̥O�3@.���k�!?�%
�o�@q�x���ٿ�5����@�6����3@ˏv��!?/���o�@q�x���ٿ�5����@�6����3@ˏv��!?/���o�@q�x���ٿ�5����@�6����3@ˏv��!?/���o�@�����ٿ`�d���@��٤�3@i:�Z��!?�=��o�@u�0�ٿ>I�����@�@
��3@[-�;��!?��E�o�@yN���ٿEk����@��>��3@k~��Ǐ!?P�.��o�@1"�]�ٿ^�f���@� ���3@���r��!?3+���o�@:�5��ٿ�D����@hod� 4@%v���!?�AΑ�o�@2��ٿ}���@Qv��M 4@:��!?1��6�o�@#�q�m�ٿt��R��@�(�3X 4@8u ��!?���^�o�@��v$יٿ��na��@�,�0 4@�`�F��!?�PK��o�@��v$יٿ��na��@�,�0 4@�`�F��!?�PK��o�@KW7�a�ٿ�F���@u��Q 4@|}�v~�!?����o�@�L��Ǘٿc	���@Hi�� 4@��ϵQ�!?i����o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@-tp6�ٿ'� ��@���� 4@�_,�!?�Ÿ�o�@^l(��ٿ�5΅ ��@��j 4@��[]��!?�Xx��o�@^l(��ٿ�5΅ ��@��j 4@��[]��!?�Xx��o�@m�����ٿh�ڌ���@?,��3@��ď!?ۢ���o�@m�����ٿh�ڌ���@?,��3@��ď!?ۢ���o�@m�����ٿh�ڌ���@?,��3@��ď!?ۢ���o�@m�����ٿh�ڌ���@?,��3@��ď!?ۢ���o�@f�rϛٿ��_Z���@�qf26�3@��
r�!?1S���o�@q��~g�ٿf������@,
X���3@�i�G��!?'����o�@q��~g�ٿf������@,
X���3@�i�G��!?'����o�@q��~g�ٿf������@,
X���3@�i�G��!?'����o�@Q۪v��ٿ�����@�^���3@<�!?=	?��o�@>4��~�ٿh�?<���@Ѓ "q�3@m��_��!?)]�>�o�@>4��~�ٿh�?<���@Ѓ "q�3@m��_��!?)]�>�o�@�EQ���ٿE�.����@�p�H�3@{벏!?V,
�o�@���ӛٿ�N����@1�����3@�L�!?V%�%�o�@�/B��ٿ3û���@T�0�3@��6ޙ�!?SMD�o�@�/B��ٿ3û���@T�0�3@��6ޙ�!?SMD�o�@�-sJ2�ٿɼ!��@g�z� 4@�`�׉�!?8R���o�@�-sJ2�ٿɼ!��@g�z� 4@�`�׉�!?8R���o�@�7˖��ٿnG�	��@"��R 4@�\�N͏!?�V�1�o�@$�e��ٿRTt
��@�y��� 4@�{A��!?�)uu�o�@،si}�ٿ�Ip���@�
�e�4@�$���!?`6���o�@��`5�ٿ�g,V%��@_�+��4@�O~�i�!?@���o�@�{���ٿR���@)��{4@$M���!?)w�o�@�{���ٿR���@)��{4@$M���!?)w�o�@�=`��ٿ��.N��@�D<1� 4@{����!? *x��o�@�=`��ٿ��.N��@�D<1� 4@{����!? *x��o�@mi�S��ٿz����@���v�3@��44��!?D��n�o�@mi�S��ٿz����@���v�3@��44��!?D��n�o�@��U��ٿ������@�����3@�M
�!?A���o�@��U��ٿ������@�����3@�M
�!?A���o�@��U��ٿ������@�����3@�M
�!?A���o�@��U��ٿ������@�����3@�M
�!?A���o�@��U��ٿ������@�����3@�M
�!?A���o�@��U��ٿ������@�����3@�M
�!?A���o�@��"v��ٿw�����@������3@������!?���o�@��"v��ٿw�����@������3@������!?���o�@��"v��ٿw�����@������3@������!?���o�@w�:|�ٿn#�����@z|D�3@ <����!?�{<��o�@w�:|�ٿn#�����@z|D�3@ <����!?�{<��o�@^Y�nS�ٿHO����@�a� ��3@}��0��!?�� �o�@c8Ve%�ٿ�z����@sX���3@��+�!?v&�o�@c8Ve%�ٿ�z����@sX���3@��+�!?v&�o�@�Isp�ٿ��}��@F�I�4@�-틏!?ٿ��o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@��L�ߜٿ�i����@I`���3@r��Ԏ�!?ώ�}�o�@	��ٿH�(���@�tXI� 4@��ӟݏ!?���o�@	��ٿH�(���@�tXI� 4@��ӟݏ!?���o�@��`���ٿ��+���@��5�N4@�~�w��!?�����o�@�z��ٿRm�\��@�y\� 4@d� G��!?�bt��o�@�z��ٿRm�\��@�y\� 4@d� G��!?�bt��o�@۫���ٿ����@�7�I��3@SX���!?a=��o�@[@�o�ٿ������@,��� 4@2>��Ǐ!?r����o�@[@�o�ٿ������@,��� 4@2>��Ǐ!?r����o�@[@�o�ٿ������@,��� 4@2>��Ǐ!?r����o�@[@�o�ٿ������@,��� 4@2>��Ǐ!?r����o�@[@�o�ٿ������@,��� 4@2>��Ǐ!?r����o�@��{͜ٿ�n)����@C�� 4@�196��!?��H�o�@j=K�Сٿr���܇�@��	&��3@<�[Ϗ!?_�S�o�@j=K�Сٿr���܇�@��	&��3@<�[Ϗ!?_�S�o�@ ��y��ٿD!Kf��@K?�$� 4@��5�Ï!?1�o�@ ��y��ٿD!Kf��@K?�$� 4@��5�Ï!?1�o�@1~��!�ٿˮUw��@��.��4@��X�P�!?n�צ�o�@1~��!�ٿˮUw��@��.��4@��X�P�!?n�צ�o�@�J~�T�ٿ�!1_��@�$��4@����!?�?QD�o�@�J~�T�ٿ�!1_��@�$��4@����!?�?QD�o�@1��V��ٿ�<����@�nt4@�,M�f�!?k��c�o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@���9�ٿ�˃��@@�d���3@��[��!?�d���o�@�A��g�ٿ���:��@-��x�3@{�i�!?n/?��o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@ol�h`�ٿ�������@� 4@!mg�n�!?y��v�o�@��赡ٿڮ����@fz:� 4@���X�!?�pV�o�@��赡ٿڮ����@fz:� 4@���X�!?�pV�o�@��赡ٿڮ����@fz:� 4@���X�!?�pV�o�@��赡ٿڮ����@fz:� 4@���X�!?�pV�o�@``����ٿcqY�ه�@�e�Z� 4@����֏!?�%�o�@``����ٿcqY�ه�@�e�Z� 4@����֏!?�%�o�@%�[�q�ٿ��b܇�@7����4@�|{Y��!?F���o�@%�[�q�ٿ��b܇�@7����4@�|{Y��!?F���o�@%�[�q�ٿ��b܇�@7����4@�|{Y��!?F���o�@�P2ip�ٿ{\���@���~4@:���!?�Gf�o�@�P2ip�ٿ{\���@���~4@:���!?�Gf�o�@�P2ip�ٿ{\���@���~4@:���!?�Gf�o�@]'�꘠ٿo!�a��@o׾=t 4@Ǟ}�!?ـɦ�o�@]'�꘠ٿo!�a��@o׾=t 4@Ǟ}�!?ـɦ�o�@�
&B��ٿF�*�܇�@nq���3@0�¾ȏ!?#eX��o�@2,���ٿ��}���@s9�g��3@���MЏ!?�����o�@2,���ٿ��}���@s9�g��3@���MЏ!?�����o�@2,���ٿ��}���@s9�g��3@���MЏ!?�����o�@2,���ٿ��}���@s9�g��3@���MЏ!?�����o�@2,���ٿ��}���@s9�g��3@���MЏ!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@z��s�ٿ7N�e��@VRh	�3@y矏͏!?�����o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@�P�a��ٿq�����@��x 4@�x��Ǐ!?��q�o�@m�@Vb�ٿn��e��@� ��4@�z�Y{�!?kL�o�@�$qݶ�ٿ������@�ps�4@s�K�X�!?���:�o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@@5ne�ٿ��Pڇ�@�,qu4@|_�U�!?9�`��o�@8��ޥٿ2�vUч�@R���{�3@% (?U�!?o�uB�o�@]Mh\��ٿ� ���@=~M=��3@?~ES�!?� �q�o�@c� Ŷ�ٿ��l���@�l����3@ّ�f�!?���;�o�@k�� <�ٿ�����@�@��" 4@�&Uʏ!?k�2�o�@k�� <�ٿ�����@�@��" 4@�&Uʏ!?k�2�o�@k�� <�ٿ�����@�@��" 4@�&Uʏ!?k�2�o�@k�� <�ٿ�����@�@��" 4@�&Uʏ!?k�2�o�@k�� <�ٿ�����@�@��" 4@�&Uʏ!?k�2�o�@'�fH'�ٿ'֞2��@�q��i 4@˵��я!?9㧐�o�@'�fH'�ٿ'֞2��@�q��i 4@˵��я!?9㧐�o�@'�fH'�ٿ'֞2��@�q��i 4@˵��я!?9㧐�o�@'�fH'�ٿ'֞2��@�q��i 4@˵��я!?9㧐�o�@>>k{Ԧٿ��f�܇�@��Ŀ�4@�^�YG�!?�N��o�@>>k{Ԧٿ��f�܇�@��Ŀ�4@�^�YG�!?�N��o�@:��y1�ٿ��4��@P	SH+ 4@�ӲL�!?��M�o�@:��y1�ٿ��4��@P	SH+ 4@�ӲL�!?��M�o�@:��y1�ٿ��4��@P	SH+ 4@�ӲL�!?��M�o�@:��y1�ٿ��4��@P	SH+ 4@�ӲL�!?��M�o�@:��y1�ٿ��4��@P	SH+ 4@�ӲL�!?��M�o�@7��l�ٿ������@&�|4@@cY�n�!?o�{��o�@7��l�ٿ������@&�|4@@cY�n�!?o�{��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@��o�ٿ�$�&���@~�b��4@���6�!?:�#��o�@����՛ٿ��k��@p־�� 4@u;�9��!?K.�}�o�@����՛ٿ��k��@p־�� 4@u;�9��!?K.�}�o�@����՛ٿ��k��@p־�� 4@u;�9��!?K.�}�o�@����՛ٿ��k��@p־�� 4@u;�9��!?K.�}�o�@����՛ٿ��k��@p־�� 4@u;�9��!?K.�}�o�@���2�ٿ6r�)���@�O�4@�Џ#��!?Eʛ��o�@���2�ٿ6r�)���@�O�4@�Џ#��!?Eʛ��o�@	<*Ć�ٿ�)�_��@�`�N. 4@2�[�i�!?/�o� p�@	<*Ć�ٿ�)�_��@�`�N. 4@2�[�i�!?/�o� p�@	<*Ć�ٿ�)�_��@�`�N. 4@2�[�i�!?/�o� p�@	<*Ć�ٿ�)�_��@�`�N. 4@2�[�i�!?/�o� p�@	<*Ć�ٿ�)�_��@�`�N. 4@2�[�i�!?/�o� p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@cB݇t�ٿx|Q���@J21@��3@9l��g�!?�s
_	p�@�4 �
�ٿ�'�����@�B.� 4@�0�9�!?�'��o�@`�,�ٿ�����@�8��6�3@��;Ԗ�!?�E4p�@`�,�ٿ�����@�8��6�3@��;Ԗ�!?�E4p�@וs�ٿ��O��@�obW�3@{�8ۏ!?��&��o�@����ٿb�$�E��@���uX�3@���d�!?xÄ�(p�@����ٿb�$�E��@���uX�3@���d�!?xÄ�(p�@,s}T!�ٿz!Db���@�O�x4@+gR̯�!?����o�@,s}T!�ٿz!Db���@�O�x4@+gR̯�!?����o�@�����ٿ=ve'��@7�����3@ٺmxÏ!?�l��p�@�����ٿ=ve'��@7�����3@ٺmxÏ!?�l��p�@�I�s��ٿ%��Շ�@��|�=4@AOYGd�!?0��N�o�@�I�s��ٿ%��Շ�@��|�=4@AOYGd�!?0��N�o�@�I�s��ٿ%��Շ�@��|�=4@AOYGd�!?0��N�o�@�V����ٿ ö̇�@<w��4@�#.���!?��U�o�@�V����ٿ ö̇�@<w��4@�#.���!?��U�o�@�V����ٿ ö̇�@<w��4@�#.���!?��U�o�@�V����ٿ ö̇�@<w��4@�#.���!?��U�o�@�V����ٿ ö̇�@<w��4@�#.���!?��U�o�@]~��J�ٿ�av߇�@)5���3@l�j�|�!?���l�o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@���*��ٿ-^
����@6�F��3@(^��=�!?�Q���o�@�1w��ٿ欯<{��@�S؁.�3@gL/��!?��{$�o�@�1w��ٿ欯<{��@�S؁.�3@gL/��!?��{$�o�@����b�ٿ½]���@��t�l�3@�Z+�ȏ!?/�c*�o�@����b�ٿ½]���@��t�l�3@�Z+�ȏ!?/�c*�o�@����b�ٿ½]���@��t�l�3@�Z+�ȏ!?/�c*�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@`ڞb�ٿ�������@3|�K��3@��y,я!?�\�o�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@o��Y՝ٿ�ugT6��@Z��q� 4@Z��;�!?s]�fp�@@�' �ٿ��1��@�7��? 4@�4MT!?�{�p�@�Q�(�ٿ�:�~V��@g����3@.�"��!?��u�o�@�Q�(�ٿ�:�~V��@g����3@.�"��!?��u�o�@�Q�(�ٿ�:�~V��@g����3@.�"��!?��u�o�@�Q�(�ٿ�:�~V��@g����3@.�"��!?��u�o�@��t��ٿq�i���@�٫�4@�/���!?���o�@��t��ٿq�i���@�٫�4@�/���!?���o�@;f�W�ٿQ�C�[��@����<4@�G�e��!?J��(#p�@Rx?�"�ٿ����و�@wY�]}4@���BK�!?�mc�sp�@��ɬ�ٿ_t�+��@z��s4@�5�h�!?��ʣ�p�@��ɬ�ٿ_t�+��@z��s4@�5�h�!?��ʣ�p�@��ɬ�ٿ_t�+��@z��s4@�5�h�!?��ʣ�p�@��ɬ�ٿ_t�+��@z��s4@�5�h�!?��ʣ�p�@�����ٿB��<N��@^:Q�4@���N�!?Jh�$�p�@�����ٿB��<N��@^:Q�4@���N�!?Jh�$�p�@�����ٿB��<N��@^:Q�4@���N�!?Jh�$�p�@�����ٿB��<N��@^:Q�4@���N�!?Jh�$�p�@��p�d�ٿAg���@����^�3@0��\��!?m�h�!q�@��p�d�ٿAg���@����^�3@0��\��!?m�h�!q�@��p�d�ٿAg���@����^�3@0��\��!?m�h�!q�@�L&T��ٿ��Cp��@D#�Ɔ�3@�Q�!͏!?$��3Bp�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@H�3Ꮰٿ������@ΘO��3@�˶Ώ!?S-�0_o�@���3�ٿ��E4���@�V���3@�"x7�!?�/[�q�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@�p9l��ٿ�ᘕ��@=#�� 4@I�ؖ�!?�ȗ8$r�@���S�ٿC�1T��@�$��3@.!��!?����r�@���S�ٿC�1T��@�$��3@.!��!?����r�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@($�[+�ٿh��>���@�o�Z 4@E��S�!?Ú�<�p�@�N����ٿ�}4N��@@���+�3@�12{�!?�5y�=s�@1
�Ф�ٿ��	#���@�[}��4@V�b(��!?�'���t�@1
�Ф�ٿ��	#���@�[}��4@V�b(��!?�'���t�@1
�Ф�ٿ��	#���@�[}��4@V�b(��!?�'���t�@1
�Ф�ٿ��	#���@�[}��4@V�b(��!?�'���t�@ڷi�ٿ2ww+��@�.,c% 4@�l�9׏!?X*�*�t�@ڷi�ٿ2ww+��@�.,c% 4@�l�9׏!?X*�*�t�@ڷi�ٿ2ww+��@�.,c% 4@�l�9׏!?X*�*�t�@�����ٿ8���ܓ�@�$���4@��蛏!?���*w�@�����ٿ8���ܓ�@�$���4@��蛏!?���*w�@�����ٿ8���ܓ�@�$���4@��蛏!?���*w�@�����ٿ8���ܓ�@�$���4@��蛏!?���*w�@�����ٿ8���ܓ�@�$���4@��蛏!?���*w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@pf�<=�ٿ �����@*��e4@��!�ݏ!?o�H�w�@�h���ٿ�n����@��>�94@�Ki��!?�����u�@J20�G�ٿ(
)7��@�~��94@ހ7�x�!?x�*v�@J20�G�ٿ(
)7��@�~��94@ހ7�x�!?x�*v�@J20�G�ٿ(
)7��@�~��94@ހ7�x�!?x�*v�@J20�G�ٿ(
)7��@�~��94@ހ7�x�!?x�*v�@J20�G�ٿ(
)7��@�~��94@ހ7�x�!?x�*v�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@nXZ�њٿ�|H��@��*t:�3@�-�R��!?�DOGw�@�Z#4��ٿ�B9���@.��	�4@!n�qj�!?��9~�@�Z#4��ٿ�B9���@.��	�4@!n�qj�!?��9~�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@'n�8�ٿ�؉�1��@�J��Y�3@r?k܏!?�̭�An�@73�ٿ㉫��@6���4@�鮈�!? ���m�@73�ٿ㉫��@6���4@�鮈�!? ���m�@73�ٿ㉫��@6���4@�鮈�!? ���m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��dk��ٿ�����@�����3@݃8�֏!?9�~��m�@��`�ٿp�@��@l�5�4@�����!?d3�j�@��`�ٿp�@��@l�5�4@�����!?d3�j�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@Y]nG\�ٿ�*�ַ��@��o�Q4@�X<���!?�#�o�@J;!���ٿnι��@:݉��3@:�i��!?���ߔn�@J;!���ٿnι��@:݉��3@:�i��!?���ߔn�@J;!���ٿnι��@:݉��3@:�i��!?���ߔn�@J;!���ٿnι��@:݉��3@:�i��!?���ߔn�@������ٿ���`{�@��y�4@�~y��!?5�nu4h�@�(ˁ�ٿ�r�u�@G,v�4@��ܡ�!?�[�d�@�(ˁ�ٿ�r�u�@G,v�4@��ܡ�!?�[�d�@�(ˁ�ٿ�r�u�@G,v�4@��ܡ�!?�[�d�@m&��פٿ��u�@�A6��3@}w�=�!?C.��Xd�@m&��פٿ��u�@�A6��3@}w�=�!?C.��Xd�@�
n2�ٿ[/N�vg�@e��� 4@�q@�!?��IG\�@�
n2�ٿ[/N�vg�@e��� 4@�q@�!?��IG\�@�
n2�ٿ[/N�vg�@e��� 4@�q@�!?��IG\�@������ٿ$mw���@W��h-4@S�& �!?�CUZ%n�@������ٿ$mw���@W��h-4@S�& �!?�CUZ%n�@������ٿ$mw���@W��h-4@S�& �!?�CUZ%n�@/�$�+�ٿ������@�i|���3@R ah�!?�@+|�@��Ia�ٿ]3���@����3@�UMя!?%�v
p�@��Ia�ٿ]3���@����3@�UMя!?%�v
p�@��Ia�ٿ]3���@����3@�UMя!?%�v
p�@��Ia�ٿ]3���@����3@�UMя!?%�v
p�@��Z��ٿS����@�Y�i� 4@0 'x�!?���Dʅ�@��Z��ٿS����@�Y�i� 4@0 'x�!?���Dʅ�@��g��ٿ�S�r��@`�ʑ4@�y����!?I���މ�@��g��ٿ�S�r��@`�ʑ4@�y����!?I���މ�@��g��ٿ�S�r��@`�ʑ4@�y����!?I���މ�@ؠ�A�ٿ����Ǉ�@-�� 4@c��Oۏ!?�9�k�o�@ؠ�A�ٿ����Ǉ�@-�� 4@c��Oۏ!?�9�k�o�@ؠ�A�ٿ����Ǉ�@-�� 4@c��Oۏ!?�9�k�o�@ؠ�A�ٿ����Ǉ�@-�� 4@c��Oۏ!?�9�k�o�@$&�k�ٿ�6(z�@�lIr&�3@2�P{ď!?/#R��g�@$&�k�ٿ�6(z�@�lIr&�3@2�P{ď!?/#R��g�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@mu�C�ٿݠD]�m�@��	p��3@�c����!?�T�]�_�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@�ZԦ,�ٿ� g�BY�@���=�4@T��W��!?�g�SS�@���+�ٿ�q���n�@g�E��3@մI�ԏ!?��}��`�@���+�ٿ�q���n�@g�E��3@մI�ԏ!?��}��`�@���+�ٿ�q���n�@g�E��3@մI�ԏ!?��}��`�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@�r}�(�ٿHF�.�@�i#� 4@]0��܏!?�a�E9�@g�c�I�ٿ�P`i*��@�h̛��3@�O�R��!?�ٕ����@g�c�I�ٿ�P`i*��@�h̛��3@�O�R��!?�ٕ����@g�c�I�ٿ�P`i*��@�h̛��3@�O�R��!?�ٕ����@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@�Tथ�ٿ*���n��@���d�3@{	�v�!?KЪ�	��@T�b�ٿ��� K;�@��/Y 4@���K�!?:4
A�@n��}�ٿ�<�@�@_�W  4@9B%�q�!??�jo;D�@n��}�ٿ�<�@�@_�W  4@9B%�q�!??�jo;D�@n��}�ٿ�<�@�@_�W  4@9B%�q�!??�jo;D�@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@ƅ̋�ٿ'/9��@�Ҡ��3@p)sH��!?$P8�i��@�E૞ٿ�j���T�@��eC��3@���F��!?l��@�E૞ٿ�j���T�@��eC��3@���F��!?l��@�E૞ٿ�j���T�@��eC��3@���F��!?l��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@r�^�g�ٿ�J>Ͱ�@�~��j�3@��!?��&�a��@�[C�˟ٿ����@��2t��3@PTw��!?�{��U��@�[C�˟ٿ����@��2t��3@PTw��!?�{��U��@X��ٿ�:?�^�@X�s�� 4@\L]�Տ!?�ߣ��V�@X��ٿ�:?�^�@X�s�� 4@\L]�Տ!?�ߣ��V�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@>Oܛٿ���G;�@���*4@c�?t��!?�M�SA�@÷3�F�ٿ]�;�@zd��� 4@G�W���!?]T삘+�@÷3�F�ٿ]�;�@zd��� 4@G�W���!?]T삘+�@÷3�F�ٿ]�;�@zd��� 4@G�W���!?]T삘+�@÷3�F�ٿ]�;�@zd��� 4@G�W���!?]T삘+�@÷3�F�ٿ]�;�@zd��� 4@G�W���!?]T삘+�@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@�,�Ѩٿ7BH���@*~m	��3@��6�z�!?Z�N!��@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@vU{CK�ٿ<������@��R1 4@
���ʏ!?�h�Lv �@s%�5T�ٿ�h�u���@�'U�4@��%�!?K����@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@@�f�ٿ�΃_�@����4@�*�u�!?|n�lX��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@����ήٿ��x��@���4@�d
��!?�0�X��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@c�fǤٿ �@o�@]B� 4@ŭ8透!?�X��A��@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@m���ٿ�&�NR��@�!��8 4@~���Տ!?��b�@�@��h���ٿ,GB����@�>}�? 4@��#��!?�����@��h���ٿ,GB����@�>}�? 4@��#��!?�����@��h���ٿ,GB����@�>}�? 4@��#��!?�����@��h���ٿ,GB����@�>}�? 4@��#��!?�����@��h���ٿ,GB����@�>}�? 4@��#��!?�����@S�'_�ٿ�;��v�@�c����3@�O����!?뷥���@���'�ٿ� ]���@E��� 4@����u�!?�b���@���'�ٿ� ]���@E��� 4@����u�!?�b���@���'�ٿ� ]���@E��� 4@����u�!?�b���@���'�ٿ� ]���@E��� 4@����u�!?�b���@���'�ٿ� ]���@E��� 4@����u�!?�b���@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�S��ٿ�x��C��@$�>���3@�5�2��!?,ȴ�h��@�X󝦙ٿ8�N�z�@{o�v 4@A�=���!?�'��g�@�X󝦙ٿ8�N�z�@{o�v 4@A�=���!?�'��g�@�X󝦙ٿ8�N�z�@{o�v 4@A�=���!?�'��g�@�X󝦙ٿ8�N�z�@{o�v 4@A�=���!?�'��g�@�y�I�ٿ����W#�@��M� 4@.��Ï!?��oH`2�@�y�I�ٿ����W#�@��M� 4@.��Ï!?��oH`2�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@>?u�`�ٿh�8�/�@A�_yR 4@7 z�!?za���9�@U����ٿSl`I���@jX�; 4@��w�C�!?$y��@U����ٿSl`I���@jX�; 4@��w�C�!?$y��@U����ٿSl`I���@jX�; 4@��w�C�!?$y��@U����ٿSl`I���@jX�; 4@��w�C�!?$y��@U����ٿSl`I���@jX�; 4@��w�C�!?$y��@G<?��ٿA�B3T�@��v��3@��a�!?N�vOIP�@����r�ٿ����x�@�����3@b%=x>�!?:Y�4��@����r�ٿ����x�@�����3@b%=x>�!?:Y�4��@����r�ٿ����x�@�����3@b%=x>�!?:Y�4��@����r�ٿ����x�@�����3@b%=x>�!?:Y�4��@���᪜ٿ�7("��@�����3@Τ<�D�!?��lL�@���᪜ٿ�7("��@�����3@Τ<�D�!?��lL�@���᪜ٿ�7("��@�����3@Τ<�D�!?��lL�@�!נٿ�<�j���@~���3@�D�\�!?-��A��@�!נٿ�<�j���@~���3@�D�\�!?-��A��@�!נٿ�<�j���@~���3@�D�\�!?-��A��@���˯�ٿO� Un��@��}�w�3@J>�z�!?S0����@�)\G�ٿM�����@}�?s14@~'�ఏ!?V`v���@�)\G�ٿM�����@}�?s14@~'�ఏ!?V`v���@jb�̤ٿ���P�@���} 4@��ى|�!?�I�JCN�@jb�̤ٿ���P�@���} 4@��ى|�!?�I�JCN�@���A��ٿ�v����@�露��3@��!?�,�p+�@���A��ٿ�v����@�露��3@��!?�,�p+�@���A��ٿ�v����@�露��3@��!?�,�p+�@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��֥��ٿ�Q����@,�4���3@
��Ϗ!?�LE�$��@��b]6�ٿ�г�w��@@h��3@�T@ c�!?�J9H���@��b]6�ٿ�г�w��@@h��3@�T@ c�!?�J9H���@��b]6�ٿ�г�w��@@h��3@�T@ c�!?�J9H���@���Ͱٿ�mKр��@\Ɩ5;�3@�/���!?'i����@���Ͱٿ�mKр��@\Ɩ5;�3@�/���!?'i����@���Ͱٿ�mKр��@\Ɩ5;�3@�/���!?'i����@���Ͱٿ�mKр��@\Ɩ5;�3@�/���!?'i����@���Ͱٿ�mKр��@\Ɩ5;�3@�/���!?'i����@b���ٿa`�5@��@�=,,��3@�1?���!?K9����@b���ٿa`�5@��@�=,,��3@�1?���!?K9����@b���ٿa`�5@��@�=,,��3@�1?���!?K9����@b���ٿa`�5@��@�=,,��3@�1?���!?K9����@�����ٿ�&���@��@� 4@��G��!?�W�~��@�����ٿ�&���@��@� 4@��G��!?�W�~��@�����ٿ�&���@��@� 4@��G��!?�W�~��@�����ٿ�&���@��@� 4@��G��!?�W�~��@�����ٿ�&���@��@� 4@��G��!?�W�~��@�����ٿ�&���@��@� 4@��G��!?�W�~��@(n'���ٿk�E0���@��v� 4@�Zӏ!? 	�˒��@��A!��ٿv2"���@�	F/��3@|�l�!?~�'�#��@��A!��ٿv2"���@�	F/��3@|�l�!?~�'�#��@��A!��ٿv2"���@�	F/��3@|�l�!?~�'�#��@��A!��ٿv2"���@�	F/��3@|�l�!?~�'�#��@�j|��ٿ7'�B�@p�QP��3@�=�U�!??��w�E�@�j|��ٿ7'�B�@p�QP��3@�=�U�!??��w�E�@�j|��ٿ7'�B�@p�QP��3@�=�U�!??��w�E�@�j|��ٿ7'�B�@p�QP��3@�=�U�!??��w�E�@Փ4�ٿ$PJU��@���Y4@��l�!?�B��$�@Փ4�ٿ$PJU��@���Y4@��l�!?�B��$�@Փ4�ٿ$PJU��@���Y4@��l�!?�B��$�@Փ4�ٿ$PJU��@���Y4@��l�!?�B��$�@Փ4�ٿ$PJU��@���Y4@��l�!?�B��$�@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��R��ٿ�l.T��@drtwr�3@�섈�!?���k��@��[���ٿ*I���@J b��3@��(Ï!?d^��X��@/����ٿ/�o7���@ռ��3@U_���!?GȒ%�@��ј�ٿ�6W��@V�:AY4@��7��!?SJ��O�@��ј�ٿ�6W��@V�:AY4@��7��!?SJ��O�@��ј�ٿ�6W��@V�:AY4@��7��!?SJ��O�@��i�ٿJ�e�5:�@5� B�3@Rm�f�!?X��d@�@��i�ٿJ�e�5:�@5� B�3@Rm�f�!?X��d@�@��i�ٿJ�e�5:�@5� B�3@Rm�f�!?X��d@�@��i�ٿJ�e�5:�@5� B�3@Rm�f�!?X��d@�@��i�ٿJ�e�5:�@5� B�3@Rm�f�!?X��d@�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@6�D�J�ٿ�t
���@9j�7��3@�d5��!?$���:�@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@C �ٿV
���@U��4@o�8a��!?Y8ݮ��@��Hȇ�ٿ/�����@�kR4@����{�!?jU~�V��@��Hȇ�ٿ/�����@�kR4@����{�!?jU~�V��@��Hȇ�ٿ/�����@�kR4@����{�!?jU~�V��@Dª���ٿ1��z��@W��4@A�!Q�!?�{���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@�9r���ٿD!,�2��@�2#N� 4@4�[��!?b
���@��d�ٿH�&����@qo�� 4@t�T�!?���Fw��@��d�ٿH�&����@qo�� 4@t�T�!?���Fw��@��d�ٿH�&����@qo�� 4@t�T�!?���Fw��@��d�ٿH�&����@qo�� 4@t�T�!?���Fw��@��d�ٿH�&����@qo�� 4@t�T�!?���Fw��@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@�1{{�ٿ���@-��&
 4@��?��!?���#%�@XcR�ٿ���h���@Ё��	�3@��K�ŏ!?d�����@���*��ٿw��k(��@�#|�3@�ekS��!?������@���*��ٿw��k(��@�#|�3@�ekS��!?������@B��ٿ���ˡV�@�����3@�� y܏!?�k��G��@��I�ٿ"2}����@���N-�3@Gl�_b�!?|�mm��@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�owW�ٿ֑O���@�|�մ�3@Y/�|�!?Z �g�@�W2�Ϟٿ�`
� ��@��pyA�3@����я!?�@�<��@H�$�ٿ�Pۉ���@����4@���랏!?w$�H�
�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@s�.�R�ٿ�n���@�:n��4@pM�O��!?����s&�@�G�J�ٿ{�A�1�@,N��4@��!h�!?ohXC;�@�G�J�ٿ{�A�1�@,N��4@��!h�!?ohXC;�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@��&�5�ٿ<h;M}/�@i���!�3@.BB&��!?b���9�@S�J1�ٿ�,��$�@���^��3@��r���!?����H-�@S�J1�ٿ�,��$�@���^��3@��r���!?����H-�@_��3�ٿ��v����@ߘF>04@�n�͎�!?ɰ�]�@_��3�ٿ��v����@ߘF>04@�n�͎�!?ɰ�]�@_��3�ٿ��v����@ߘF>04@�n�͎�!?ɰ�]�@_��3�ٿ��v����@ߘF>04@�n�͎�!?ɰ�]�@_��3�ٿ��v����@ߘF>04@�n�͎�!?ɰ�]�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@7��#��ٿM�dX7S�@�Ř 4@��ӫ�!?�\�o�O�@ڭL<˦ٿP�;��@NO%��3@hx�Hя!?��\7i��@ڭL<˦ٿP�;��@NO%��3@hx�Hя!?��\7i��@ڭL<˦ٿP�;��@NO%��3@hx�Hя!?��\7i��@ڭL<˦ٿP�;��@NO%��3@hx�Hя!?��\7i��@��a���ٿ���J�@]�霱�3@���ߏ!?2�]J�@�g����ٿe#7��'�@�)�� 4@/�/���!?<9���4�@mV�*��ٿ$Ȯ��@�G��3@@	�$9�!?�ށ!�@�>詸�ٿ(�����@v��k4@ ު��!?/�r.��@�>詸�ٿ(�����@v��k4@ ު��!?/�r.��@����ٿ{��c�w�@�/��)4@��F��!?�E`߭��@����ٿ{��c�w�@�/��)4@��F��!?�E`߭��@iq ��ٿ��~pl��@���4@/1�P��!?� (����@iq ��ٿ��~pl��@���4@/1�P��!?� (����@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�*�tX�ٿ֧d���@��pS�4@ƕ*�֏!?���j��@�ԏ�;�ٿ�zTJ7�@��q�Z 4@���!?�[3�3��@�ԏ�;�ٿ�zTJ7�@��q�Z 4@���!?�[3�3��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@��σߤٿ�9�/.�@� gՖ�3@���ަ�!?�m�.H��@I����ٿ���#��@���˿�3@.	�1��!?�j���@I����ٿ���#��@���˿�3@.	�1��!?�j���@I����ٿ���#��@���˿�3@.	�1��!?�j���@I����ٿ���#��@���˿�3@.	�1��!?�j���@I����ٿ���#��@���˿�3@.	�1��!?�j���@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@���Ȩٿn�W�;$�@K2��#�3@�U}�!?+"=�c��@A9M:��ٿ�R��K�@�����3@��Y}�!?K���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@p��-�ٿ|ј��r�@>�X'4@�:��!?�͜T���@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@>�RwJ�ٿ
�X؇��@C��T��3@�p���!?X�0M|��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@ct��ٿ5�7ar��@�����3@ɦ�h��!?GЄ[K��@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@�>�&%�ٿOz&v,��@�8P��4@�~�x��!?T�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@SP,P�ٿjB���@��n���3@���p��!?�j�����@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@^��l�ٿ� � ���@g>?e�4@�I�AS�!?8�K�Q�@�s�5�ٿPkK�!��@���4@�=f�!?�+���@�s�5�ٿPkK�!��@���4@�=f�!?�+���@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@Z�yB�ٿ�MD4�@��k��3@י����!?� ��,)�@�:!�U�ٿ�AB���@X��4@;��Վ�!?Rj&�g(�@�:!�U�ٿ�AB���@X��4@;��Վ�!?Rj&�g(�@&�*��ٿ�������@��0�)�3@�]ˆ�!?R���9�@&�*��ٿ�������@��0�)�3@�]ˆ�!?R���9�@�	�I�ٿo�w=��@Ei(ݞ�3@�\�L�!?��K7r+�@�	�I�ٿo�w=��@Ei(ݞ�3@�\�L�!?��K7r+�@�	�I�ٿo�w=��@Ei(ݞ�3@�\�L�!?��K7r+�@w�z�[�ٿ�M�Ç�@�����3@��;�!?�%����@w�z�[�ٿ�M�Ç�@�����3@��;�!?�%����@w�z�[�ٿ�M�Ç�@�����3@��;�!?�%����@w�z�[�ٿ�M�Ç�@�����3@��;�!?�%����@f����ٿ�_fā�@Ϣï*�3@zې�u�!?~�� ��@f����ٿ�_fā�@Ϣï*�3@zې�u�!?~�� ��@f����ٿ�_fā�@Ϣï*�3@zې�u�!?~�� ��@f����ٿ�_fā�@Ϣï*�3@zې�u�!?~�� ��@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@:%�`O�ٿ�Hk݃�@wf� 4@ ���ˏ!?�k�u*�@�_����ٿMQ�z�@N��5�3@E7�lʏ!?&CTD.�@�_����ٿMQ�z�@N��5�3@E7�lʏ!?&CTD.�@IAZ<#�ٿ\��B�@)�k$��3@1�[Ϗ!?%�c�*E�@IAZ<#�ٿ\��B�@)�k$��3@1�[Ϗ!?%�c�*E�@IAZ<#�ٿ\��B�@)�k$��3@1�[Ϗ!?%�c�*E�@;�I��ٿ=*�o�d�@���D!�3@�U؟��!?���mYZ�@\����ٿ�g]�~�@��S˗�3@�~7p��!?�ub��@\����ٿ�g]�~�@��S˗�3@�~7p��!?�ub��@\����ٿ�g]�~�@��S˗�3@�~7p��!?�ub��@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@%	�Q��ٿ9�
 ���@C_�� 4@�7���!?(�����@�����ٿْv����@%~cL@�3@��Z`�!?"��TS��@�����ٿْv����@%~cL@�3@��Z`�!?"��TS��@�����ٿْv����@%~cL@�3@��Z`�!?"��TS��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@�``�S�ٿ�v�yt�@�y�a�3@`=�ӑ�!?�c��A��@F(4�ٿ@���u��@ت�Ue�3@���H��!?>p=��@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@���)��ٿ�P��@� 4@��L��!?�S'��	�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@$���ٿ�V�@_nh��3@:h���!?�^�X!�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@H��V��ٿ��~b��@���2�3@5�F1��!?:���#�@%�Y�8�ٿ�Ef�@]�͛[�3@��=�!?�n.g\��@�$��!�ٿ��l���@�K� 4@c.���!?��+��@�$��!�ٿ��l���@�K� 4@c.���!?��+��@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@��i�F�ٿ�8�����@fح'4@8����!?�ޫ����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@E��E��ٿ�g$S��@�l�G+4@�� m{�!?IG�����@��=���ٿ�c�����@�Xf�3@NZo��!?�4��_�@��=���ٿ�c�����@�Xf�3@NZo��!?�4��_�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�7���ٿ>�x��@��� | 4@�E��!?~/f
�@�Ƴ�ٿ�5s���@5�����3@�,�͐�!?������@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@*D{ʗٿ��-�>�@ד�4@Fh���!?s<뷧A�@𥳐�خٿ����@h&4-r�3@�|~��!?�[{���@Vnk��ٿÓ�g'�@3|)��3@Iz��!?<੔�1�@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@bj���ٿfo�y��@�{�[� 4@���>��!?ky�2^��@�O�ކ�ٿ9TA�Ȅ�@������3@p�	�x�!?��L���@�O�ކ�ٿ9TA�Ȅ�@������3@p�	�x�!?��L���@�O�ކ�ٿ9TA�Ȅ�@������3@p�	�x�!?��L���@�o��ٿۓ9���@
\c���3@�g3��!?Ʊ����@�o��ٿۓ9���@
\c���3@�g3��!?Ʊ����@�o��ٿۓ9���@
\c���3@�g3��!?Ʊ����@B��$v�ٿhg(��@������3@��zd�!?�b�!�@B��$v�ٿhg(��@������3@��zd�!?�b�!�@ [�j��ٿ�2ّ�.�@�&�� 4@C
��Q�!?��=j1�@ [�j��ٿ�2ّ�.�@�&�� 4@C
��Q�!?��=j1�@ [�j��ٿ�2ّ�.�@�&�� 4@C
��Q�!?��=j1�@ [�j��ٿ�2ّ�.�@�&�� 4@C
��Q�!?��=j1�@=�ކ��ٿ��g'���@�{
o�4@}J��!?UE1��@=�ކ��ٿ��g'���@�{
o�4@}J��!?UE1��@=�ކ��ٿ��g'���@�{
o�4@}J��!?UE1��@=�ކ��ٿ��g'���@�{
o�4@}J��!?UE1��@t&��ٿֿ����@�fb�� 4@���A�!?U�>H���@t&��ٿֿ����@�fb�� 4@���A�!?U�>H���@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@]qe�ٿ�ԩ��@y�"� 4@�U�B��!?mb��M��@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@͠e6��ٿ�����@�]�� 4@~���ݏ!?��C[�	�@�q얥ٿ�8m�w�@k�3&�3@�<J{��!?Wg�C��@OZ�\��ٿE����@�!���3@�0߼��!?:
h���@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@��(�̟ٿGQ�R���@,OH2h�3@�~^��!?8\�@�7c�L�ٿݰ� ��@zrWi�3@9I���!?65N�c��@�7c�L�ٿݰ� ��@zrWi�3@9I���!?65N�c��@�7c�L�ٿݰ� ��@zrWi�3@9I���!?65N�c��@�7c�L�ٿݰ� ��@zrWi�3@9I���!?65N�c��@�I���ٿ��	�"�@�R�c�3@��h�ˏ!?����>�@Q�*�Ϩٿ⻪�x(�@U;N��3@e�]��!?-�2��=�@Q�*�Ϩٿ⻪�x(�@U;N��3@e�]��!?-�2��=�@Q�*�Ϩٿ⻪�x(�@U;N��3@e�]��!?-�2��=�@�\z�b�ٿ0�����@��%� 4@��<���!?ֶdq���@�\z�b�ٿ0�����@��%� 4@��<���!?ֶdq���@�\z�b�ٿ0�����@��%� 4@��<���!?ֶdq���@�\z�b�ٿ0�����@��%� 4@��<���!?ֶdq���@�\z�b�ٿ0�����@��%� 4@��<���!?ֶdq���@��hJ:�ٿ�ϛ�@��b���3@�9a�s�!?:[LE��@��hJ:�ٿ�ϛ�@��b���3@�9a�s�!?:[LE��@�/!�|�ٿ�Q�!���@t[��3@�.MEK�!?>zp��@�/!�|�ٿ�Q�!���@t[��3@�.MEK�!?>zp��@h���z�ٿ���?�@c�����3@jav���!?�F���@h���z�ٿ���?�@c�����3@jav���!?�F���@h���z�ٿ���?�@c�����3@jav���!?�F���@h���z�ٿ���?�@c�����3@jav���!?�F���@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@_Q���ٿu���c�@������3@G�;��!?��3�>�@���K	�ٿ�IWܣ�@*[��Y 4@ƇF ��!?��^qh��@���K	�ٿ�IWܣ�@*[��Y 4@ƇF ��!?��^qh��@���K	�ٿ�IWܣ�@*[��Y 4@ƇF ��!?��^qh��@���K	�ٿ�IWܣ�@*[��Y 4@ƇF ��!?��^qh��@���K	�ٿ�IWܣ�@*[��Y 4@ƇF ��!?��^qh��@��1CL�ٿE!� *�@����� 4@)2ʂ�!?C��={�@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�6�j�ٿ��S��@d�B4@$|�ӏ!?�^l��@�VEf�ٿ�F��Ɏ�@�m�$� 4@��L���!?��3���@ �O���ٿ���1Y��@FG�� 4@!��ݏ!?es�P��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@9�s�ٿ�-!K��@KL"�^�3@4�~f��!?��6�1��@���H�ٿ�jW��@�φug 4@4X���!?�Cm���@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@�?��/�ٿB��S���@�;�4@_�b�ԏ!?ŢNڤ��@	>�;�ٿ��o#���@�dC��3@~Z*5��!?���<��@mQHez�ٿ�'Q�pz�@y�"�& 4@�U��ޏ!?���w�&�@mQHez�ٿ�'Q�pz�@y�"�& 4@�U��ޏ!?���w�&�@mQHez�ٿ�'Q�pz�@y�"�& 4@�U��ޏ!?���w�&�@mQHez�ٿ�'Q�pz�@y�"�& 4@�U��ޏ!?���w�&�@2i�JǙٿ����%��@�����3@�Z�g.�!?��^��Z�@2i�JǙٿ����%��@�����3@�Z�g.�!?��^��Z�@�$#5�ٿ��$��u�@�g3�4@+I�z�!?�C4m���@�$#5�ٿ��$��u�@�g3�4@+I�z�!?�C4m���@�$#5�ٿ��$��u�@�g3�4@+I�z�!?�C4m���@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@�	�V�ٿTH�� �@��gm4@]j׏!?�\�r��@
a�R�ٿ�* �'�@�����3@��׿�!?O�((�@
a�R�ٿ�* �'�@�����3@��׿�!?O�((�@]ϰ�ٿ6[�[#�@�`����3@�I̏!?�3�3)-�@�]�&o�ٿ�7�_Ѓ�@�� ?��3@�nC?��!?L(�FP�@�]�&o�ٿ�7�_Ѓ�@�� ?��3@�nC?��!?L(�FP�@[1�p�ٿm$E�o)�@���3@������!?�,`c(�@@�����ٿ������@?=6�� 4@��z��!?�������@@�����ٿ������@?=6�� 4@��z��!?�������@@�����ٿ������@?=6�� 4@��z��!?�������@@�����ٿ������@?=6�� 4@��z��!?�������@@�����ٿ������@?=6�� 4@��z��!?�������@@�����ٿ������@?=6�� 4@��z��!?�������@���vu�ٿ������@��Nio�3@�Tmy��!?�����@}w�ٿ�� r�C�@��=4@r\AϏ!?�R�~�<�@�7=�ۦٿ���:�@!�M��3@{�q䎏!?��(P9�@�7=�ۦٿ���:�@!�M��3@{�q䎏!?��(P9�@9��O��ٿ�_z����@�Ֆq4@k7�Eq�!?�դ�W��@9��O��ٿ�_z����@�Ֆq4@k7�Eq�!?�դ�W��@9��O��ٿ�_z����@�Ֆq4@k7�Eq�!?�դ�W��@9��O��ٿ�_z����@�Ֆq4@k7�Eq�!?�դ�W��@9��O��ٿ�_z����@�Ֆq4@k7�Eq�!?�դ�W��@���B��ٿ�� �//�@��U�� 4@'���!?p@W��v�@���B��ٿ�� �//�@��U�� 4@'���!?p@W��v�@���B��ٿ�� �//�@��U�� 4@'���!?p@W��v�@���B��ٿ�� �//�@��U�� 4@'���!?p@W��v�@���5��ٿ����@�X"4@J0��3�!?�DO�c��@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@e�\��ٿTѫ���@�ԗ��4@Rt8橏!?E)�He�@���N�ٿ?�T����@�yNR4@6��O�!?:4�۬�@���N�ٿ?�T����@�yNR4@6��O�!?:4�۬�@���N�ٿ?�T����@�yNR4@6��O�!?:4�۬�@���N�ٿ?�T����@�yNR4@6��O�!?:4�۬�@E�pi�ٿ��\�@S��� 4@��}ʏ!?�L�\ǻ�@E�pi�ٿ��\�@S��� 4@��}ʏ!?�L�\ǻ�@E�pi�ٿ��\�@S��� 4@��}ʏ!?�L�\ǻ�@E�pi�ٿ��\�@S��� 4@��}ʏ!?�L�\ǻ�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@͕o�!�ٿV��ʄ��@t�kۂ 4@SZY��!?��` �z�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@�綻��ٿ�5�����@�L�ޟ4@���ɐ�!?��\��F�@����ٿ{��ۚ��@4�j 4@tӀ�!? �dd�@����ٿ{��ۚ��@4�j 4@tӀ�!? �dd�@�Q8�Ѭٿm������@~����3@x ��!?�{����@�Q8�Ѭٿm������@~����3@x ��!?�{����@�Q8�Ѭٿm������@~����3@x ��!?�{����@6b"Ȼ�ٿ+y��L��@�5�) 4@�$V5�!?�ǜb�"�@6b"Ȼ�ٿ+y��L��@�5�) 4@�$V5�!?�ǜb�"�@I���ϛٿg�h�@�
��.4@oG�U�!?�>a�j��@I���ϛٿg�h�@�
��.4@oG�U�!?�>a�j��@I���ϛٿg�h�@�
��.4@oG�U�!?�>a�j��@n��M�ٿ��"��@�I�!�3@��u�!?"�;Kf�@@����ٿ����c��@tj!$� 4@.��G��!?�i1:a��@@����ٿ����c��@tj!$� 4@.��G��!?�i1:a��@@����ٿ����c��@tj!$� 4@.��G��!?�i1:a��@@����ٿ����c��@tj!$� 4@.��G��!?�i1:a��@_��b�ٿIԣ����@nCQ( 4@���䀏!?���?�^�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@�w��ٿ4Y�V�@��*���3@U3#�=�!?�j<n�@��(��ٿvD�W��@�(�y�3@z5�G��!?|���Q�@��(��ٿvD�W��@�(�y�3@z5�G��!?|���Q�@��(��ٿvD�W��@�(�y�3@z5�G��!?|���Q�@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@����ٿ7�!�q�@R���v�3@5v��!?�ӂ�c��@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@���V�ٿ
�Bؚ�@}Ħ;��3@g�躏!?̪���@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@�V����ٿ�Bn���@|���3@��d���!?��.(:��@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@e@%�ٿB����@[� 4@}2EV��!?٦�t�@O�ܫٿ`�^���@��t� 4@���'��!?^�}�xD�@O�ܫٿ`�^���@��t� 4@���'��!?^�}�xD�@O�ܫٿ`�^���@��t� 4@���'��!?^�}�xD�@O�ܫٿ`�^���@��t� 4@���'��!?^�}�xD�@O�ܫٿ`�^���@��t� 4@���'��!?^�}�xD�@�1��y�ٿq��ث�@qԳs4@Rs��!?���L@��@�1��y�ٿq��ث�@qԳs4@Rs��!?���L@��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@ǉzäٿ� ��A�@d��o94@��I!?��BLk��@�>;�ڭٿ��0��@I�h�] 4@�M檑�!?�3�i��@�>;�ڭٿ��0��@I�h�] 4@�M檑�!?�3�i��@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@���o*�ٿ������@}.�C� 4@C�G_��!?�s\���@�_�=שٿڋ�x���@o�m�� 4@u�cF��!?u}��A �@�_�=שٿڋ�x���@o�m�� 4@u�cF��!?u}��A �@l@,��ٿ�u��]�@�Mkk�4@mܖ���!?א�����@l@,��ٿ�u��]�@�Mkk�4@mܖ���!?א�����@l@,��ٿ�u��]�@�Mkk�4@mܖ���!?א�����@l@,��ٿ�u��]�@�Mkk�4@mܖ���!?א�����@l@,��ٿ�u��]�@�Mkk�4@mܖ���!?א�����@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@�ڗ�D�ٿ9o��q��@NN� 4@����!?i�,9��@[?ÐG�ٿ9л]���@{lS�N4@w�S�!?�'�sR�@�Ks���ٿ�xS���@���(4@	/D"��!?��Þ�@�Ks���ٿ�xS���@���(4@	/D"��!?��Þ�@�Ks���ٿ�xS���@���(4@	/D"��!?��Þ�@�Ks���ٿ�xS���@���(4@	/D"��!?��Þ�@�#�>3�ٿ\�����@�@�J 4@p��m�!?�ġpׄ�@�S����ٿ~˛�֢�@���� 4@l��wk�!?�@�L�@y3�w�ٿ�����@���p/4@�d��m�!?(�y�+�@y3�w�ٿ�����@���p/4@�d��m�!?(�y�+�@n��:�ٿk_p����@M\��24@}\�&�!?��ׁ��@n��:�ٿk_p����@M\��24@}\�&�!?��ׁ��@�p��̡ٿ��)c+�@�1Ր�4@Za6D�!?eڻ.�j�@���M[�ٿK�;v��@�x�<4@�l�4��!?�6܌z2�@���M[�ٿK�;v��@�x�<4@�l�4��!?�6܌z2�@Z� S�ٿ��.,�U�@g>�
\4@��L�\�!?���^a�@Z� S�ٿ��.,�U�@g>�
\4@��L�\�!?���^a�@Z� S�ٿ��.,�U�@g>�
\4@��L�\�!?���^a�@��اڢٿ���Ԏr�@7F}�3�3@��7�h�!?Ϩ���T�@��اڢٿ���Ԏr�@7F}�3�3@��7�h�!?Ϩ���T�@��اڢٿ���Ԏr�@7F}�3�3@��7�h�!?Ϩ���T�@��اڢٿ���Ԏr�@7F}�3�3@��7�h�!?Ϩ���T�@��اڢٿ���Ԏr�@7F}�3�3@��7�h�!?Ϩ���T�@^0:��ٿ2��A׍�@��@�.�3@,���E�!?����1��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@O	�+��ٿ<`%E^�@t��)��3@�^JYG�!?>�G��@�Wv�+�ٿEPh��@<?���3@��L��!?�k\v[6�@M���٠ٿ�(�".�@��&��3@>ߘ�!?�֫/�U�@M���٠ٿ�(�".�@��&��3@>ߘ�!?�֫/�U�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@'>�(ԗٿt��x(��@W�� 4@%Ls�B�!?פ<ЙJ�@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@zMLZ��ٿ�����@�:�&��3@�?�Մ�!?$�d �@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@�3&6�ٿD��r3��@�H<X�3@��zA��!?��r��@<X��ٿ���!u�@hƙE��3@���|{�!?'ԍ��@<X��ٿ���!u�@hƙE��3@���|{�!?'ԍ��@<X��ٿ���!u�@hƙE��3@���|{�!?'ԍ��@<X��ٿ���!u�@hƙE��3@���|{�!?'ԍ��@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@��9J�ٿh������@a��>4@Z���Џ!?| �Ȇk�@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@�Fаm�ٿ���@��,�4@�;�k��!?�6���@������ٿ�bVZ���@T���3@#�g:\�!?�"2����@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@Ne�ٿ��tq�@B,T��3@f��l�!?�������@���9�ٿŉ_���@� G��3@8),Ò�!?ۧ��y�@���9�ٿŉ_���@� G��3@8),Ò�!?ۧ��y�@���9�ٿŉ_���@� G��3@8),Ò�!?ۧ��y�@���9�ٿŉ_���@� G��3@8),Ò�!?ۧ��y�@j��g=�ٿsS���@S,����3@��Bȏ!??bax��@8:5�ʞٿ�y8OG�@���A��3@�l-��!?ȋ�����@8:5�ʞٿ�y8OG�@���A��3@�l-��!?ȋ�����@���ٿ�ǐد%�@Q����3@P�e��!?$X;|ޚ�@���ٿ�ǐد%�@Q����3@P�e��!?$X;|ޚ�@��w���ٿ�8q����@(	�5��3@������!?��L���@��w���ٿ�8q����@(	�5��3@������!?��L���@��w���ٿ�8q����@(	�5��3@������!?��L���@��w���ٿ�8q����@(	�5��3@������!?��L���@��w���ٿ�8q����@(	�5��3@������!?��L���@��w���ٿ�8q����@(	�5��3@������!?��L���@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@-N[˱ٿd�%S���@�!З* 4@�z�܏!?j��G�@8!�|�ٿ���>+�@G�m�� 4@�!$ Y�!?C���)i�@8!�|�ٿ���>+�@G�m�� 4@�!$ Y�!?C���)i�@8!�|�ٿ���>+�@G�m�� 4@�!$ Y�!?C���)i�@K�ߕ�ٿ$��K�n�@�G�<�3@mM�K�!?�2�,��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@$+�M�ٿ?a+e�@����I�3@3��d�!?�w�p��@�@ʝ
�ٿ�놦��@�Q�A4@�E;��!?�B��e�@���ٿ�̛�a��@���.64@@���!?��ఉ~�@���ٿ�̛�a��@���.64@@���!?��ఉ~�@���ٿ�̛�a��@���.64@@���!?��ఉ~�@���ٿ�̛�a��@���.64@@���!?��ఉ~�@���ٿ�̛�a��@���.64@@���!?��ఉ~�@�k�.C�ٿ����8�@��R�H 4@U�L�!?�o�d0��@�k�.C�ٿ����8�@��R�H 4@U�L�!?�o�d0��@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�f�a�ٿ�/~����@!�2� 4@ȴ�|E�!?���_�@�5�ٿ�C����@�t����3@
V�޷�!?pvf@���@�5�ٿ�C����@�t����3@
V�޷�!?pvf@���@�5�ٿ�C����@�t����3@
V�޷�!?pvf@���@�5�ٿ�C����@�t����3@
V�޷�!?pvf@���@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@�[E�ٿ�k�#���@�Y̪�3@��	�Ə!??k�j�F�@C̝���ٿ��;蚭�@�w˛S�3@��߬�!?�e��~�@q0����ٿ�|�p�@EF��[ 4@;�l@��!?-�E�q�@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@21O��ٿi!B'C�@�&-��3@�tu0Ə!?d\e�P��@tǣ*/�ٿ�9B�Py�@͗X�U 4@nݤM�!?/�lOk��@tǣ*/�ٿ�9B�Py�@͗X�U 4@nݤM�!?/�lOk��@tǣ*/�ٿ�9B�Py�@͗X�U 4@nݤM�!?/�lOk��@tǣ*/�ٿ�9B�Py�@͗X�U 4@nݤM�!?/�lOk��@tǣ*/�ٿ�9B�Py�@͗X�U 4@nݤM�!?/�lOk��@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@��F3T�ٿ�LYhl��@]�
6y�3@I�$�F�!?;]L���@�,$��ٿ|�ϬW�@�^ �| 4@�骂"�!?�Y�^.��@�,$��ٿ|�ϬW�@�^ �| 4@�骂"�!?�Y�^.��@�,$��ٿ|�ϬW�@�^ �| 4@�骂"�!?�Y�^.��@׿	:�ٿ_��x���@*<|9�3@G��?�!?&���B�@׿	:�ٿ_��x���@*<|9�3@G��?�!?&���B�@׿	:�ٿ_��x���@*<|9�3@G��?�!?&���B�@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@
����ٿ��g׆�@�zN`9�3@[�`Z�!?�,/-���@i��A^�ٿ1��e�-�@���w�3@1ԯRX�!?X�Bv�@i��A^�ٿ1��e�-�@���w�3@1ԯRX�!?X�Bv�@i��A^�ٿ1��e�-�@���w�3@1ԯRX�!?X�Bv�@i��A^�ٿ1��e�-�@���w�3@1ԯRX�!?X�Bv�@i��A^�ٿ1��e�-�@���w�3@1ԯRX�!?X�Bv�@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@{ �o�ٿ�z9X�X�@�vR���3@�ٖ��!?3�A���@��&��ٿ؍^�ł�@�/�*�3@�v��!?V=y�Ҵ�@��&��ٿ؍^�ł�@�/�*�3@�v��!?V=y�Ҵ�@��&��ٿ؍^�ł�@�/�*�3@�v��!?V=y�Ҵ�@��&��ٿ؍^�ł�@�/�*�3@�v��!?V=y�Ҵ�@N���ٿ$���ٗ�@J< i��3@<47ﳏ!?Th�;i�@N���ٿ$���ٗ�@J< i��3@<47ﳏ!?Th�;i�@N���ٿ$���ٗ�@J< i��3@<47ﳏ!?Th�;i�@N���ٿ$���ٗ�@J< i��3@<47ﳏ!?Th�;i�@��Gb�ٿ��(��@�d ���3@���y�!?U��0�@��Gb�ٿ��(��@�d ���3@���y�!?U��0�@��Gb�ٿ��(��@�d ���3@���y�!?U��0�@J�=U�ٿC�8���@M_H�`4@T+�sď!?��i���@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@ōxO�ٿjL�\�@/�&,�4@ԏ�ټ�!??�<"o��@T���ٿ������@���Y�4@��.8��!?�36i]�@ʬ6H٢ٿ�� ��@-R�6�3@���&_�!?ђԠ�(�@!9��ٿ��M]d��@���)� 4@�"#��!?'��(`�@!9��ٿ��M]d��@���)� 4@�"#��!?'��(`�@!9��ٿ��M]d��@���)� 4@�"#��!?'��(`�@!9��ٿ��M]d��@���)� 4@�"#��!?'��(`�@l!�8��ٿj�i=��@���_m4@��.t�!?�v�j��@l!�8��ٿj�i=��@���_m4@��.t�!?�v�j��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@��S̰�ٿ�׳L��@���4@���픏!?!k毌��@M4�?�ٿ�W*C%�@w;�{ 4@�]���!?�6v�6��@M4�?�ٿ�W*C%�@w;�{ 4@�]���!?�6v�6��@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�a�b0�ٿV�{N7��@mh�� �3@:�+���!?9K�����@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@�fb�ٿ�V_4��@ �v�Z 4@y���!?�eb>�l�@��؂_�ٿg�Co���@�d�4@|��\W�!??o'~�@��؂_�ٿg�Co���@�d�4@|��\W�!??o'~�@ԅ9	u�ٿ8�F���@�U~�4@H��P�!?�(��'�@ԅ9	u�ٿ8�F���@�U~�4@H��P�!?�(��'�@�m����ٿ�w����@��l�4@A�g�	�!?���}�@�m����ٿ�w����@��l�4@A�g�	�!?���}�@ MZ(��ٿJ�- ��@�M_�%4@�p�ɏ!?��F`̰�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@��q7�ٿ�� s�9�@��m+4@�CT:ۏ!?RSU��O�@�ląٿ�B#�9��@�J=4@gM&ˏ!?R�ۣ�@�ląٿ�B#�9��@�J=4@gM&ˏ!?R�ۣ�@�}̘�ٿ�_D��@&��3�4@�=���!?ϟ�R~4�@�}̘�ٿ�_D��@&��3�4@�=���!?ϟ�R~4�@�}̘�ٿ�_D��@&��3�4@�=���!?ϟ�R~4�@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�I�'�ٿ�J����@�� l��3@�u�_�!?�f�=��@�e�z�ٿ��:���@Qp`�] 4@�}iS�!?���-��@�e�z�ٿ��:���@Qp`�] 4@�}iS�!?���-��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@�Z:�
�ٿ��-�@��K-4@C�����!?��>�o��@"�ݡ�ٿ�5��@PQ%�4@�Pv�!?����SU�@"�ݡ�ٿ�5��@PQ%�4@�Pv�!?����SU�@"�ݡ�ٿ�5��@PQ%�4@�Pv�!?����SU�@"�ݡ�ٿ�5��@PQ%�4@�Pv�!?����SU�@f|O�\�ٿA(���_�@I}���3@�FD�y�!?�Ǩ#Π�@f|O�\�ٿA(���_�@I}���3@�FD�y�!?�Ǩ#Π�@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@�]*L�ٿ�F۱n��@�����3@��{��!?��g��@��%E�ٿ'K���@.J�4@3\'���!?K�a֍��@��%E�ٿ'K���@.J�4@3\'���!?K�a֍��@��%E�ٿ'K���@.J�4@3\'���!?K�a֍��@��%E�ٿ'K���@.J�4@3\'���!?K�a֍��@��%E�ٿ'K���@.J�4@3\'���!?K�a֍��@�1^Ƭٿ0DcD��@�����4@��R��!?6�W���@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�m]��ٿ���8��@U"}4@�I�Ϣ�!?��Ee�>�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�7m2�ٿ �X0���@ݵ��/ 4@�X􅎏!?`?n�4�@�N�IK�ٿY��م��@�f�[g4@N~	�ݏ!?A�u�>�@�N�IK�ٿY��م��@�f�[g4@N~	�ݏ!?A�u�>�@�N�IK�ٿY��م��@�f�[g4@N~	�ݏ!?A�u�>�@��ŵ��ٿ�Iݤ�@����4@�2;���!?ND��h�@��ŵ��ٿ�Iݤ�@����4@�2;���!?ND��h�@��ŵ��ٿ�Iݤ�@����4@�2;���!?ND��h�@��ŵ��ٿ�Iݤ�@����4@�2;���!?ND��h�@�٦xv�ٿ�-�{�@P4b@4@�_�{�!?�m�i�J�@�٦xv�ٿ�-�{�@P4b@4@�_�{�!?�m�i�J�@�٦xv�ٿ�-�{�@P4b@4@�_�{�!?�m�i�J�@�٦xv�ٿ�-�{�@P4b@4@�_�{�!?�m�i�J�@�٦xv�ٿ�-�{�@P4b@4@�_�{�!?�m�i�J�@�n�{�ٿ��}D_�@��5B�4@,"\`��!?�_���@�V�-x�ٿ��ht��@*�&�'4@�ӊ��!?h�����@�V�-x�ٿ��ht��@*�&�'4@�ӊ��!?h�����@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�-���ٿF�8D��@��4@k�cL��!?E��@�t��u�ٿ8���l�@ǀM`4@^D�T؏!?*���@�t��u�ٿ8���l�@ǀM`4@^D�T؏!?*���@�t��u�ٿ8���l�@ǀM`4@^D�T؏!?*���@��Z%��ٿ�fN���@�G��2 4@Ԡ=x��!?a��D���@��Z%��ٿ�fN���@�G��2 4@Ԡ=x��!?a��D���@��Z%��ٿ�fN���@�G��2 4@Ԡ=x��!?a��D���@��Z%��ٿ�fN���@�G��2 4@Ԡ=x��!?a��D���@��Z%��ٿ�fN���@�G��2 4@Ԡ=x��!?a��D���@ַ�R]�ٿ����6��@	�=�*4@ǔ7.��!?פ.��
�@ַ�R]�ٿ����6��@	�=�*4@ǔ7.��!?פ.��
�@ַ�R]�ٿ����6��@	�=�*4@ǔ7.��!?פ.��
�@��cq�ٿ����y��@��zz��3@].��~�!?e �J��@BP[qF�ٿ��-��@���^ 4@N�ꛏ!?�3J_���@BP[qF�ٿ��-��@���^ 4@N�ꛏ!?�3J_���@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�V�ٿ'������@�0b���3@�(Ǔ�!?�.~j_��@�3�ٿ%���Վ�@<����3@c}��Ϗ!?�18�r�@�3�ٿ%���Վ�@<����3@c}��Ϗ!?�18�r�@�3�ٿ%���Վ�@<����3@c}��Ϗ!?�18�r�@�H���ٿ-2 �y�@�U��.�3@�y�T��!?��7|��@�H���ٿ-2 �y�@�U��.�3@�y�T��!?��7|��@�H���ٿ-2 �y�@�U��.�3@�y�T��!?��7|��@�H���ٿ-2 �y�@�U��.�3@�y�T��!?��7|��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@W���?�ٿ+oX2y�@���+�3@�ܺ�x�!?�t�l��@����ٿ�K �m�@y7|u�3@c��P�!?�c�t{,�@��Kh�ٿ��R���@ j���3@^��y�!?u%瀷�@��Kh�ٿ��R���@ j���3@^��y�!?u%瀷�@P2u�1�ٿ�Q���'�@��,��3@�K�g��!?�c*6���@@ύs��ٿ�#�@ZZ�@1���J 4@/���Ə!?cƇ����@}��w(�ٿ��3˯��@�e�ff 4@#����!?<�����@}��w(�ٿ��3˯��@�e�ff 4@#����!?<�����@��U�)�ٿ����mL�@m֫I� 4@%A3���!?�ϯ�B�@��U�)�ٿ����mL�@m֫I� 4@%A3���!?�ϯ�B�@��U�)�ٿ����mL�@m֫I� 4@%A3���!?�ϯ�B�@��U�)�ٿ����mL�@m֫I� 4@%A3���!?�ϯ�B�@��U�)�ٿ����mL�@m֫I� 4@%A3���!?�ϯ�B�@��c�ٿAb.,��@��٩� 4@�mr��!?�Hq�>��@��c�ٿAb.,��@��٩� 4@�mr��!?�Hq�>��@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@!i���ٿ	�KPҦ�@>�.4@�H�#��!?��h:6�@�dQ���ٿ� w�t�@������3@i�V���!?h�*�c��@{�a� �ٿÄE���@�^�S�3@��Ï!?O&�2�@{�a� �ٿÄE���@�^�S�3@��Ï!?O&�2�@{�a� �ٿÄE���@�^�S�3@��Ï!?O&�2�@{�a� �ٿÄE���@�^�S�3@��Ï!?O&�2�@̭F�,�ٿ�����@��<w 4@Wǿϻ�!?R��2?�@̭F�,�ٿ�����@��<w 4@Wǿϻ�!?R��2?�@��ե��ٿg]E�
v�@zz��< 4@����m�!?:���Gs�@��ե��ٿg]E�
v�@zz��< 4@����m�!?:���Gs�@��ե��ٿg]E�
v�@zz��< 4@����m�!?:���Gs�@��P�ٿ����@ʸ�{� 4@\}��!?�[��3N�@��P�ٿ����@ʸ�{� 4@\}��!?�[��3N�@��P�ٿ����@ʸ�{� 4@\}��!?�[��3N�@��P�ٿ����@ʸ�{� 4@\}��!?�[��3N�@��P�ٿ����@ʸ�{� 4@\}��!?�[��3N�@=�w�ٿ�����@Ɉ;�4@�}g�!?@ޡ����@=�w�ٿ�����@Ɉ;�4@�}g�!?@ޡ����@=�w�ٿ�����@Ɉ;�4@�}g�!?@ޡ����@=�w�ٿ�����@Ɉ;�4@�}g�!?@ޡ����@=�w�ٿ�����@Ɉ;�4@�}g�!?@ޡ����@��1Y�ٿ�C&�F�@PgF(��3@<8Ʌ��!?]|��b�@��1Y�ٿ�C&�F�@PgF(��3@<8Ʌ��!?]|��b�@��1Y�ٿ�C&�F�@PgF(��3@<8Ʌ��!?]|��b�@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@A�#h��ٿ���r=h�@}n-�4 4@��BLɏ!?o�f�x��@m_��ٿZ�l��J�@��M/��3@��ˏ!?�SM����@m_��ٿZ�l��J�@��M/��3@��ˏ!?�SM����@����ٿD��l�@�./��3@�|}��!?�3aŌ�@����ٿD��l�@�./��3@�|}��!?�3aŌ�@����ٿD��l�@�./��3@�|}��!?�3aŌ�@����ٿD��l�@�./��3@�|}��!?�3aŌ�@7��V��ٿH=-p\�@d��)� 4@L,�Ə!?�'*
u�@7��V��ٿH=-p\�@d��)� 4@L,�Ə!?�'*
u�@7��V��ٿH=-p\�@d��)� 4@L,�Ə!?�'*
u�@o�밟ٿ�M�t�@� b���3@��y���!?龻���@o�밟ٿ�M�t�@� b���3@��y���!?龻���@�}�ʫٿ��N��@��f3" 4@Hs@���!?��D_��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@�=u�x�ٿ(�5���@B<;���3@�%~��!?�1��Y��@(��dQ�ٿY^�^�}�@��@SP�3@�ޗ�܏!?��C�.y�@�����ٿ��W�h��@���_�3@�����!?,�6�Xf�@�����ٿ��W�h��@���_�3@�����!?,�6�Xf�@�����ٿ��W�h��@���_�3@�����!?,�6�Xf�@�����ٿ��W�h��@���_�3@�����!?,�6�Xf�@�����ٿ��W�h��@���_�3@�����!?,�6�Xf�@x}H��ٿ8q���P�@��{+g�3@G
y���!?m�>k�@���$p�ٿyf��n�@ߌ�m� 4@X`?Х�!?d#{B��@F~��ڢٿ_m�$���@s�Q4@r�t���!?�_�n���@F~��ڢٿ_m�$���@s�Q4@r�t���!?�_�n���@F~��ڢٿ_m�$���@s�Q4@r�t���!?�_�n���@F~��ڢٿ_m�$���@s�Q4@r�t���!?�_�n���@F~��ڢٿ_m�$���@s�Q4@r�t���!?�_�n���@�U�-�ٿ�˪no�@��B�4@��;7؏!?ld-8�@�U�-�ٿ�˪no�@��B�4@��;7؏!?ld-8�@f��*)�ٿT��F��@#<���3@v����!?�0E�se�@9*;���ٿ�GVt���@CϮ�� 4@_�Xz-�!?	Z
���@j��D �ٿF�Z�s��@�}�) 4@����!?�3�G�j�@j��D �ٿF�Z�s��@�}�) 4@����!?�3�G�j�@�Y�1�ٿP� b�@������3@���z��!?����QJ�@�Y�1�ٿP� b�@������3@���z��!?����QJ�@�Y�1�ٿP� b�@������3@���z��!?����QJ�@�����ٿ�	v��@��N2��3@��� ��!?� j�R�@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@q���ٿ�2^=#p�@�X�3@�X����!? >�g��@��_�ٿ����D��@�����3@M��x��!?��M����@��_�ٿ����D��@�����3@M��x��!?��M����@��_�ٿ����D��@�����3@M��x��!?��M����@��ieݩٿ2�߷{�@;�K3�3@vp�ҏ!?R�o��*�@��ieݩٿ2�߷{�@;�K3�3@vp�ҏ!?R�o��*�@�qKj��ٿO�GnO)�@���S[�3@�Q�׏!?!��L���@�fDu�ٿ�=��0��@��*] 4@���Ï!?�@Uj�k�@�fDu�ٿ�=��0��@��*] 4@���Ï!?�@Uj�k�@�fDu�ٿ�=��0��@��*] 4@���Ï!?�@Uj�k�@���4��ٿ��SK�@FǷQ��3@5
��!?��ڝ���@���4��ٿ��SK�@FǷQ��3@5
��!?��ڝ���@���4��ٿ��SK�@FǷQ��3@5
��!?��ڝ���@���4��ٿ��SK�@FǷQ��3@5
��!?��ڝ���@]�ϗٿ���,�@��;�)�3@ͣ����!?�B53�\�@]�ϗٿ���,�@��;�)�3@ͣ����!?�B53�\�@]�ϗٿ���,�@��;�)�3@ͣ����!?�B53�\�@�vr@�ٿ��O��f�@��� 4@��ࡏ!?p�.����@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�2�5�ٿ`m}��@�a&�4@�d�(��!?���}QI�@�4��B�ٿ"ʸ��v�@�FV!4@�s�՞�!?��r���@�4��B�ٿ"ʸ��v�@�FV!4@�s�՞�!?��r���@�4��B�ٿ"ʸ��v�@�FV!4@�s�՞�!?��r���@�4��B�ٿ"ʸ��v�@�FV!4@�s�՞�!?��r���@�4��B�ٿ"ʸ��v�@�FV!4@�s�՞�!?��r���@,�y�ٿ9S�Vy�@F�����3@��1��!?����7��@,�y�ٿ9S�Vy�@F�����3@��1��!?����7��@,�y�ٿ9S�Vy�@F�����3@��1��!?����7��@,�y�ٿ9S�Vy�@F�����3@��1��!?����7��@��#�ٿ�������@Og��� 4@��9|o�!?�[����@��#�ٿ�������@Og��� 4@��9|o�!?�[����@��#�ٿ�������@Og��� 4@��9|o�!?�[����@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@镬�E�ٿܪx��@Fj���3@�7Ew(�!?��4�1�@ܷP-?�ٿ��#�q�@�{j�� 4@��o���!?&�=��F�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@;\*.�ٿ��^��@&���� 4@�����!?C�0�@u:�ɥ�ٿ�4����@	��>4@|�C��!?�p�;��@u:�ɥ�ٿ�4����@	��>4@|�C��!?�p�;��@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�����ٿr�^���@��X* 4@29AEm�!?m�/�@�I7P��ٿ�����@�ml[Y4@{���!?|�|$��@�I7P��ٿ�����@�ml[Y4@{���!?|�|$��@�^B�;�ٿ��k���@�FR�� 4@���!?�z�
)�@�^B�;�ٿ��k���@�FR�� 4@���!?�z�
)�@�^B�;�ٿ��k���@�FR�� 4@���!?�z�
)�@�^B�;�ٿ��k���@�FR�� 4@���!?�z�
)�@�r^Ǐٿa�4l���@��0�H 4@f����!?��� M�@�r^Ǐٿa�4l���@��0�H 4@f����!?��� M�@�r^Ǐٿa�4l���@��0�H 4@f����!?��� M�@�r^Ǐٿa�4l���@��0�H 4@f����!?��� M�@^��
#�ٿ�XO8���@>[lQ��3@ �Vu��!?a�$����@�̀��ٿ��uI�`�@����. 4@(�p[�!?�F͐��@�̀��ٿ��uI�`�@����. 4@(�p[�!?�F͐��@�̀��ٿ��uI�`�@����. 4@(�p[�!?�F͐��@�h��3�ٿ�>�l�@76E`;4@ړ�Mc�!?-)����@�dq��ٿ���P��@=9���3@���Qo�!?ԇ��m��@�dq��ٿ���P��@=9���3@���Qo�!?ԇ��m��@�dq��ٿ���P��@=9���3@���Qo�!?ԇ��m��@�dq��ٿ���P��@=9���3@���Qo�!?ԇ��m��@�dq��ٿ���P��@=9���3@���Qo�!?ԇ��m��@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@|�㌣ٿ])�Т��@J�~\��3@�ݶE��!?3�x��G�@���̥ٿcO�D���@B��8��3@e2��͏!?�{��w�@���̥ٿcO�D���@B��8��3@e2��͏!?�{��w�@���̥ٿcO�D���@B��8��3@e2��͏!?�{��w�@���̥ٿcO�D���@B��8��3@e2��͏!?�{��w�@� 4=)�ٿu����^�@�ۇ�4@�5��!?c5�q���@� 4=)�ٿu����^�@�ۇ�4@�5��!?c5�q���@���>��ٿ���j���@oZ:4@��x'ޏ!?z�_�>��@���>��ٿ���j���@oZ:4@��x'ޏ!?z�_�>��@���>��ٿ���j���@oZ:4@��x'ޏ!?z�_�>��@���>��ٿ���j���@oZ:4@��x'ޏ!?z�_�>��@���>��ٿ���j���@oZ:4@��x'ޏ!?z�_�>��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@_guz��ٿ\�\�XE�@}� 4@��1�ߏ!?�F��v��@g�zӣٿ"�k��@��H�� 4@.�$��!?)H��@V#���ٿQpp�k�@�Y5µ 4@��:���!?��]� �@V#���ٿQpp�k�@�Y5µ 4@��:���!?��]� �@V#���ٿQpp�k�@�Y5µ 4@��:���!?��]� �@V#���ٿQpp�k�@�Y5µ 4@��:���!?��]� �@V#���ٿQpp�k�@�Y5µ 4@��:���!?��]� �@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@-N���ٿ�(��:��@��4@��
��!?��J��@	jÕt�ٿf��=���@w�fϰ�3@��*��!?��BVu~�@	jÕt�ٿf��=���@w�fϰ�3@��*��!?��BVu~�@���Nd�ٿmn����@���/��3@�d����!?X>Z����@���Nd�ٿmn����@���/��3@�d����!?X>Z����@���Nd�ٿmn����@���/��3@�d����!?X>Z����@Xs�Xk�ٿw��^Hi�@3�rj��3@��^���!?b��Ʌ�@Xs�Xk�ٿw��^Hi�@3�rj��3@��^���!?b��Ʌ�@Xs�Xk�ٿw��^Hi�@3�rj��3@��^���!?b��Ʌ�@Xs�Xk�ٿw��^Hi�@3�rj��3@��^���!?b��Ʌ�@Xs�Xk�ٿw��^Hi�@3�rj��3@��^���!?b��Ʌ�@)�ٓ��ٿ	О�Y�@��ew)�3@~��׏!?�^H>R��@)�ٓ��ٿ	О�Y�@��ew)�3@~��׏!?�^H>R��@)�ٓ��ٿ	О�Y�@��ew)�3@~��׏!?�^H>R��@)�ٓ��ٿ	О�Y�@��ew)�3@~��׏!?�^H>R��@)�ٓ��ٿ	О�Y�@��ew)�3@~��׏!?�^H>R��@ �"�T�ٿ��So��@х����3@�Q<]
�!?A��@Sa��ϬٿYj��@�(���3@�����!?y����|�@
�s��ٿ���5��@Ҷ"	b�3@�Cͼ�!?_���y�@
�s��ٿ���5��@Ҷ"	b�3@�Cͼ�!?_���y�@
�s��ٿ���5��@Ҷ"	b�3@�Cͼ�!?_���y�@���e��ٿ����@��X��3@#j*���!?l@U���@���e��ٿ����@��X��3@#j*���!?l@U���@���e��ٿ����@��X��3@#j*���!?l@U���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@�ed�ٿ�ߒA*J�@��|�1�3@/3aƏ!?�ص���@Ղa�ٿX�ݛ�@7F!	g�3@>��͏!?�|�O��@Ղa�ٿX�ݛ�@7F!	g�3@>��͏!?�|�O��@Ղa�ٿX�ݛ�@7F!	g�3@>��͏!?�|�O��@A$g�z�ٿtR�����@7aOdc�3@ڨ�ˏ!?�р5�@�A�!�ٿ���jԬ�@�O��e�3@s�T���!?6���B�@�A�!�ٿ���jԬ�@�O��e�3@s�T���!?6���B�@�A�!�ٿ���jԬ�@�O��e�3@s�T���!?6���B�@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@��%�ϡٿ����t�@
�ٟ�3@fT�L�!?��p��@t@>��ٿ_����R�@��l�"�3@�ɻVo�!?�Q �d�@,Gߨٿ?�r�?�@��5�� 4@:����!?�fJC��@,Gߨٿ?�r�?�@��5�� 4@:����!?�fJC��@,Gߨٿ?�r�?�@��5�� 4@:����!?�fJC��@,Gߨٿ?�r�?�@��5�� 4@:����!?�fJC��@,Gߨٿ?�r�?�@��5�� 4@:����!?�fJC��@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�F�ז�ٿ����U��@�Ґ�4@K����!?���@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@�%�A�ٿ���N��@�uz��4@pE�ɬ�!?D�ps��@H�D'��ٿ�T�-��@2Şf��3@�y:���!? j���X�@H�D'��ٿ�T�-��@2Şf��3@�y:���!? j���X�@H�D'��ٿ�T�-��@2Şf��3@�y:���!? j���X�@H�D'��ٿ�T�-��@2Şf��3@�y:���!? j���X�@|��B�ٿ�L�p�w�@�B�E 4@.��Q_�!?���pT��@|��B�ٿ�L�p�w�@�B�E 4@.��Q_�!?���pT��@|��B�ٿ�L�p�w�@�B�E 4@.��Q_�!?���pT��@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@�W-�d�ٿ�b�e���@����� 4@#�^�(�!?� ��}�@e_�dZ�ٿ��J���@���4@�fd�!?��f����@yYm�*�ٿ������@����4@D˳*)�!?E�)G)�@yYm�*�ٿ������@����4@D˳*)�!?E�)G)�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@6p���ٿ�zf�?��@��V�4@�s{�8�!?�Z,��|�@|[����ٿ;%�����@�?��4@��#N|�!?E�nD�@|[����ٿ;%�����@�?��4@��#N|�!?E�nD�@|[����ٿ;%�����@�?��4@��#N|�!?E�nD�@Tr"0?�ٿ�j��b�@2���3@�H8�!?aw����@Tr"0?�ٿ�j��b�@2���3@�H8�!?aw����@������ٿ� �b�@��Ѥ��3@{�w`�!?*}�Ь�@������ٿ� �b�@��Ѥ��3@{�w`�!?*}�Ь�@J-)��ٿS_�+C��@�ۯ80 4@#��*|�!?��ԑ��@J-)��ٿS_�+C��@�ۯ80 4@#��*|�!?��ԑ��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@H�ȱ��ٿ�,rچ��@]B:p4@s&�Ï!?���)��@#�z᭕ٿ���	��@�;_�B4@<=�ŏ!?�m,r��@#�z᭕ٿ���	��@�;_�B4@<=�ŏ!?�m,r��@J�k��ٿ��_�@�B�UY4@�#��!?��1VŪ�@J�k��ٿ��_�@�B�UY4@�#��!?��1VŪ�@��e�àٿ-ӧ�`��@f�f���3@�&ov�!?��q�S8�@��e�àٿ-ӧ�`��@f�f���3@�&ov�!?��q�S8�@��e�àٿ-ӧ�`��@f�f���3@�&ov�!?��q�S8�@����3�ٿ�c~���@-no���3@$�e���!?f'[_ĝ�@����3�ٿ�c~���@-no���3@$�e���!?f'[_ĝ�@����3�ٿ�c~���@-no���3@$�e���!?f'[_ĝ�@����3�ٿ�c~���@-no���3@$�e���!?f'[_ĝ�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@�5��ٿ�&
:�J�@x��L�4@�m���!?����E�@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@//1�^�ٿn,"j�*�@f2T\ 4@�C��!?�=��@@�錩ٿ#� l�E�@/��4@�X_�o�!?V�e�rG�@�f�0:�ٿ�lD<�	�@��
Fe4@�ǅc��!?���$�@�f�0:�ٿ�lD<�	�@��
Fe4@�ǅc��!?���$�@�f�0:�ٿ�lD<�	�@��
Fe4@�ǅc��!?���$�@��p;�ٿ�ܴv���@�sq��3@Մh��!?x;�P\��@��p;�ٿ�ܴv���@�sq��3@Մh��!?x;�P\��@��p;�ٿ�ܴv���@�sq��3@Մh��!?x;�P\��@��p;�ٿ�ܴv���@�sq��3@Մh��!?x;�P\��@]�R��ٿeq\͘�@����3@G$�Gk�!?�b:�|�@]�R��ٿeq\͘�@����3@G$�Gk�!?�b:�|�@]�R��ٿeq\͘�@����3@G$�Gk�!?�b:�|�@]�R��ٿeq\͘�@����3@G$�Gk�!?�b:�|�@]�R��ٿeq\͘�@����3@G$�Gk�!?�b:�|�@?R�`��ٿrgH#��@�+0?�3@�8�1U�!?)w9�?�@?R�`��ٿrgH#��@�+0?�3@�8�1U�!?)w9�?�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@,]3ď�ٿ��4G�@Q��Q��3@�\�za�!?~�k/�J�@Þ���ٿ��2`�;�@�K@/ 4@�☧��!?�aҖn��@Þ���ٿ��2`�;�@�K@/ 4@�☧��!?�aҖn��@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@��]_��ٿ�@!�h�@;U<F��3@��hs��!?Sn�T�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�;�H��ٿKR���@(4@���P��!?D���w4�@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@�B�Jd�ٿ�w����@��]�4@h��s��!?Ew���@&��B��ٿRI��+�@j�S4@��~�!?[��E�@&��B��ٿRI��+�@j�S4@��~�!?[��E�@&��B��ٿRI��+�@j�S4@��~�!?[��E�@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@+�{�ٿ�V��@��8�Q 4@g�,�؏!?��F����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@ղ�A�ٿ���s c�@�9�\4@=�B|�!?�q�����@Ѓ!k��ٿ&>.a=b�@vnt��4@[�s�Տ!?f���(�@Ѓ!k��ٿ&>.a=b�@vnt��4@[�s�Տ!?f���(�@Ѓ!k��ٿ&>.a=b�@vnt��4@[�s�Տ!?f���(�@Q;���ٿ[R�2��@τ��� 4@��
��!?������@Q;���ٿ[R�2��@τ��� 4@��
��!?������@Q;���ٿ[R�2��@τ��� 4@��
��!?������@Q;���ٿ[R�2��@τ��� 4@��
��!?������@Q;���ٿ[R�2��@τ��� 4@��
��!?������@Q;���ٿ[R�2��@τ��� 4@��
��!?������@n7��Z�ٿe2�Y��@g�[ � 4@��W��!?&Z0�i�@2@Th�ٿ:��N��@P�ȯT4@�Ց��!?��Sz�@2@Th�ٿ:��N��@P�ȯT4@�Ց��!?��Sz�@2@Th�ٿ:��N��@P�ȯT4@�Ց��!?��Sz�@2@Th�ٿ:��N��@P�ȯT4@�Ց��!?��Sz�@�tZ�ٿ�x����@��
*� 4@J�+ο�!?�����@�tZ�ٿ�x����@��
*� 4@J�+ο�!?�����@?�k,�ٿ���J	��@�0U%b4@�(��s�!?��v=��@#���[�ٿ�$���@�"	��4@ヺ㾏!?�h�-�@#���[�ٿ�$���@�"	��4@ヺ㾏!?�h�-�@#���[�ٿ�$���@�"	��4@ヺ㾏!?�h�-�@#���[�ٿ�$���@�"	��4@ヺ㾏!?�h�-�@#���[�ٿ�$���@�"	��4@ヺ㾏!?�h�-�@
���)�ٿoK����@�	y�?4@�e��!?�����@
���)�ٿoK����@�	y�?4@�e��!?�����@
���)�ٿoK����@�	y�?4@�e��!?�����@�P&Πٿ=�w���@����~4@+sa�!?���Q�@�P&Πٿ=�w���@����~4@+sa�!?���Q�@�P&Πٿ=�w���@����~4@+sa�!?���Q�@���K��ٿ��=�	�@��go4@�����!?�Q���@���K��ٿ��=�	�@��go4@�����!?�Q���@���K��ٿ��=�	�@��go4@�����!?�Q���@���K��ٿ��=�	�@��go4@�����!?�Q���@���K��ٿ��=�	�@��go4@�����!?�Q���@���K��ٿ��=�	�@��go4@�����!?�Q���@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@ק/���ٿ㞢���@޴�_�3@'��ʃ�!?�x�Dk�@�`n���ٿ�U�HL��@��/2�4@^N��֏!?eL ��@�`n���ٿ�U�HL��@��/2�4@^N��֏!?eL ��@�`n���ٿ�U�HL��@��/2�4@^N��֏!?eL ��@�`n���ٿ�U�HL��@��/2�4@^N��֏!?eL ��@�`n���ٿ�U�HL��@��/2�4@^N��֏!?eL ��@]YC7|�ٿm��r�N�@�r�'� 4@:��d��!?�*l��@ig+�m�ٿ�4��@U$�+�4@����]�!?W>,��@ig+�m�ٿ�4��@U$�+�4@����]�!?W>,��@ig+�m�ٿ�4��@U$�+�4@����]�!?W>,��@ig+�m�ٿ�4��@U$�+�4@����]�!?W>,��@�G-�a�ٿ{@�ͱ��@����3@�Y�W�!?:��p�@�G-�a�ٿ{@�ͱ��@����3@�Y�W�!?:��p�@8�B�4�ٿ��x�g��@�=�ݢ4@c�!?�9�8��@
s/�ٿ�{X�.��@]�ٛp4@���J��!?�yU\�U�@
s/�ٿ�{X�.��@]�ٛp4@���J��!?�yU\�U�@?�_���ٿ+�Ly)�@����4@XH����!?1�$�D�@?�_���ٿ+�Ly)�@����4@XH����!?1�$�D�@�YM���ٿB�^c��@cؽ<4@����!?⚘U.t�@�YM���ٿB�^c��@cؽ<4@����!?⚘U.t�@�YM���ٿB�^c��@cؽ<4@����!?⚘U.t�@�YM���ٿB�^c��@cؽ<4@����!?⚘U.t�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@|:�6�ٿ��+��p�@�أ � 4@q��DǏ!?��:�T�@&��w�ٿ�hRf��@�F��4@�V��Ϗ!?�u����@&��w�ٿ�hRf��@�F��4@�V��Ϗ!?�u����@&��w�ٿ�hRf��@�F��4@�V��Ϗ!?�u����@�K?���ٿ?fD�!��@Nt|=e 4@�#�#r�!?є,�4�@�K?���ٿ?fD�!��@Nt|=e 4@�#�#r�!?є,�4�@�K?���ٿ?fD�!��@Nt|=e 4@�#�#r�!?є,�4�@�K?���ٿ?fD�!��@Nt|=e 4@�#�#r�!?є,�4�@_��e�ٿ���!34�@ϭ>B0 4@�=P��!?�6�- 8�@��{���ٿ�O'��;�@N-l���3@��Q��!?���:�@��{���ٿ�O'��;�@N-l���3@��Q��!?���:�@���2"�ٿ��9`��@dRh��3@�Txe	�!?8��x��@�qI��ٿ��a�?�@~�9�� 4@���BG�!?��+x��@�qI��ٿ��a�?�@~�9�� 4@���BG�!?��+x��@�qI��ٿ��a�?�@~�9�� 4@���BG�!?��+x��@�qI��ٿ��a�?�@~�9�� 4@���BG�!?��+x��@��Mњٿ|�Z����@�v_U.4@�B��J�!?�����@��Mњٿ|�Z����@�v_U.4@�B��J�!?�����@�����ٿ��EX�@��h��3@��m�7�!?��n�4z�@�����ٿ��EX�@��h��3@��m�7�!?��n�4z�@�����ٿ��EX�@��h��3@��m�7�!?��n�4z�@��L>8�ٿw���#��@f�{k�3@8��S�!?>� b���@^8��ٿ��@'F��@�d8���3@�
	\�!?W�م�@^8��ٿ��@'F��@�d8���3@�
	\�!?W�م�@7�*4ǯٿ��?y.�@
@���3@���!?i��\6n�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@�ϻưٿ�b9"��@���D��3@��Ȍ!?4�d� q�@��ؤ��ٿ
'�����@�I��3@Y����!?fp�1��@��ؤ��ٿ
'�����@�I��3@Y����!?fp�1��@��ؤ��ٿ
'�����@�I��3@Y����!?fp�1��@n��H��ٿ#��0E�@�LQ�
�3@A�/�U�!?(Ɩu(��@n��H��ٿ#��0E�@�LQ�
�3@A�/�U�!?(Ɩu(��@����ٿ	�C3�@�,|�4@/�4�Ə!?�s����@����ٿ	�C3�@�,|�4@/�4�Ə!?�s����@����ٿ	�C3�@�,|�4@/�4�Ə!?�s����@@��.^�ٿU�m�z>�@�� 4@ϐ�~��!?)����@@��.^�ٿU�m�z>�@�� 4@ϐ�~��!?)����@@��.^�ٿU�m�z>�@�� 4@ϐ�~��!?)����@�t}� �ٿ�������@�nk� 4@[&�R��!?3]�'��@�t}� �ٿ�������@�nk� 4@[&�R��!?3]�'��@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@ʬl�ٿ�A�og�@f��� 4@a>�Ə!?w�:�L7�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@޶���ٿ�d���@�(�݃�3@d��`ӏ!?.�.b:l�@��s�]�ٿ9c�,��@�-.�� 4@H����!?���tx�@��s�]�ٿ9c�,��@�-.�� 4@H����!?���tx�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@!�ݔٿ����(��@�F�e 4@�K��!?���Pm�@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�0�<�ٿ),�u\��@;���4@9%}�)�!?�'N#���@�}�0��ٿk7Y��@�� �t�3@sh�׏!?I0�\�)�@3'*��ٿȼf�>�@%C3v9 4@�Em���!?����@��@3'*��ٿȼf�>�@%C3v9 4@�Em���!?����@��@3'*��ٿȼf�>�@%C3v9 4@�Em���!?����@��@��:�¡ٿ���k4��@;_G:4@s��؏!?�E�&6��@��:�¡ٿ���k4��@;_G:4@s��؏!?�E�&6��@��:�¡ٿ���k4��@;_G:4@s��؏!?�E�&6��@��:�¡ٿ���k4��@;_G:4@s��؏!?�E�&6��@��:�¡ٿ���k4��@;_G:4@s��؏!?�E�&6��@�@J��ٿ�C:����@>��ȹ 4@hI��ʏ!?�	��_��@�@J��ٿ�C:����@>��ȹ 4@hI��ʏ!?�	��_��@r�Dݑ�ٿ�'�<�2�@qȁ� 4@� �ŏ!?����@r�Dݑ�ٿ�'�<�2�@qȁ� 4@� �ŏ!?����@����t�ٿ{�*��#�@�5�S4@?.��ɏ!?������@����t�ٿ{�*��#�@�5�S4@?.��ɏ!?������@����t�ٿ{�*��#�@�5�S4@?.��ɏ!?������@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@4O=P�ٿ��[5��@��� 4@L�7|�!?���[��@6ToG��ٿ�|��	��@,��� 4@�b"綏!?�sª�Y�@E��""�ٿ�����@����� 4@ߣ��!?|\��F�@E��""�ٿ�����@����� 4@ߣ��!?|\��F�@E��""�ٿ�����@����� 4@ߣ��!?|\��F�@E��""�ٿ�����@����� 4@ߣ��!?|\��F�@E��""�ٿ�����@����� 4@ߣ��!?|\��F�@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@��&��ٿ���xŜ�@l}8��3@m`�R֏!?�c$���@E�����ٿ$b�m�@*�� K�3@����	�!?�.w���@�J��e�ٿ�6J�˲�@U�<���3@�t����!?%��|)��@�q7���ٿ��ɷ��@�{�n4@�t;�~�!?�+�I�~�@�q7���ٿ��ɷ��@�{�n4@�t;�~�!?�+�I�~�@�q7���ٿ��ɷ��@�{�n4@�t;�~�!?�+�I�~�@�q7���ٿ��ɷ��@�{�n4@�t;�~�!?�+�I�~�@�}��ٿ1�'�b��@!���4@ �2#�!?Hj�O�W�@�}��ٿ1�'�b��@!���4@ �2#�!?Hj�O�W�@�}��ٿ1�'�b��@!���4@ �2#�!?Hj�O�W�@�rfy�ٿ�u�␥�@~�&�g4@^5S�ߏ!?��:�3�@��c�ٿj�,;��@��� 4@���S�!?���Ba��@��Pm��ٿg�N��@a |� 4@nni�!?�@��"N�@��Pm��ٿg�N��@a |� 4@nni�!?�@��"N�@��Pm��ٿg�N��@a |� 4@nni�!?�@��"N�@�����ٿ����O�@�<��� 4@E�Ze�!?%�`[���@�����ٿ����O�@�<��� 4@E�Ze�!?%�`[���@�����ٿ����O�@�<��� 4@E�Ze�!?%�`[���@�����ٿ����O�@�<��� 4@E�Ze�!?%�`[���@�|��/�ٿ�3ޟl��@+-�l 4@@��'�!?Ԃ|���@�|��/�ٿ�3ޟl��@+-�l 4@@��'�!?Ԃ|���@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@�Φ�ٿ5n�	���@�,L��4@>����!?�����@����h�ٿ,S�j��@[07�� 4@�|촏!?�)Ee���@����h�ٿ,S�j��@[07�� 4@�|촏!?�)Ee���@����h�ٿ,S�j��@[07�� 4@�|촏!?�)Ee���@����h�ٿ,S�j��@[07�� 4@�|촏!?�)Ee���@����h�ٿ,S�j��@[07�� 4@�|촏!?�)Ee���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@L�h3�ٿg�lB��@̦�� 4@���!��!?g-]���@~���ٿA����@�bH�� 4@�(�׏!?��*��@~���ٿA����@�bH�� 4@�(�׏!?��*��@~���ٿA����@�bH�� 4@�(�׏!?��*��@~���ٿA����@�bH�� 4@�(�׏!?��*��@~���ٿA����@�bH�� 4@�(�׏!?��*��@~���ٿA����@�bH�� 4@�(�׏!?��*��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@"� +)�ٿ\M:v���@%\�x4@�����!?2Y1x}��@ʓ����ٿ�p]���@��A�4@�1 <�!?[�Xfѷ�@��3Φٿ]MI� �@�ˑ�S4@N��[��!?[f��[��@��M� �ٿ���[c��@y��H��3@�	ьϏ!?�9�Ώ�@��M� �ٿ���[c��@y��H��3@�	ьϏ!?�9�Ώ�@��M� �ٿ���[c��@y��H��3@�	ьϏ!?�9�Ώ�@��M� �ٿ���[c��@y��H��3@�	ьϏ!?�9�Ώ�@��M� �ٿ���[c��@y��H��3@�	ьϏ!?�9�Ώ�@d�[�`�ٿ��)�w�@K+�<4@�ܫظ�!?��d��@��WMh�ٿnA�-e��@�6��f 4@l��~�!?>ꊶ1��@u�N��ٿ)A�p��@4���4@f�����!?W^�W��@u�N��ٿ)A�p��@4���4@f�����!?W^�W��@u�N��ٿ)A�p��@4���4@f�����!?W^�W��@u�N��ٿ)A�p��@4���4@f�����!?W^�W��@�h��Q�ٿ� Y����@��`4@�0M���!?}���v��@�h��Q�ٿ� Y����@��`4@�0M���!?}���v��@�h��Q�ٿ� Y����@��`4@�0M���!?}���v��@���F�ٿ=�(A&��@ӷg�d 4@���"��!?'�j]��@���F�ٿ=�(A&��@ӷg�d 4@���"��!?'�j]��@���F�ٿ=�(A&��@ӷg�d 4@���"��!?'�j]��@���F�ٿ=�(A&��@ӷg�d 4@���"��!?'�j]��@���F�ٿ=�(A&��@ӷg�d 4@���"��!?'�j]��@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@֫�%�ٿ���D�h�@a5^P 4@��3숏!?࠰x���@�2�i��ٿ?�rޥn�@��I=\ 4@�ɒ�!?XݚƵ�@�2�i��ٿ?�rޥn�@��I=\ 4@�ɒ�!?XݚƵ�@�2�i��ٿ?�rޥn�@��I=\ 4@�ɒ�!?XݚƵ�@�2�i��ٿ?�rޥn�@��I=\ 4@�ɒ�!?XݚƵ�@�2�i��ٿ?�rޥn�@��I=\ 4@�ɒ�!?XݚƵ�@o��םٿ�Z���e�@�.�� 4@h���!?���zC�@x��b�ٿ����;1�@�_U��3@�}8Ԯ�!?Q\��"�@"u�E�ٿk��'j�@L����4@�[Փ��!?y��_.��@"u�E�ٿk��'j�@L����4@�[Փ��!?y��_.��@`'�i��ٿ�1�4���@�����4@X���l�!?em�Չ[�@`'�i��ٿ�1�4���@�����4@X���l�!?em�Չ[�@#cW���ٿ�ۆz���@���R4@��Wq�!?�l-�&�@��5�ٿ�F�}���@;u���4@�.2���!?�����P�@��5�ٿ�F�}���@;u���4@�.2���!?�����P�@��5�ٿ�F�}���@;u���4@�.2���!?�����P�@��5�ٿ�F�}���@;u���4@�.2���!?�����P�@����ٿ~���@^;��4@x�k_��!?�J��1�@����ٿ~���@^;��4@x�k_��!?�J��1�@����ٿ~���@^;��4@x�k_��!?�J��1�@����ٿ~���@^;��4@x�k_��!?�J��1�@����ٿ~���@^;��4@x�k_��!?�J��1�@�@��ٿbH����@�s�� 4@����!?k��֧�@G.;��ٿ�",��@{�(+f4@E�.{��!?h�f!y��@G.;��ٿ�",��@{�(+f4@E�.{��!?h�f!y��@G.;��ٿ�",��@{�(+f4@E�.{��!?h�f!y��@G.;��ٿ�",��@{�(+f4@E�.{��!?h�f!y��@G.;��ٿ�",��@{�(+f4@E�.{��!?h�f!y��@�y��ٿ^����2�@>`~��4@���.��!?����@Uћ�%�ٿ�}����@4j�V4@��薏!?ۮyN�@Uћ�%�ٿ�}����@4j�V4@��薏!?ۮyN�@Uћ�%�ٿ�}����@4j�V4@��薏!?ۮyN�@Uћ�%�ٿ�}����@4j�V4@��薏!?ۮyN�@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@�?�T��ٿ&��_O(�@���ר4@z��Uď!?r�u���@C_�y�ٿw�
,�i�@���0��3@5��ӏ!?pu�dQ�@C_�y�ٿw�
,�i�@���0��3@5��ӏ!?pu�dQ�@C_�y�ٿw�
,�i�@���0��3@5��ӏ!?pu�dQ�@C_�y�ٿw�
,�i�@���0��3@5��ӏ!?pu�dQ�@C_�y�ٿw�
,�i�@���0��3@5��ӏ!?pu�dQ�@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@���u�ٿ��&}��@{�J��4@�*�Mm�!?*
�u��@�<�牥ٿN'����@̇�H�4@������!?r��4��@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@0���ٿ&��lX��@�億 4@{cù�!?� r���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�ʉbp�ٿiY���@��t	��3@f�Х�!?k���@�#ئ��ٿ�5�L�p�@Qy6k 4@�a��t�!?Bp��8�@�? �o�ٿ��d>~*�@n��ז�3@ _���!?��}b �@����ٿ��G���@ɬ�� 4@�����!?��o@�@0�6{"�ٿ�˼����@>C	5��3@r�}齏!?����r�@Ȼ��l�ٿ)��	Wz�@�G'���3@A�ٿ�!??��t�@Ȼ��l�ٿ)��	Wz�@�G'���3@A�ٿ�!??��t�@����ٿ7�	���@��'M��3@��K���!?*���@����ٿ7�	���@��'M��3@��K���!?*���@����ٿ7�	���@��'M��3@��K���!?*���@����ٿ7�	���@��'M��3@��K���!?*���@����ٿ7�	���@��'M��3@��K���!?*���@�H�~�ٿɆg�p��@���� 4@������!?meDe���@�H�~�ٿɆg�p��@���� 4@������!?meDe���@�H�~�ٿɆg�p��@���� 4@������!?meDe���@�H�~�ٿɆg�p��@���� 4@������!?meDe���@� �8�ٿ�P�W��@��;�4@>t��!?4���+�@� �8�ٿ�P�W��@��;�4@>t��!?4���+�@� �8�ٿ�P�W��@��;�4@>t��!?4���+�@�7*�ٿ#��.���@���f��3@P�>Ƞ�!?%�]�L�@�7*�ٿ#��.���@���f��3@P�>Ƞ�!?%�]�L�@�7*�ٿ#��.���@���f��3@P�>Ƞ�!?%�]�L�@�7*�ٿ#��.���@���f��3@P�>Ƞ�!?%�]�L�@�Vf7��ٿ,��!��@D� � 4@df-%��!?y�^�3��@V��=b�ٿlfE��v�@R#��  4@��˱�!?F
�x��@V��=b�ٿlfE��v�@R#��  4@��˱�!?F
�x��@��\B��ٿ��E>�@mR,���3@B�]�!?�9uS��@��ZȩٿlI���@h�6z� 4@ؘpEK�!?���:ъ�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�qL���ٿ�sR���@\> �� 4@8�p«�!?���	�@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@�b� �ٿ/ 9���@8.�"4@��/��!?Ƚ�4��@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@׬)]�ٿ�#�c��@�>b	�4@y@ܭ�!?p��"�8�@�'GĨٿY� �\�@^��S^ 4@�F/D��!?���-�@�'GĨٿY� �\�@^��S^ 4@�F/D��!?���-�@O����ٿ҇w�L"�@HN-� 4@|�귏!?Xcbє�@O����ٿ҇w�L"�@HN-� 4@|�귏!?Xcbє�@?�����ٿF�y�X��@f�#M 4@-\.c��!?rakl�@?�����ٿF�y�X��@f�#M 4@-\.c��!?rakl�@�M�\-�ٿ��V>��@y�h%U 4@��5X�!?��*ͩ�@.7a�ٿ� �	���@/��,q4@n���N�!?��@���@.7a�ٿ� �	���@/��,q4@n���N�!?��@���@.7a�ٿ� �	���@/��,q4@n���N�!?��@���@�1"�}�ٿ��~o�@��7�R4@����L�!?N��<��@^A���ٿ��aѱ��@ұ�Mf4@�c�'�!?��<[�@�ԉQ$�ٿ]���V�@X��� 4@��:�O�!? �uI���@�ԉQ$�ٿ]���V�@X��� 4@��:�O�!? �uI���@&ت�\�ٿv?�A`�@�Wb�|4@?j��a�!?�QJ�n�@&ت�\�ٿv?�A`�@�Wb�|4@?j��a�!?�QJ�n�@&ت�\�ٿv?�A`�@�Wb�|4@?j��a�!?�QJ�n�@���߯ٿ�w�ɹ�@�k�1�4@��l^�!?�.2���@���߯ٿ�w�ɹ�@�k�1�4@��l^�!?�.2���@���߯ٿ�w�ɹ�@�k�1�4@��l^�!?�.2���@�X\ٮٿ�k\��\�@�@Q��4@S�X�Z�!?��l;�@�X\ٮٿ�k\��\�@�@Q��4@S�X�Z�!?��l;�@�X\ٮٿ�k\��\�@�@Q��4@S�X�Z�!?��l;�@�X\ٮٿ�k\��\�@�@Q��4@S�X�Z�!?��l;�@�X\ٮٿ�k\��\�@�@Q��4@S�X�Z�!?��l;�@5���;�ٿYQ&gKq�@W6���4@AF����!?�x��^��@5���;�ٿYQ&gKq�@W6���4@AF����!?�x��^��@5���;�ٿYQ&gKq�@W6���4@AF����!?�x��^��@�\�&�ٿ��:���@�6���4@U�!d�!?i�W�@�\�&�ٿ��:���@�6���4@U�!d�!?i�W�@a�G �ٿfؕ�c�@n�E�4@4���`�!?v� �A�@a�G �ٿfؕ�c�@n�E�4@4���`�!?v� �A�@:sX&�ٿ]%��QY�@�0� 4@�J�gx�!?������@:sX&�ٿ]%��QY�@�0� 4@�J�gx�!?������@:sX&�ٿ]%��QY�@�0� 4@�J�gx�!?������@���
�ٿ�����}�@#|�d�4@��dT��!?�@&�?�@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@�I����ٿ�8����@7�� � 4@���!?G���g��@s����ٿ��I�z��@�b�W 4@���r�!?7?m<�@s����ٿ��I�z��@�b�W 4@���r�!?7?m<�@s����ٿ��I�z��@�b�W 4@���r�!?7?m<�@s����ٿ��I�z��@�b�W 4@���r�!?7?m<�@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@��x@��ٿ�"1��@�쿧 4@Z�j�L�!?o0d`��@�؈н�ٿ��|5�U�@�#���4@h��6g�!?=!��
�@�؈н�ٿ��|5�U�@�#���4@h��6g�!?=!��
�@�؈н�ٿ��|5�U�@�#���4@h��6g�!?=!��
�@�؈н�ٿ��|5�U�@�#���4@h��6g�!?=!��
�@p�y7�ٿ�x�d���@L�0#4@D�20O�!?�m���@��u>*�ٿ�.�0��@K23��3@������!?����C�@��u>*�ٿ�.�0��@K23��3@������!?����C�@��).�ٿR���{0�@�.�W� 4@d/o)u�!?��C{��@��).�ٿR���{0�@�.�W� 4@d/o)u�!?��C{��@f�Vj��ٿ��9F;<�@i���4@ͷ/���!?��~��@���\��ٿi�UU�@o��q�4@L+�6��!?�{�nL��@���\��ٿi�UU�@o��q�4@L+�6��!?�{�nL��@���\��ٿi�UU�@o��q�4@L+�6��!?�{�nL��@���\��ٿi�UU�@o��q�4@L+�6��!?�{�nL��@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@o�h�u�ٿI���(�@�,k6� 4@Y�v���!?�S�?���@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@z�P6��ٿ49����@��)f� 4@� ���!?xu2]l�@Q'g~��ٿ0W� i`�@<H�;��3@{0�̏!?����@��n���ٿ��s|��@�1uv6�3@Z��Տ!?�ǃ,ē�@��n���ٿ��s|��@�1uv6�3@Z��Տ!?�ǃ,ē�@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@�`z8��ٿ����qS�@�0��3@������!?6�����@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@"i)��ٿ�5����@ꣷ>: 4@J��!?�Zka$�@���T�ٿn�Gu�@�$���3@ez�7�!?t�>#��@���T�ٿn�Gu�@�$���3@ez�7�!?t�>#��@+��w)�ٿ�K�Uy��@Fw�!M�3@kP�Vۏ!?��<6j�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@�#"�ԫٿ3:)�Ɗ�@�O����3@��� 	�!?Ϸ��>�@~ �E�ٿ᠑D���@��~=�3@p���!?b�m���@~ �E�ٿ᠑D���@��~=�3@p���!?b�m���@~ �E�ٿ᠑D���@��~=�3@p���!?b�m���@~ �E�ٿ᠑D���@��~=�3@p���!?b�m���@~ �E�ٿ᠑D���@��~=�3@p���!?b�m���@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@�ѫᑤٿC'�5� �@�^��3@��n ԏ!?���ۑ[�@m�:d�ٿ���`&*�@H#>�3@��@�!?a���)�@��Ni��ٿ~�h����@* ���3@V��7��!?d�sj%�@��Ni��ٿ~�h����@* ���3@V��7��!?d�sj%�@��Ni��ٿ~�h����@* ���3@V��7��!?d�sj%�@��Ni��ٿ~�h����@* ���3@V��7��!?d�sj%�@��Ni��ٿ~�h����@* ���3@V��7��!?d�sj%�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@�uȢ��ٿeZ�I��@�E6�^�3@��l���!?�XY�W�@c���D�ٿ	h��h��@(��9�3@�S�}��!?oD�|��@c���D�ٿ	h��h��@(��9�3@�S�}��!?oD�|��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@���F�ٿ O/�ٚ�@L�� 4@���ף�!?_���4��@[͏!�ٿ�?�"P�@S-�T� 4@8 ���!?�������@�y:�s�ٿnv��M�@n>9O 4@`���!?¹ԑ= �@�y:�s�ٿnv��M�@n>9O 4@`���!?¹ԑ= �@�y:�s�ٿnv��M�@n>9O 4@`���!?¹ԑ= �@�y:�s�ٿnv��M�@n>9O 4@`���!?¹ԑ= �@�y:�s�ٿnv��M�@n>9O 4@`���!?¹ԑ= �@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@k?o�
�ٿm1�6V�@~��� 4@�O�Z��!?��#��E�@�����ٿ��ȟ� �@�l4@	�ER��!?�[/�<�@�����ٿ��ȟ� �@�l4@	�ER��!?�[/�<�@��I���ٿ�s�	���@k���d4@��q�u�!?���k���@y�r3�ٿ���)��@k&�05 4@>Ǫ+��!?�?���h�@y�r3�ٿ���)��@k&�05 4@>Ǫ+��!?�?���h�@y�r3�ٿ���)��@k&�05 4@>Ǫ+��!?�?���h�@����T�ٿ�Gj��O�@�$۱ 4@���tz�!?↼+�@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@:�0n�ٿ�Ǥ_u�@8����3@�!1 r�!?�����@'%��ٿt�A�s�@�X��q�3@�mF^~�!?��S�@ȕ睩ٿ	=��sJ�@�
�N#�3@���HY�!?k#���@�'8��ٿTV
��@���J 4@G>b��!?�[u��|�@�'8��ٿTV
��@���J 4@G>b��!?�[u��|�@��ޜٿ���V(k�@�얟4@��"���!?={�<�@����I�ٿ񘘰Ɵ�@�ܲ�4@��i�d�!?�p��t`�@�4�fY�ٿS�5Z���@]t��/4@c-�]̏!?�ZӠ��@�z;i7�ٿ���P��@�5��4@��u�׏!?$��'�@�P���ٿ{���Q�@W�[�4@�ݡt�!?),���)�@�P���ٿ{���Q�@W�[�4@�ݡt�!?),���)�@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@)����ٿ���5�q�@LG���3@+�z=��!?"�F���@d���"�ٿ[��h��@[�1n 4@�	c�!?�"-��@d���"�ٿ[��h��@[�1n 4@�	c�!?�"-��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@����ʝٿ��a���@L�� 4@��tv�!?�ʜ!x��@�!R��ٿ/e�ܐv�@���k4@��jR�!?���D��@vM���ٿ]:���@����4@gp�0�!?��l�p�@y�=0�ٿt]����@�2�}E 4@y�8;�!?���W�4�@y�=0�ٿt]����@�2�}E 4@y�8;�!?���W�4�@y�=0�ٿt]����@�2�}E 4@y�8;�!?���W�4�@y�=0�ٿt]����@�2�}E 4@y�8;�!?���W�4�@yI(�ٿ�Y��:��@6��1J�3@PC4峏!?�������@yI(�ٿ�Y��:��@6��1J�3@PC4峏!?�������@yI(�ٿ�Y��:��@6��1J�3@PC4峏!?�������@yI(�ٿ�Y��:��@6��1J�3@PC4峏!?�������@yI(�ٿ�Y��:��@6��1J�3@PC4峏!?�������@s���Z�ٿh�a��G�@�t��3@�h�q�!?������@s���Z�ٿh�a��G�@�t��3@�h�q�!?������@s���Z�ٿh�a��G�@�t��3@�h�q�!?������@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@ނGQ�ٿ�r���g�@�LD� 4@���w�!?��Hb�@�n�z:�ٿMB�i���@D�Ґ�4@�(ab��!?���`�t�@�n�z:�ٿMB�i���@D�Ґ�4@�(ab��!?���`�t�@�n�z:�ٿMB�i���@D�Ґ�4@�(ab��!?���`�t�@�n�z:�ٿMB�i���@D�Ґ�4@�(ab��!?���`�t�@�����ٿ���i׺�@���4�4@V���}�!?3cb���@�����ٿ���i׺�@���4�4@V���}�!?3cb���@�����ٿ���i׺�@���4�4@V���}�!?3cb���@�73W�ٿ��l�ݮ�@u��6�4@5�[�!?��β��@�73W�ٿ��l�ݮ�@u��6�4@5�[�!?��β��@�73W�ٿ��l�ݮ�@u��6�4@5�[�!?��β��@�73W�ٿ��l�ݮ�@u��6�4@5�[�!?��β��@6�ާٿ���`�`�@UNP+� 4@eXY*��!?E�G�d�@>��ٿ���k��@�� 4@����!?�qU�Z�@#�/�'�ٿ�W<�1��@_���!4@��v���!?��nd�<�@#�/�'�ٿ�W<�1��@_���!4@��v���!?��nd�<�@#�/�'�ٿ�W<�1��@_���!4@��v���!?��nd�<�@#�/�'�ٿ�W<�1��@_���!4@��v���!?��nd�<�@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@͗�Bɚٿ�J����@�%-t4@gϳڏ!?=�0��@M�n���ٿuߺ�K�@�?�|{4@�E�x��!?�=Y���@M�n���ٿuߺ�K�@�?�|{4@�E�x��!?�=Y���@(%���ٿO<'@��@V�\�34@A$c�!?���p���@(%���ٿO<'@��@V�\�34@A$c�!?���p���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@�!��ٿpA�䩽�@���\�4@$���`�!?1���@h�ʙٿ���G���@�s6(J 4@�&���!?�W�.���@h�ʙٿ���G���@�s6(J 4@�&���!?�W�.���@h�ʙٿ���G���@�s6(J 4@�&���!?�W�.���@h�ʙٿ���G���@�s6(J 4@�&���!?�W�.���@�5���ٿ|p3J���@ط�kU 4@˼pm��!?f���$M�@�EtfY�ٿr"�'�k�@Sw��b 4@�=�W�!?�CO���@�EtfY�ٿr"�'�k�@Sw��b 4@�=�W�!?�CO���@�EtfY�ٿr"�'�k�@Sw��b 4@�=�W�!?�CO���@= ����ٿ�����@ɔTC�4@�Ż�
�!?g��~:�@= ����ٿ�����@ɔTC�4@�Ż�
�!?g��~:�@= ����ٿ�����@ɔTC�4@�Ż�
�!?g��~:�@= ����ٿ�����@ɔTC�4@�Ż�
�!?g��~:�@����x�ٿ������@f�m��3@f���ӏ!?�7}��@����x�ٿ������@f�m��3@f���ӏ!?�7}��@����x�ٿ������@f�m��3@f���ӏ!?�7}��@����x�ٿ������@f�m��3@f���ӏ!?�7}��@����x�ٿ������@f�m��3@f���ӏ!?�7}��@2��C��ٿ+�n��@:'ڥ�4@�{���!?����5l�@4�M+h�ٿ櫧��y�@臌��4@^��k�!?dUA��@4�M+h�ٿ櫧��y�@臌��4@^��k�!?dUA��@��9�M�ٿ��Yב^�@���i4@|��HK�!?�l�<�@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@OCxʥٿևZ�U�@�M��) 4@k���@�!?)�R��@^��N�ٿ$q� ��@�� �_ 4@ֈ0H��!? 娂�)�@^��N�ٿ$q� ��@�� �_ 4@ֈ0H��!? 娂�)�@^��N�ٿ$q� ��@�� �_ 4@ֈ0H��!? 娂�)�@����&�ٿۑl%�N�@2��q 4@i/�Ϗ!?�P	̦��@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@7�)@�ٿ`�����@e�Aq�4@�i����!?�"{p�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���R�ٿ���(��@l񈧣4@�ß��!?�@��'�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@���Iw�ٿ�-md��@c��>7 4@8���!?IW4dd�@��s�ٿ�&+e��@�L�.��3@���M��!?.���@��s�ٿ�&+e��@�L�.��3@���M��!?.���@��s�ٿ�&+e��@�L�.��3@���M��!?.���@��s�ٿ�&+e��@�L�.��3@���M��!?.���@��s�ٿ�&+e��@�L�.��3@���M��!?.���@�� �ٿ&k�`	�@$�@Y�4@�j&��!?�5���~�@�<�I��ٿ�*����@��e��3@���u~�!?ŵ���<�@w#�9��ٿ��c�&�@��(���3@������!?%����@��8�ٿ���iO*�@YZM;�3@���XN�!?���6d��@��8�ٿ���iO*�@YZM;�3@���XN�!?���6d��@��8�ٿ���iO*�@YZM;�3@���XN�!?���6d��@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@�#I��ٿ�76��@�j�j��3@�\�(n�!?C�f�L�@4j'�ٿ	`E��@⥿��3@��c��!?3��Z!��@4j'�ٿ	`E��@⥿��3@��c��!?3��Z!��@4j'�ٿ	`E��@⥿��3@��c��!?3��Z!��@7��[�ٿ&�2C�@��,��3@\{��Џ!?#���v�@0n��ٿ�xB��@a�K0 4@B���!?c)\���@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@�28z��ٿP�3��f�@1�_�J 4@!
e� �!?�ثr��@*^��q�ٿ��A7�@��G�4@��
8{�!?�R���/�@*^��q�ٿ��A7�@��G�4@��
8{�!?�R���/�@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@P�Ґ�ٿ���]��@��Ԛ4@Zsfj�!?�s&D��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@�㛔ٿ�cP�o��@O�f�� 4@A�h��!?��4(��@��afJ�ٿ(�RJKv�@��#6s 4@,\�t��!?��"����@��_V��ٿzoѾKZ�@:~ݿ`�3@���4�!?�ig{*��@�)O�k�ٿY������@��!��3@�����!?����M��@i����ٿ��%	��@��f]��3@�KW嫏!?������@i����ٿ��%	��@��f]��3@�KW嫏!?������@i����ٿ��%	��@��f]��3@�KW嫏!?������@i����ٿ��%	��@��f]��3@�KW嫏!?������@i����ٿ��%	��@��f]��3@�KW嫏!?������@i����ٿ��%	��@��f]��3@�KW嫏!?������@������ٿ��l���@����4@[�����!?�/�7�@������ٿ��l���@����4@[�����!?�/�7�@������ٿ��l���@����4@[�����!?�/�7�@������ٿ��l���@����4@[�����!?�/�7�@������ٿ��l���@����4@[�����!?�/�7�@��7�ٿ�W����@@/ܡ4@D����!?�"�H��@��7�ٿ�W����@@/ܡ4@D����!?�"�H��@��7�ٿ�W����@@/ܡ4@D����!?�"�H��@��6L�ٿ�T n*��@�q~�N4@�+��!?�м����@��6L�ٿ�T n*��@�q~�N4@�+��!?�м����@��wg�ٿ��ـLF�@F���4�3@�����!?��K��@C��^��ٿi��a���@�g٬�3@�Rj줏!?_LH�ʊ�@C��^��ٿi��a���@�g٬�3@�Rj줏!?_LH�ʊ�@C��^��ٿi��a���@�g٬�3@�Rj줏!?_LH�ʊ�@�f?C�ٿ��l$��@��e��4@1�1��!?�R�����@�f?C�ٿ��l$��@��e��4@1�1��!?�R�����@�.�{0�ٿz�p�uN�@?J���3@�n_S͏!?`�'��@�.�{0�ٿz�p�uN�@?J���3@�n_S͏!?`�'��@�.�{0�ٿz�p�uN�@?J���3@�n_S͏!?`�'��@�&ȡ �ٿ�CL�/�@A�����3@P�M3̏!?9Y�G��@�&ȡ �ٿ�CL�/�@A�����3@P�M3̏!?9Y�G��@�&ȡ �ٿ�CL�/�@A�����3@P�M3̏!?9Y�G��@�&ȡ �ٿ�CL�/�@A�����3@P�M3̏!?9Y�G��@�&ȡ �ٿ�CL�/�@A�����3@P�M3̏!?9Y�G��@_@f��ٿN�0�c��@e�����3@$�Dя!?/L���@�OǍc�ٿ-�]pG�@�� ��3@d��Ǐ!?�(S��@�OǍc�ٿ-�]pG�@�� ��3@d��Ǐ!?�(S��@�OǍc�ٿ-�]pG�@�� ��3@d��Ǐ!?�(S��@�OǍc�ٿ-�]pG�@�� ��3@d��Ǐ!?�(S��@�OǍc�ٿ-�]pG�@�� ��3@d��Ǐ!?�(S��@�kW �ٿ���w���@4�� 4@I��*h�!?7����@�kW �ٿ���w���@4�� 4@I��*h�!?7����@nF(s�ٿ�=ܼ*�@�,��_4@&f8��!?�2Fu�@nF(s�ٿ�=ܼ*�@�,��_4@&f8��!?�2Fu�@�jRg��ٿ�ދ0x|�@���4@<�W��!?�������@�jRg��ٿ�ދ0x|�@���4@<�W��!?�������@�jRg��ٿ�ދ0x|�@���4@<�W��!?�������@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@�ߞ��ٿ��2���@,�TBG 4@̳�V�!?d�c,])�@��5hy�ٿ���]d�@�N9��3@+�U�!?�cFw{j�@��5hy�ٿ���]d�@�N9��3@+�U�!?�cFw{j�@��5hy�ٿ���]d�@�N9��3@+�U�!?�cFw{j�@��5hy�ٿ���]d�@�N9��3@+�U�!?�cFw{j�@7�AD��ٿF�x�@���r`�3@��W�6�!?�o����@7�AD��ٿF�x�@���r`�3@��W�6�!?�o����@W�:�ٿh�t=�@�Ȓ���3@�9����!?��/k�k�@W�:�ٿh�t=�@�Ȓ���3@�9����!?��/k�k�@W�:�ٿh�t=�@�Ȓ���3@�9����!?��/k�k�@W�:�ٿh�t=�@�Ȓ���3@�9����!?��/k�k�@W�:�ٿh�t=�@�Ȓ���3@�9����!?��/k�k�@Q�7�x�ٿ��3{�Y�@K��` 4@�ᖨq�!?S$�D���@�zC��ٿ�ۻb��@Gݭk��3@ΣX�:�!?�ݧK��@�zC��ٿ�ۻb��@Gݭk��3@ΣX�:�!?�ݧK��@�zC��ٿ�ۻb��@Gݭk��3@ΣX�:�!?�ݧK��@�zC��ٿ�ۻb��@Gݭk��3@ΣX�:�!?�ݧK��@�zC��ٿ�ۻb��@Gݭk��3@ΣX�:�!?�ݧK��@���̻�ٿ�,�Y��@�)4@������!?�m*aF��@���̻�ٿ�,�Y��@�)4@������!?�m*aF��@���̻�ٿ�,�Y��@�)4@������!?�m*aF��@xV#���ٿokO;��@��s�o4@t�$�B�!?��X���@xV#���ٿokO;��@��s�o4@t�$�B�!?��X���@xV#���ٿokO;��@��s�o4@t�$�B�!?��X���@����Z�ٿ�(����@�D�?4@d2�VR�!?ﴚ�i��@����ٿLɯ�ev�@�հ!4@B��B�!?�x0	��@����ٿLɯ�ev�@�հ!4@B��B�!?�x0	��@����ٿLɯ�ev�@�հ!4@B��B�!?�x0	��@����ٿLɯ�ev�@�հ!4@B��B�!?�x0	��@��EwݥٿL�����@�B�ߨ4@�����!?���0�@7ı�ٿF��~<��@���3@� �ޏ!?MC���@�P�=�ٿ2wA���@���^4@^�ڤ�!?@z�b�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�Y�z�ٿ)l��=�@d� 4@�Y�dˏ!?��Fd4J�@�@M\��ٿ$z����@q��� 4@�ש�W�!?\�|H�@�@M\��ٿ$z����@q��� 4@�ש�W�!?\�|H�@�@M\��ٿ$z����@q��� 4@�ש�W�!?\�|H�@�@M\��ٿ$z����@q��� 4@�ש�W�!?\�|H�@%Hca��ٿ.�j�M�@�U�Q 4@x~��!?w�=�m��@����ɟٿYCn���@z>~���3@.��1�!?VzOߋ��@����ɟٿYCn���@z>~���3@.��1�!?VzOߋ��@����ɟٿYCn���@z>~���3@.��1�!?VzOߋ��@����ɟٿYCn���@z>~���3@.��1�!?VzOߋ��@����ʧٿk5x�N�@	Ý�4@E��R �!?W���@l��8��ٿ���Y��@J�w��3@TLحd�!?�#-j>��@l��8��ٿ���Y��@J�w��3@TLحd�!?�#-j>��@l��8��ٿ���Y��@J�w��3@TLحd�!?�#-j>��@#�4[�ٿ�����@��KF��3@�e!?��&��@#�4[�ٿ�����@��KF��3@�e!?��&��@#�4[�ٿ�����@��KF��3@�e!?��&��@#�4[�ٿ�����@��KF��3@�e!?��&��@#�4[�ٿ�����@��KF��3@�e!?��&��@#�4[�ٿ�����@��KF��3@�e!?��&��@��C4v�ٿ(�+��n�@H�>� 4@�Xr��!?u�Z?R�@��C4v�ٿ(�+��n�@H�>� 4@�Xr��!?u�Z?R�@��C4v�ٿ(�+��n�@H�>� 4@�Xr��!?u�Z?R�@��C4v�ٿ(�+��n�@H�>� 4@�Xr��!?u�Z?R�@��C4v�ٿ(�+��n�@H�>� 4@�Xr��!?u�Z?R�@[i�1�ٿ�z��@@.�w� 4@�n3ꄏ!?ףQ?%K�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@*�n=Φٿ�Y��V��@V�چ� 4@�]�2��!?�<�7*�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@���G4�ٿ�Ð�@�����3@�B�~�!?���zP�@A;�ըٿ8��u��@\g/)��3@�D͜�!?��(�a_�@A;�ըٿ8��u��@\g/)��3@�D͜�!?��(�a_�@A;�ըٿ8��u��@\g/)��3@�D͜�!?��(�a_�@A;�ըٿ8��u��@\g/)��3@�D͜�!?��(�a_�@A;�ըٿ8��u��@\g/)��3@�D͜�!?��(�a_�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@_�!���ٿV,�s��@��.�D4@N��F��!?�C�P�@�z��ٿF2:ux�@�߷74@֏����!?m��;�X�@���_�ٿp�-y�?�@���+�4@SX_�!?�a���@��b�ٿk��x�H�@TT���4@6*9�z�!?U�u��@y��Iܧٿ���tR�@\\��3@�ĉ�!?yw@����@y��Iܧٿ���tR�@\\��3@�ĉ�!?yw@����@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�l���ٿY�H@�@��W�� 4@�'���!?�G3Q�@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@�J��ٿ����F�@���� 4@\f�`z�!?;a���@4�=q��ٿ�!K�[��@�3�c4@�P\�~�!?Iܝ��&�@~uD��ٿf����@8��8V4@�"�,��!?��zAG�@�i�b�ٿ�'Q�R��@�ۢ4@;V�#r�!?@obj�c�@�i�b�ٿ�'Q�R��@�ۢ4@;V�#r�!?@obj�c�@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@���4��ٿ��bj)�@䖩��4@
�ȏ!?5[[MR��@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@�DTȣٿ3�O=j��@	c���4@���R��!?b_�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@+����ٿ�D�����@P@�� 4@'�Gz{�!?g��t�@�i�Ҵ�ٿ��V
�@�H���3@��k��!?�1����@�i�Ҵ�ٿ��V
�@�H���3@��k��!?�1����@�i�Ҵ�ٿ��V
�@�H���3@��k��!?�1����@�i�Ҵ�ٿ��V
�@�H���3@��k��!?�1����@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@,�?�ٿ�(DM�5�@2���K�3@�[��Ώ!?d�#�%z�@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@�wW��ٿ���#
��@���3@�����!?P�[����@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@$�:�èٿ����ϴ�@�ˢ�4@}����!?���T���@��ٿ��t�Ih�@�Ш�J 4@�Y�.ޏ!?�,����@��ٿ��t�Ih�@�Ш�J 4@�Y�.ޏ!?�,����@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@��t�{�ٿ�M�V�@��p>� 4@���ʗ�!?�R�4�@m�6�g�ٿ� /!/9�@��e2�4@��,V�!?WV���P�@��¡ٿ��a6���@���4@D[p9H�!?�(���d�@3~
�ٿq��h��@J_4@&��W>�!?1���5��@0z5�$�ٿ�Fkܡ��@2���4@�5-�!?��\��@0z5�$�ٿ�Fkܡ��@2���4@�5-�!?��\��@��ى��ٿ+l:���@Բ���4@��a�v�!?������@��ى��ٿ+l:���@Բ���4@��a�v�!?������@�Y=뚫ٿG�k-��@��RRI4@d	 ���!?�7T�O�@R��ڂ�ٿ�N����@�v��4@��5̏!? ����k�@�\G��ٿ�X�s�@�@���b��3@as��ُ!?�}�2��@�ܼ��ٿ%���C�@p-S�4@��M��!?y~��p�@Gd1B�ٿ��Mތ��@Tnf݇4@��Q^�!?��	T�s�@Gd1B�ٿ��Mތ��@Tnf݇4@��Q^�!?��	T�s�@Gd1B�ٿ��Mތ��@Tnf݇4@��Q^�!?��	T�s�@Gd1B�ٿ��Mތ��@Tnf݇4@��Q^�!?��	T�s�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@D��7�ٿ�� (�%�@�l� 4@������!?�����o�@�oj�˟ٿ��}$��@�c��3@c��nӏ!?�J��0�@�oj�˟ٿ��}$��@�c��3@c��nӏ!?�J��0�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@�_���ٿ�Kxh���@3��6��3@R��(��!?%��<�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@k�Ԭٿ�B��j�@��9��3@��͏!?����T�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@ș�	D�ٿ���e���@E."� 4@HmN�!?��C�Q<�@��j��ٿz�P����@ l� 4@,��z�!?�������@��j��ٿz�P����@ l� 4@,��z�!?�������@��j��ٿz�P����@ l� 4@,��z�!?�������@K��5{�ٿ��7���@gͦ�4@�[ڡ�!?�������@	=���ٿ���S���@�8��4@�f%�r�!?p��C��@;����ٿ!I���2�@LD�bm4@faL~�!?:����@;����ٿ!I���2�@LD�bm4@faL~�!?:����@2t�鯰ٿe��;�e�@�<4@7��⻏!?�:33&��@2t�鯰ٿe��;�e�@�<4@7��⻏!?�:33&��@2t�鯰ٿe��;�e�@�<4@7��⻏!?�:33&��@�.��ٿ����R��@j{��4@�k���!?��V�Z��@�.��ٿ����R��@j{��4@�k���!?��V�Z��@�.��ٿ����R��@j{��4@�k���!?��V�Z��@�]��ٿ�$�,���@烱g4@:a�<Ə!?�������@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@s��6�ٿi N-���@��� 4@v����!?�&S%��@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@����[�ٿ4~D���@���%�3@"5�E��!?�A�r�[�@O��t�ٿ���(��@�,����3@$bE��!?�I3�@��r�ٿ���>�z�@�J��^ 4@i��!?�P�v���@��r�ٿ���>�z�@�J��^ 4@i��!?�P�v���@��r�ٿ���>�z�@�J��^ 4@i��!?�P�v���@zC�B��ٿK["Ii�@�7�q 4@,�' ��!?��ˍ��@zC�B��ٿK["Ii�@�7�q 4@,�' ��!?��ˍ��@\9q�ٿ"2'ٵ��@(r0�4@����W�!?���{���@\9q�ٿ"2'ٵ��@(r0�4@����W�!?���{���@\9q�ٿ"2'ٵ��@(r0�4@����W�!?���{���@\9q�ٿ"2'ٵ��@(r0�4@����W�!?���{���@��m�`�ٿ0��a���@����*4@���X�!?R�5���@��m�`�ٿ0��a���@����*4@���X�!?R�5���@��m�`�ٿ0��a���@����*4@���X�!?R�5���@��m�`�ٿ0��a���@����*4@���X�!?R�5���@��m�`�ٿ0��a���@����*4@���X�!?R�5���@�<�֞ٿ|��O�@��'��4@�(�N�!?;\9����@F�ޗ�ٿ\6D�W-�@��p��4@m_���!?v|�:SE�@F�ޗ�ٿ\6D�W-�@��p��4@m_���!?v|�:SE�@F�ޗ�ٿ\6D�W-�@��p��4@m_���!?v|�:SE�@F�ޗ�ٿ\6D�W-�@��p��4@m_���!?v|�:SE�@���o\�ٿ8K�)���@Z�����3@\8
/�!?	S����@���o\�ٿ8K�)���@Z�����3@\8
/�!?	S����@���o\�ٿ8K�)���@Z�����3@\8
/�!?	S����@�654�ٿË?�H��@A)"���3@�ue ׏!?C�����@�654�ٿË?�H��@A)"���3@�ue ׏!?C�����@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@+�bb��ٿ�^ϳ��@I[�54@�b#⚏!?�I��Zm�@�AI�˜ٿ��
�ћ�@��	4@5��rd�!?�dX?(��@]��텚ٿ��<%��@q�u�4@\m��?�!?_����*�@]��텚ٿ��<%��@q�u�4@\m��?�!?_����*�@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�W����ٿ�执*��@��� �4@d��J3�!?Xg%t8��@�Ûتٿ���#�@�"F,�4@�I�2�!?^3����@�Ûتٿ���#�@�"F,�4@�I�2�!?^3����@�Ûتٿ���#�@�"F,�4@�I�2�!?^3����@�Ûتٿ���#�@�"F,�4@�I�2�!?^3����@oZ}B��ٿه��N��@����4@��}�Q�!?�.���@oZ}B��ٿه��N��@����4@��}�Q�!?�.���@oZ}B��ٿه��N��@����4@��}�Q�!?�.���@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@���g�ٿ���4a�@Q���$ 4@�=$�!?a�f5k��@6��4��ٿ��{��#�@T'�� 4@lM*
��!?�<~��@6��4��ٿ��{��#�@T'�� 4@lM*
��!?�<~��@6��4��ٿ��{��#�@T'�� 4@lM*
��!?�<~��@��*�U�ٿ���D1��@8����3@��
�!?����*��@��*�U�ٿ���D1��@8����3@��
�!?����*��@��*�U�ٿ���D1��@8����3@��
�!?����*��@.���ٿZ�撉�@����2�3@|6>Տ!?t�Bb�@��<�ٿ`��C���@��B��3@�.C��!?�M�k��@��<�ٿ`��C���@��B��3@�.C��!?�M�k��@���F�ٿA*����@�9�M�3@�_���!?<XOܻ��@���F�ٿA*����@�9�M�3@�_���!?<XOܻ��@���F�ٿA*����@�9�M�3@�_���!?<XOܻ��@���F�ٿA*����@�9�M�3@�_���!?<XOܻ��@���F�ٿA*����@�9�M�3@�_���!?<XOܻ��@r���ٿ %��M �@7ۘ�3�3@K�˔��!?�i�T��@r���ٿ %��M �@7ۘ�3�3@K�˔��!?�i�T��@r���ٿ %��M �@7ۘ�3�3@K�˔��!?�i�T��@�R�x�ٿ$��w�_�@��B~�3@����	�!?�t��@�R�x�ٿ$��w�_�@��B~�3@����	�!?�t��@��
��ٿ<5�����@�qo�2 4@M��k�!?�_�ޖ��@��
��ٿ<5�����@�qo�2 4@M��k�!?�_�ޖ��@��
��ٿ<5�����@�qo�2 4@M��k�!?�_�ޖ��@��
��ٿ<5�����@�qo�2 4@M��k�!?�_�ޖ��@��
��ٿ<5�����@�qo�2 4@M��k�!?�_�ޖ��@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@c�B
��ٿf�W����@��	e�3@�9��c�!?w/��)�@�A!t�ٿ:51�=�@c�Re 4@P=r]�!?�\i��#�@1�$6�ٿ0�uN���@�|� 4@�󺌈�!?�+�F�\�@1�$6�ٿ0�uN���@�|� 4@�󺌈�!?�+�F�\�@1�$6�ٿ0�uN���@�|� 4@�󺌈�!?�+�F�\�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@�+y��ٿ]O�����@�̦s��3@��-J�!?�T­ߪ�@.�Q`F�ٿ��~�ת�@V-� 4@^8���!?�^\���@.�Q`F�ٿ��~�ת�@V-� 4@^8���!?�^\���@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���5��ٿ�{ŋ��@�S%� 4@0=���!?��m�.��@���
��ٿ0��Xσ�@b�9��3@u"uRԏ!?�3j����@���
��ٿ0��Xσ�@b�9��3@u"uRԏ!?�3j����@���
��ٿ0��Xσ�@b�9��3@u"uRԏ!?�3j����@���
��ٿ0��Xσ�@b�9��3@u"uRԏ!?�3j����@&�"��ٿ6Q,<Fd�@C��h��3@\��_d�!?�phz�q�@&�"��ٿ6Q,<Fd�@C��h��3@\��_d�!?�phz�q�@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@1�Ƨ2�ٿ *�2��@�sR���3@Ykv�n�!?&N�X��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@��S6,�ٿ���M:��@��^>* 4@(ɏ!?���ˉ��@�G�ͮٿ.���b��@w��\\ 4@H���ď!?���ۨ��@�G�ͮٿ.���b��@w��\\ 4@H���ď!?���ۨ��@�G�ͮٿ.���b��@w��\\ 4@H���ď!?���ۨ��@�G�ͮٿ.���b��@w��\\ 4@H���ď!?���ۨ��@\���%�ٿ_��v�@�
�!P�3@���͏!?�G�9L��@\���%�ٿ_��v�@�
�!P�3@���͏!?�G�9L��@\���%�ٿ_��v�@�
�!P�3@���͏!?�G�9L��@\���%�ٿ_��v�@�
�!P�3@���͏!?�G�9L��@\���%�ٿ_��v�@�
�!P�3@���͏!?�G�9L��@S:n���ٿKOd,���@n�]L 4@63?|�!?e�![�-�@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@FT��ٿv�?���@8�{�b 4@,Gr�!?
D,{��@4��-�ٿ��4�@�q��� 4@���f�!?w��0 �@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@�3B��ٿ:-gO�W�@I.� 4@qXkD��!?�ӓ���@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@V�/Si�ٿ�@�^���@u�_�4@�\U�!?�1Ch��@�B	Ϟٿ�r|̅-�@����3@X���a�!?G۬�8��@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@�dĝٿ��ܞ3�@���!� 4@�C�b�!? ���@)V��v�ٿO̾z��@m��Yf 4@ֳ��!?��AiI �@)V��v�ٿO̾z��@m��Yf 4@ֳ��!?��AiI �@)V��v�ٿO̾z��@m��Yf 4@ֳ��!?��AiI �@)V��v�ٿO̾z��@m��Yf 4@ֳ��!?��AiI �@�%��A�ٿy)o���@�)��� 4@Lk����!?Nc�qK��@�%��A�ٿy)o���@�)��� 4@Lk����!?Nc�qK��@�%��A�ٿy)o���@�)��� 4@Lk����!?Nc�qK��@�%��A�ٿy)o���@�)��� 4@Lk����!?Nc�qK��@�%��A�ٿy)o���@�)��� 4@Lk����!?Nc�qK��@��I�ٿ(3P�ы�@%�BoL�3@k�o͏!?;i�4u��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@4}66%�ٿ7�AEP�@#�% 4@�B��ڏ!?�Q�d��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@>�@��ٿxM�@^�@L��f~�3@�+��ُ!?H��V(��@|�3[��ٿ2�-0��@��Fj�3@J���׏!?]aG���@|�3[��ٿ2�-0��@��Fj�3@J���׏!?]aG���@|�3[��ٿ2�-0��@��Fj�3@J���׏!?]aG���@|�3[��ٿ2�-0��@��Fj�3@J���׏!?]aG���@3ܻ��ٿ�@D,���@pk/���3@�{_t��!?�!x����@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@��ɄZ�ٿ�zo�`�@�K�o9�3@H�(ꃏ!?�<�[`�@z�R*�ٿ��T��@6�2K 4@Ł
B��!?�5@��"�@z�R*�ٿ��T��@6�2K 4@Ł
B��!?�5@��"�@{����ٿt���o��@�ȧ�� 4@�a����!?�ō�1�@t�Ҍ>�ٿ��Np�@�5��64@��w��!?}�Z����@t�Ҍ>�ٿ��Np�@�5��64@��w��!?}�Z����@t�Ҍ>�ٿ��Np�@�5��64@��w��!?}�Z����@t�Ҍ>�ٿ��Np�@�5��64@��w��!?}�Z����@t�Ҍ>�ٿ��Np�@�5��64@��w��!?}�Z����@̐sX��ٿ�t>g~%�@V{�?�3@�:�Z�!?��/V��@̐sX��ٿ�t>g~%�@V{�?�3@�:�Z�!?��/V��@̐sX��ٿ�t>g~%�@V{�?�3@�:�Z�!?��/V��@��V+��ٿc�Ѡ�@)�BTW�3@���P{�!?�����@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@]�Lu�ٿ�G;�r6�@��_ˀ�3@���P�!?ִr�FZ�@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�e7>ʥٿ�L�p^I�@c�ˡ��3@�K�0a�!?GG���@�;u]�ٿ#����I�@� �iA�3@M�	MB�!?�`�)%�@�;u]�ٿ#����I�@� �iA�3@M�	MB�!?�`�)%�@�;u]�ٿ#����I�@� �iA�3@M�	MB�!?�`�)%�@��誋�ٿ�K�ă��@.��� 4@4�)�!?��3�'�@��誋�ٿ�K�ă��@.��� 4@4�)�!?��3�'�@��誋�ٿ�K�ă��@.��� 4@4�)�!?��3�'�@��誋�ٿ�K�ă��@.��� 4@4�)�!?��3�'�@4���J�ٿ�>�W��@Ϫ��� 4@��H+�!?=�ip��@4���J�ٿ�>�W��@Ϫ��� 4@��H+�!?=�ip��@�4� ٿYXY���@K���8�3@9�s�^�!?�A��e�@6��>�ٿ(Q\��n�@��M��3@�P��Y�!?ſ���@jZ~�;�ٿ���@�W94@���qs�!?�w�ώQ�@jZ~�;�ٿ���@�W94@���qs�!?�w�ώQ�@jZ~�;�ٿ���@�W94@���qs�!?�w�ώQ�@jZ~�;�ٿ���@�W94@���qs�!?�w�ώQ�@t�l�C�ٿ�������@]3��x�3@g�:��!?�K����@��5�[�ٿv枇V��@��� 4@j�MY��!?����� �@:1H�F�ٿ�-<޼g�@>y�W��3@V5L:܏!?ڶ�^��@:1H�F�ٿ�-<޼g�@>y�W��3@V5L:܏!?ڶ�^��@:1H�F�ٿ�-<޼g�@>y�W��3@V5L:܏!?ڶ�^��@:1H�F�ٿ�-<޼g�@>y�W��3@V5L:܏!?ڶ�^��@:1H�F�ٿ�-<޼g�@>y�W��3@V5L:܏!?ڶ�^��@����g�ٿ����G�@$�� �4@(��͏!?_-$��9�@����g�ٿ����G�@$�� �4@(��͏!?_-$��9�@����g�ٿ����G�@$�� �4@(��͏!?_-$��9�@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@)���ٿ�]���l�@.�4@!�i��!?�PHd���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@^���ٿi�P���@\���3@��G���!?�r�V���@~�y@�ٿ0iו��@�~K!,4@s�K}�!?��z;N��@~�y@�ٿ0iו��@�~K!,4@s�K}�!?��z;N��@~�y@�ٿ0iו��@�~K!,4@s�K}�!?��z;N��@~�y@�ٿ0iו��@�~K!,4@s�K}�!?��z;N��@~�y@�ٿ0iו��@�~K!,4@s�K}�!?��z;N��@�-c׬ٿ�V<�v�@��]N��3@X�����!?,fo���@�-c׬ٿ�V<�v�@��]N��3@X�����!?,fo���@�-c׬ٿ�V<�v�@��]N��3@X�����!?,fo���@�-c׬ٿ�V<�v�@��]N��3@X�����!?,fo���@�-c׬ٿ�V<�v�@��]N��3@X�����!?,fo���@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@��霨�ٿ�_�Ն��@n��mg 4@d�.v��!?S,�Lz��@S�`Xi�ٿ��h����@ƒ��3@������!?J�e�L�@!<r�ٿ��HS���@A9U��3@�=ɏ!?\G9�<��@!<r�ٿ��HS���@A9U��3@�=ɏ!?\G9�<��@!<r�ٿ��HS���@A9U��3@�=ɏ!?\G9�<��@���LH�ٿ�Nۮ���@yh0�0�3@$����!?��[��@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@��)���ٿ�&�٩��@����% 4@t� �!?����~�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@����ٿ��]C5i�@��x�G4@g�����!?�N��b�@{�3w��ٿW��l�@�㪜�4@�`r���!?�	�;)�@L��Z�ٿ�f�ɿs�@���X�4@�M,N~�!?q����@L��Z�ٿ�f�ɿs�@���X�4@�M,N~�!?q����@L��Z�ٿ�f�ɿs�@���X�4@�M,N~�!?q����@L��Z�ٿ�f�ɿs�@���X�4@�M,N~�!?q����@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@j�M�ٿ����@�@���i�4@���Q��!?�Kgp��@�׆L+�ٿt�@nb;�@�7��3@6$���!?������@�׆L+�ٿt�@nb;�@�7��3@6$���!?������@�׆L+�ٿt�@nb;�@�7��3@6$���!?������@6L��ٿMH!��@"�V�� 4@g ��)�!?�~��2��@6L��ٿMH!��@"�V�� 4@g ��)�!?�~��2��@6L��ٿMH!��@"�V�� 4@g ��)�!?�~��2��@��g���ٿ��,#h�@j�/4@���L�!?�ئE�@��S�m�ٿßD�@���+ 4@r0lJL�!?����
�@u�,\a�ٿKc���@	k��4@�=3l�!?��߬�@u�,\a�ٿKc���@	k��4@�=3l�!?��߬�@u�,\a�ٿKc���@	k��4@�=3l�!?��߬�@�k�Oݲٿ�D0���@�׹E 4@I�)��!?B�����@(�:ȩٿ˾m�F��@-�[Ȓ4@v�G��!?��Pq��@(�:ȩٿ˾m�F��@-�[Ȓ4@v�G��!?��Pq��@(�:ȩٿ˾m�F��@-�[Ȓ4@v�G��!?��Pq��@(�:ȩٿ˾m�F��@-�[Ȓ4@v�G��!?��Pq��@��y�H�ٿ&<5�k�@Q+T 4@x�;��!?�$7�y�@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@�a�
��ٿW��G�&�@�oA�4@4��}��!?������@2�D�ٿn���-�@t��4@�>�1��!?W<��@!����ٿ��1
��@�2*B�4@�[tT�!?��T��@!����ٿ��1
��@�2*B�4@�[tT�!?��T��@��wk�ٿ�JG��@U(%�G4@�H�D�!?X�`�`�@��wk�ٿ�JG��@U(%�G4@�H�D�!?X�`�`�@���}\�ٿ7���G^�@� � 4@��a��!?M�
�3N�@���}\�ٿ7���G^�@� � 4@��a��!?M�
�3N�@���}\�ٿ7���G^�@� � 4@��a��!?M�
�3N�@_�Aڦٿh�A�w�@z��4@���	h�!?Rl+�nL�@_�Aڦٿh�A�w�@z��4@���	h�!?Rl+�nL�@_�Aڦٿh�A�w�@z��4@���	h�!?Rl+�nL�@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@B���Ģٿ�P�i��@��M�4@?��.��!?����O��@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@������ٿ튱���@I���>4@"�lԏ!?�%����@��g2M�ٿ�òߩY�@���L4@�)����!?1dz�ڸ�@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@���)y�ٿi�w��@i���4@�E s�!?0�<_���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@�4��ٿ���ie�@*UFD��3@Ws�Ə!?���@;k��ٿ셁=��@�7 4@'E�ʏ!?���xw{�@;k��ٿ셁=��@�7 4@'E�ʏ!?���xw{�@EoK��ٿ*�z(��@i�w4@�~;g�!?	o����@h�%鋰ٿ��]${��@ؘee� 4@pP+^�!?�@NŁ�@h�%鋰ٿ��]${��@ؘee� 4@pP+^�!?�@NŁ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@c�@��ٿZ�0.�@q��% 4@�KM�y�!?n�6�ӷ�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@��ջ��ٿf~"t��@ƶ4]{4@J��I��!?�s��>�@�氰��ٿe�w	�@�O�24@�qwQ�!?x�>	�@Oȥٿ8��x��@�&ɩ��3@�e���!?`>����@Oȥٿ8��x��@�&ɩ��3@�e���!?`>����@9�p���ٿW�C�@ �@m۲fy�3@r�"�ӏ!?��6�8�@�m���ٿ�p���@�ih̃4@x�r���!?�K����@�m���ٿ�p���@�ih̃4@x�r���!?�K����@�m���ٿ�p���@�ih̃4@x�r���!?�K����@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@�nP���ٿ�$MA\�@L��4@�>Q͏!? ���=��@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@8�`���ٿ�.�c���@�m]��4@�Z����!?x򗕸/�@'y0A�ٿڌ�|��@��Y���3@����Ï!?�0�����@'y0A�ٿڌ�|��@��Y���3@����Ï!?�0�����@'y0A�ٿڌ�|��@��Y���3@����Ï!?�0�����@'y0A�ٿڌ�|��@��Y���3@����Ï!?�0�����@'y0A�ٿڌ�|��@��Y���3@����Ï!?�0�����@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@���+�ٿ��M���@1�9�� 4@���ֺ�!?X�X�G��@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@.���ٿ���w��@.o$D 4@�x`��!?h��!� �@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@�\IH?�ٿR����@���p 4@�s���!?�e+��@���fɗٿ��P���@w��F��3@�@�3��!?�/�%Ձ�@���fɗٿ��P���@w��F��3@�@�3��!?�/�%Ձ�@��pR��ٿ��t����@�cJe� 4@��I���!?����V�@'�-+��ٿP+2�³�@ˑ�3@�d���!?��1��@'�-+��ٿP+2�³�@ˑ�3@�d���!?��1��@O���)�ٿƿo�h��@��(%S 4@�M�r�!?�0R�u�@ISt��ٿ��u\��@L؆O� 4@A�Y�!?F�z)�@)��ЖٿS�LA��@T�7��4@�^�6��!?B�#.���@)��ЖٿS�LA��@T�7��4@�^�6��!?B�#.���@)��ЖٿS�LA��@T�7��4@�^�6��!?B�#.���@)��ЖٿS�LA��@T�7��4@�^�6��!?B�#.���@w]���ٿy�K	?��@>E364@AH�!?(�SiI�@���M��ٿ�uג�o�@�|x� 4@vL��׏!?�z|���@���M��ٿ�uג�o�@�|x� 4@vL��׏!?�z|���@�=�Ud�ٿa_��E��@V#B�F 4@ECr���!?�k��'�@�=�Ud�ٿa_��E��@V#B�F 4@ECr���!?�k��'�@�=�Ud�ٿa_��E��@V#B�F 4@ECr���!?�k��'�@.���ٿ�G�O�`�@�:���3@�D:��!?��e�JY�@.���ٿ�G�O�`�@�:���3@�D:��!?��e�JY�@.���ٿ�G�O�`�@�:���3@�D:��!?��e�JY�@.���ٿ�G�O�`�@�:���3@�D:��!?��e�JY�@~O��}�ٿ��ڭ��@��� 4@|E���!?�zj����@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@��<ۥٿ��>���@�pm�$4@- �	��!?�6k{��@/*\, �ٿ��l����@#���4@;bє�!?̍�\�#�@�"b�Y�ٿ��k���@�/w�14@�s���!?9����.�@�"b�Y�ٿ��k���@�/w�14@�s���!?9����.�@�"b�Y�ٿ��k���@�/w�14@�s���!?9����.�@�"b�Y�ٿ��k���@�/w�14@�s���!?9����.�@�"b�Y�ٿ��k���@�/w�14@�s���!?9����.�@t`�Q�ٿ��f�+4�@��u3�4@7W,]�!?U���K��@t`�Q�ٿ��f�+4�@��u3�4@7W,]�!?U���K��@t`�Q�ٿ��f�+4�@��u3�4@7W,]�!?U���K��@t`�Q�ٿ��f�+4�@��u3�4@7W,]�!?U���K��@t`�Q�ٿ��f�+4�@��u3�4@7W,]�!?U���K��@���A�ٿ���P��@e�?s�4@'Zޜg�!?K��8N�@���A�ٿ���P��@e�?s�4@'Zޜg�!?K��8N�@���A�ٿ���P��@e�?s�4@'Zޜg�!?K��8N�@��@?�ٿK�@R��@�qT�; 4@���(;�!?�9@z��@� ֟ٿA?�N�@u�f�4@A��j�!?s�ԭ���@� ֟ٿA?�N�@u�f�4@A��j�!?s�ԭ���@R�_�ٿ�Q��@����4@�fُ!?��3��P�@R�_�ٿ�Q��@����4@�fُ!?��3��P�@R�_�ٿ�Q��@����4@�fُ!?��3��P�@R�_�ٿ�Q��@����4@�fُ!?��3��P�@R�_�ٿ�Q��@����4@�fُ!?��3��P�@s�;�_�ٿ5�7�w�@p�h�4@���W�!?�@�v��@s�;�_�ٿ5�7�w�@p�h�4@���W�!?�@�v��@s�;�_�ٿ5�7�w�@p�h�4@���W�!?�@�v��@s�;�_�ٿ5�7�w�@p�h�4@���W�!?�@�v��@l�vÀ�ٿ��?8��@I�y824@k�
(�!?�y��B!�@l�vÀ�ٿ��?8��@I�y824@k�
(�!?�y��B!�@l�vÀ�ٿ��?8��@I�y824@k�
(�!?�y��B!�@�4�zS�ٿ��4����@�XV��4@~]Cߏ!?.�l�!�@�4�zS�ٿ��4����@�XV��4@~]Cߏ!?.�l�!�@qUV��ٿ��W����@���N4@l�3�!?ܲ�[��@qUV��ٿ��W����@���N4@l�3�!?ܲ�[��@�����ٿ��[�@ؿ؍1 4@�}�Kԏ!?�v�Sy�@�����ٿ��[�@ؿ؍1 4@�}�Kԏ!?�v�Sy�@�����ٿ��[�@ؿ؍1 4@�}�Kԏ!?�v�Sy�@�����ٿ��[�@ؿ؍1 4@�}�Kԏ!?�v�Sy�@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@��6�ٿ~��1c5�@j?��4@��]��!?a��J��@���4;�ٿ4{�u�@��e4@g;ŏ!?j^C��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@�R[;�ٿ!!['�@�9�W��3@x�,���!?���l��@� �I[�ٿ4M
k�g�@��?[�4@�(�ʏ!?��Y@
U�@� �I[�ٿ4M
k�g�@��?[�4@�(�ʏ!?��Y@
U�@� �I[�ٿ4M
k�g�@��?[�4@�(�ʏ!?��Y@
U�@� �I[�ٿ4M
k�g�@��?[�4@�(�ʏ!?��Y@
U�@� �I[�ٿ4M
k�g�@��?[�4@�(�ʏ!?��Y@
U�@�+�b�ٿ��?���@�'е/4@�ԟď!?h~��G4�@�+�b�ٿ��?���@�'е/4@�ԟď!?h~��G4�@�+�b�ٿ��?���@�'е/4@�ԟď!?h~��G4�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@,�^�6�ٿ�!K�d��@���F�4@�O`͏!?�r�D
V�@�-�[�ٿ=�h�P��@G�l�' 4@�<=��!?Q���D�@�-�[�ٿ=�h�P��@G�l�' 4@�<=��!?Q���D�@�-�[�ٿ=�h�P��@G�l�' 4@�<=��!?Q���D�@�Ԩ(�ٿ�q�&x��@[>�h�3@F��!?��(�'�@�Ԩ(�ٿ�q�&x��@[>�h�3@F��!?��(�'�@�Ԩ(�ٿ�q�&x��@[>�h�3@F��!?��(�'�@�Ԩ(�ٿ�q�&x��@[>�h�3@F��!?��(�'�@�Ԩ(�ٿ�q�&x��@[>�h�3@F��!?��(�'�@�����ٿ#s�u�+�@�z��� 4@E��Ao�!?M81٨�@�����ٿ#s�u�+�@�z��� 4@E��Ao�!?M81٨�@�����ٿ#s�u�+�@�z��� 4@E��Ao�!?M81٨�@�����ٿ#s�u�+�@�z��� 4@E��Ao�!?M81٨�@�����ٿ#s�u�+�@�z��� 4@E��Ao�!?M81٨�@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��B�Щٿ�]�]J��@ 5�o4@�̇o�!?����@��S�2�ٿ%�-��@�4{��4@�y6|��!?�N���@��S�2�ٿ%�-��@�4{��4@�y6|��!?�N���@#Af���ٿ�Ӏf���@�3. 4@���G��!?h�V��@#Af���ٿ�Ӏf���@�3. 4@���G��!?h�V��@#Af���ٿ�Ӏf���@�3. 4@���G��!?h�V��@#Af���ٿ�Ӏf���@�3. 4@���G��!?h�V��@o̊L��ٿOCј��@'��4@�b&��!?�K��.T�@o̊L��ٿOCј��@'��4@�b&��!?�K��.T�@o̊L��ٿOCј��@'��4@�b&��!?�K��.T�@o̊L��ٿOCј��@'��4@�b&��!?�K��.T�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@U�\q*�ٿ��Om��@�B �94@��]/ɏ!?���Fs�@���<�ٿ��]�>��@�f 4@?Hb~��!?b��̚-�@����ڠٿ{j��T��@![\4� 4@�GH��!?$�a�u+�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@���!�ٿ������@*��s��3@љ���!?#] 30�@}�*���ٿ��5��@��*4@*?��ȏ!?���x���@}�*���ٿ��5��@��*4@*?��ȏ!?���x���@}�*���ٿ��5��@��*4@*?��ȏ!?���x���@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@J���#�ٿt	�9 ��@A�)Lk 4@�Z$�!?��8�Bb�@Tʑ�o�ٿ4Ɲ��D�@��!�4@!S^b�!?�4��	�@�b�n�ٿl���%�@��y64@`�͏!?X�����@�b�n�ٿl���%�@��y64@`�͏!?X�����@�b�n�ٿl���%�@��y64@`�͏!?X�����@�b�n�ٿl���%�@��y64@`�͏!?X�����@�b�n�ٿl���%�@��y64@`�͏!?X�����@�b�n�ٿl���%�@��y64@`�͏!?X�����@�����ٿ꜇V��@�I&��4@7[`ɏ!?�٘U0��@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�A���ٿf��	��@-$pj 4@TݮOɏ!?g�*�L�@�HL�;�ٿ�B����@���j� 4@�G+��!??��H��@Y깮9�ٿ����O�@A��	 4@���q��!? ���@m�4ϴ�ٿGf1|+�@}�$ 4@A�o���!?L���]�@m�4ϴ�ٿGf1|+�@}�$ 4@A�o���!?L���]�@��@�
�ٿX��1��@�$'cq 4@h�=B��!?�4�F2�@��@�
�ٿX��1��@�$'cq 4@h�=B��!?�4�F2�@A��v�ٿ��г�@�T���3@S�S�!?`����@�@��E�s�ٿ`A�֒�@U�0���3@)��-�!?C�Ei�@����{�ٿ��'4�@����3@kW�É�!?;n�6���@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@P�=5��ٿ��*�@�,����3@=��岏!?��3�
�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@͐n���ٿ�@���@=�h� 4@�᭟_�!?�=L�~?�@;��"�ٿԯ@B�
�@�6ۄ�4@q|1h~�!?�Y��=�@jL2��ٿ5�"�- �@��!�4@z�(ɏ!? ~��A��@jL2��ٿ5�"�- �@��!�4@z�(ɏ!? ~��A��@��XD�ٿ����A�@�=���4@����d�!?;��o�:�@,����ٿfVq����@�.�9-4@qjm���!?�i�l@�@,����ٿfVq����@�.�9-4@qjm���!?�i�l@�@,����ٿfVq����@�.�9-4@qjm���!?�i�l@�@�B��ٿB�-9�k�@�Y�4@�y�eG�!?�N\8�@�B��ٿB�-9�k�@�Y�4@�y�eG�!?�N\8�@~��~�ٿ�$�f�t�@�5�4@���9�!?5).��@~��~�ٿ�$�f�t�@�5�4@���9�!?5).��@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@P��q��ٿ�n]̌�@଄��4@�g�!?/O����@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@�t��ٿwp����@�-��� 4@��qE�!?�KXHă�@��cW�ٿ�ԓ���@^/B(�3@g �c�!?G� ����@��cW�ٿ�ԓ���@^/B(�3@g �c�!?G� ����@��cW�ٿ�ԓ���@^/B(�3@g �c�!?G� ����@�^_���ٿ|����@T�f���3@�l��u�!?Yi����@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@u�Zb��ٿ�y9���@<Y� 14@b����!? �&��~�@P���ٿ�`+Vl�@'#�{�4@�z嚏!?�5P�k��@]ҩ%�ٿ�/�R��@sk3?!4@ܥ iߏ!?W����j�@]ҩ%�ٿ�/�R��@sk3?!4@ܥ iߏ!?W����j�@�)q��ٿ�Y����@>bg�4@m�R��!?{v�����@�)q��ٿ�Y����@>bg�4@m�R��!?{v�����@D�
c��ٿ�a<e#�@��s��4@�	���!?1+@�ˑ�@D�
c��ٿ�a<e#�@��s��4@�	���!?1+@�ˑ�@նM�9�ٿwAڼRc�@��Z��3@`kݵ�!?3K*���@նM�9�ٿwAڼRc�@��Z��3@`kݵ�!?3K*���@նM�9�ٿwAڼRc�@��Z��3@`kݵ�!?3K*���@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@7Ķ���ٿ�7\a�&�@�Q�x��3@��^��!?���v��@8T���ٿ��,jփ�@]�`O�4@��v���!?��!����@8T���ٿ��,jփ�@]�`O�4@��v���!?��!����@8T���ٿ��,jփ�@]�`O�4@��v���!?��!����@8T���ٿ��,jփ�@]�`O�4@��v���!?��!����@����ٿl(
줽�@��	�4@/cyk�!?�4�կ�@����ٿl(
줽�@��	�4@/cyk�!?�4�կ�@����ٿl(
줽�@��	�4@/cyk�!?�4�կ�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@�h����ٿ�z.���@PC�� 4@���!?���	�@��{�P�ٿ�3��m�@�k�ȧ�3@:�_D�!?A���Û�@��{�P�ٿ�3��m�@�k�ȧ�3@:�_D�!?A���Û�@��{�P�ٿ�3��m�@�k�ȧ�3@:�_D�!?A���Û�@f���ٿl����_�@�0��M 4@��ࡏ!?���'��@f���ٿl����_�@�0��M 4@��ࡏ!?���'��@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@��07��ٿ��٪@�@�W�� 4@⪨&r�!?����j�@�� � �ٿ���(�@���V��3@A\���!?�t��m��@�����ٿ � Y���@�K�!��3@��gϢ�!?0�?���@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@�R�?�ٿ���*j��@Pt�%��3@�O���!?���،�@���3M�ٿ���)˱�@�����3@� �f�!?ؾ�&�T�@���3M�ٿ���)˱�@�����3@� �f�!?ؾ�&�T�@���3M�ٿ���)˱�@�����3@� �f�!?ؾ�&�T�@���3M�ٿ���)˱�@�����3@� �f�!?ؾ�&�T�@�v谣ٿ��Wr6��@�	��'�3@�ͪ^�!?���7�@�v谣ٿ��Wr6��@�	��'�3@�ͪ^�!?���7�@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@U�,�ٿELC~�@'o>�� 4@���s�!?�|T���@�CV��ٿ��@��W�4@z�Mi��!?-m�\��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@5y8��ٿH3j0%��@=r�-4@ּH��!?^�(��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@��5g��ٿ�,��p�@;��sn 4@ �j��!?0��G*��@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@Ea&��ٿR�s`F{�@�<�c 4@IK�Jq�!?��:�Ĥ�@�P�Ų�ٿ�+�dZ�@	����3@����!?�ȇ(1�@�P�Ų�ٿ�+�dZ�@	����3@����!?�ȇ(1�@�P�Ų�ٿ�+�dZ�@	����3@����!?�ȇ(1�@�P�Ų�ٿ�+�dZ�@	����3@����!?�ȇ(1�@�P�Ų�ٿ�+�dZ�@	����3@����!?�ȇ(1�@�:��F�ٿ*G�nk�@I�6],�3@���!?7:b_�@�:��F�ٿ*G�nk�@I�6],�3@���!?7:b_�@�:��F�ٿ*G�nk�@I�6],�3@���!?7:b_�@�:��F�ٿ*G�nk�@I�6],�3@���!?7:b_�@E4��ٿ�'��@��˥ 4@�����!?[6I�`�@E4��ٿ�'��@��˥ 4@�����!?[6I�`�@E4��ٿ�'��@��˥ 4@�����!?[6I�`�@E4��ٿ�'��@��˥ 4@�����!?[6I�`�@E4��ٿ�'��@��˥ 4@�����!?[6I�`�@���y��ٿ���I�@�(����3@=����!?��ⷯ��@���y��ٿ���I�@�(����3@=����!?��ⷯ��@;;�v�ٿx#5�|�@tˆ�(�3@�xZ4��!?B��V��@;;�v�ٿx#5�|�@tˆ�(�3@�xZ4��!?B��V��@;;�v�ٿx#5�|�@tˆ�(�3@�xZ4��!?B��V��@��%W[�ٿ7p=LW�@ �J�� 4@���I�!?ؼ�1�R�@g�r�'�ٿ/"��1�@x�Y��4@#��И�!?.��*��@˩��ٿʎ�8(�@�L���3@��<Xӏ!?M�©�)�@��&�ٿge�@d�ht�3@���!?�?�����@����ٿ��P��@qLԖ��3@���!?�>����@Ķ5�;�ٿ�<j��u�@��q��3@�1K>�!?ʬΨO�@���Śٿ��T>;�@��ˬ�3@ܯc��!?8{�����@���Śٿ��T>;�@��ˬ�3@ܯc��!?8{�����@���Śٿ��T>;�@��ˬ�3@ܯc��!?8{�����@��2�ٿ� �#B��@�y��H�3@z���4�!?�7���}�@�3�/ �ٿ�/?:��@�Qȝ; 4@X�����!?ZnE��@�3�/ �ٿ�/?:��@�Qȝ; 4@X�����!?ZnE��@�3�/ �ٿ�/?:��@�Qȝ; 4@X�����!?ZnE��@�3�/ �ٿ�/?:��@�Qȝ; 4@X�����!?ZnE��@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@��-��ٿ�P�l�@���F) 4@o�b��!?�b��	�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@^=G8�ٿ�h:X~��@���x� 4@������!?ա��E�@��r�M�ٿ;p�o)��@�=紷�3@?̄ϓ�!?�`�l���@��r�M�ٿ;p�o)��@�=紷�3@?̄ϓ�!?�`�l���@��r�M�ٿ;p�o)��@�=紷�3@?̄ϓ�!?�`�l���@:�0�;�ٿ��
}��@Xu��<�3@Έ�Q}�!?�=U����@:�0�;�ٿ��
}��@Xu��<�3@Έ�Q}�!?�=U����@:�0�;�ٿ��
}��@Xu��<�3@Έ�Q}�!?�=U����@:�0�;�ٿ��
}��@Xu��<�3@Έ�Q}�!?�=U����@7�P4�ٿ������@��'r��3@��h�
�!?�k�~o�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@�L��=�ٿ~ yG�@VRw/F 4@�QL�U�!?���K�K�@o޸s�ٿ(G�n��@u�F��3@]�{ԏ!?dz+/�@o޸s�ٿ(G�n��@u�F��3@]�{ԏ!?dz+/�@o޸s�ٿ(G�n��@u�F��3@]�{ԏ!?dz+/�@o޸s�ٿ(G�n��@u�F��3@]�{ԏ!?dz+/�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@��r�ٿ�C=`p�@�*��3@���	��!?4;�˝�@Z��M�ٿR�l��t�@e�d� 4@N����!?����@Z��M�ٿR�l��t�@e�d� 4@N����!?����@P��#�ٿ�I��q�@6��5 4@���� �!?��`j��@P��#�ٿ�I��q�@6��5 4@���� �!?��`j��@P��#�ٿ�I��q�@6��5 4@���� �!?��`j��@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@������ٿ����y�@��
V 4@l�R/�!?7�w�ZP�@b�7�ٿ��*�W�@o#)���3@��
�!?D������@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@��x6_�ٿ�h��9�@���ڵ 4@�qXu{�!?�h? q�@Y�8��ٿ�;��!�@~���P4@�e��a�!?wM��
�@Y�8��ٿ�;��!�@~���P4@�e��a�!?wM��
�@Y�8��ٿ�;��!�@~���P4@�e��a�!?wM��
�@Y�8��ٿ�;��!�@~���P4@�e��a�!?wM��
�@Y�8��ٿ�;��!�@~���P4@�e��a�!?wM��
�@���U��ٿf"�u�`�@L	�4@3
7�o�!?S:%���@���U��ٿf"�u�`�@L	�4@3
7�o�!?S:%���@���U��ٿf"�u�`�@L	�4@3
7�o�!?S:%���@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�䵠H�ٿ�/: 9.�@��3��3@��ք��!?�ܦx��@�ZOp��ٿ�y�-�@G���! 4@���X\�!?2���X�@�ZOp��ٿ�y�-�@G���! 4@���X\�!?2���X�@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@�H{]�ٿ�.�uHg�@���>7 4@�F#���!?�m�I��@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��o<�ٿٛ�|0t�@jF�� 4@�~���!?r�Ԗ�@��Y�ٿ9�R����@�ߜ;�4@�A����!?�n���@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@��Ȕ��ٿ�ڗ����@7TmCK4@G{�e�!?��&
F�@�g��ٿ�}���@Hh��u4@�gi��!?�QO����@�g��ٿ�}���@Hh��u4@�gi��!?�QO����@�4���ٿ�I0at%�@�V��F4@�s��ߏ!?b�9v|��@�4���ٿ�I0at%�@�V��F4@�s��ߏ!?b�9v|��@z��ȯٿ22�N���@��f| 4@���U��!?�����<�@�7=g�ٿ���V;�@���W�3@Z&v�o�!?�YI�E�@�7=g�ٿ���V;�@���W�3@Z&v�o�!?�YI�E�@�;�3y�ٿ��Z��@���	&�3@?�{v�!?�چ�@�h����ٿ7�i��I�@��5r	 4@�v�Y��!?��=#�S�@�h����ٿ7�i��I�@��5r	 4@�v�Y��!?��=#�S�@�h����ٿ7�i��I�@��5r	 4@�v�Y��!?��=#�S�@�h����ٿ7�i��I�@��5r	 4@�v�Y��!?��=#�S�@i�?I�ٿ�\����@��) 4@2�*6�!?��͊�@�`�*�ٿd,7��U�@�8�� 4@,sHƏ!?&���[�@�`�*�ٿd,7��U�@�8�� 4@,sHƏ!?&���[�@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@��Wm�ٿ��g#��@�����3@Dg��!?�]�N��@�އ5�ٿL��=�@�/HZ�3@�Qj�!?@��Ȅ��@�އ5�ٿL��=�@�/HZ�3@�Qj�!?@��Ȅ��@�އ5�ٿL��=�@�/HZ�3@�Qj�!?@��Ȅ��@U'���ٿ��=�
��@\: ���3@��ď!?EV~٧��@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@�ݤn�ٿ|�#�E3�@�er 4@�.����!?��S�>N�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@l�In[�ٿ�F���@�;1 4@Asf_�!?��{�ٰ�@w�@���ٿ��{u��@c�բ� 4@�g?��!?�yI��@w�@���ٿ��{u��@c�բ� 4@�g?��!?�yI��@�x�4��ٿ��yK�E�@�(�� 4@\J8���!?��3��g�@�x�4��ٿ��yK�E�@�(�� 4@\J8���!?��3��g�@�x�4��ٿ��yK�E�@�(�� 4@\J8���!?��3��g�@���Z�ٿW�����@��U 4@ �>�!?E���.�@�X��ٿ<��o��@:y���3@�I�!�!?8i�t���@�X��ٿ<��o��@:y���3@�I�!�!?8i�t���@�X��ٿ<��o��@:y���3@�I�!�!?8i�t���@�m�G�ٿ<v%�v��@��V� 4@ qPO�!?�}��aI�@�}�ٿ����:�@�,��`4@���{6�!?�^�i��@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@�v���ٿ�����@�?�F� 4@{�h�/�!?�%�_���@��*�"�ٿ(�!����@uuk�� 4@�SV��!?�-�t�@h�OT/�ٿg�`W���@���Ü 4@>���$�!?ϔ3�):�@h�OT/�ٿg�`W���@���Ü 4@>���$�!?ϔ3�):�@h�OT/�ٿg�`W���@���Ü 4@>���$�!?ϔ3�):�@C��ޥٿd+0�q�@ܺ�`��3@(#�R��!?�M���@L���ٿd�%6X�@5aF�� 4@�'�G��!?%Z�@��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@y�℥ٿ�'l�q\�@i0�@� 4@��]_Տ!?��
yT��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@���ʤٿ���_*�@ep�(4@�V"�Ə!?�}�H��@�({6t�ٿ&z�!��@)Jғ1 4@��Ñ�!?�>��/��@�-��u�ٿ��w���@~w��4@�Mj�ŏ!?��Z���@�-��u�ٿ��w���@~w��4@�Mj�ŏ!?��Z���@�-��u�ٿ��w���@~w��4@�Mj�ŏ!?��Z���@�-��u�ٿ��w���@~w��4@�Mj�ŏ!?��Z���@(���ٿ4��k�@ZS0��4@��4w�!?�$����@Oxݫ��ٿ��9���@��cb4@e ���!?bJ��~[�@Oxݫ��ٿ��9���@��cb4@e ���!?bJ��~[�@n갧Ŕٿ�.�%H&�@�}�o 4@Ei�IǏ!?������@n갧Ŕٿ�.�%H&�@�}�o 4@Ei�IǏ!?������@n갧Ŕٿ�.�%H&�@�}�o 4@Ei�IǏ!?������@n갧Ŕٿ�.�%H&�@�}�o 4@Ei�IǏ!?������@n갧Ŕٿ�.�%H&�@�}�o 4@Ei�IǏ!?������@��:���ٿ������@V�&���3@�%.x��!?A)�y�%�@��:���ٿ������@V�&���3@�%.x��!?A)�y�%�@��:���ٿ������@V�&���3@�%.x��!?A)�y�%�@��:���ٿ������@V�&���3@�%.x��!?A)�y�%�@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@�2��h�ٿ�o=���@v��K?�3@Qy�*��!?���9��@J���ٿ��4l�@��Fe�3@V]i�!?�����@�t�*ʙٿ�rل��@�ߙZy 4@�g��!?�
SbH�@w�殥ٿ&S�}���@c� (>4@~E��!?N��a�@=r��ٿ�/�-���@��HQ4@�����!?�ɐ�s�@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@i~�w�ٿ�p��e�@q�J�4@�Qຏ!?��S��@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@��ڼb�ٿ*>��j�@ٌ��i4@�gZ[Ï!?@JJ��Y�@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@�uс�ٿ�)��}�@�ù�y4@� >=��!?�`Ϯ���@ں��ٿ���Cz��@Q��cy4@,��w�!?�	�	���@ں��ٿ���Cz��@Q��cy4@,��w�!?�	�	���@ں��ٿ���Cz��@Q��cy4@,��w�!?�	�	���@�#��ͩٿ��k%�@&��t 4@jUҏ!?\�w����@Vb�@��ٿ��R����@�޽�4@�����!?�����-�@Vb�@��ٿ��R����@�޽�4@�����!?�����-�@Vb�@��ٿ��R����@�޽�4@�����!?�����-�@Vb�@��ٿ��R����@�޽�4@�����!?�����-�@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@�*�L�ٿ��QU~�@^x�04@ �u֏!?�pf�P��@ܶfn�ٿ6�0 hb�@&��H4@�����!?�k�N���@ܶfn�ٿ6�0 hb�@&��H4@�����!?�k�N���@
Ċs�ٿ�i,�Vz�@��� 4@�F���!?���d�@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@��fB*�ٿ&c��;��@�� 4@qT�k�!?�ȟ���@U�?�ٿ�-`=0�@���}^ 4@R�250�!?�7E��D�@U�?�ٿ�-`=0�@���}^ 4@R�250�!?�7E��D�@U�?�ٿ�-`=0�@���}^ 4@R�250�!?�7E��D�@U�?�ٿ�-`=0�@���}^ 4@R�250�!?�7E��D�@U�?�ٿ�-`=0�@���}^ 4@R�250�!?�7E��D�@]5Z�ٿ� W���@��ͧ! 4@������!?�0[$0h�@]5Z�ٿ� W���@��ͧ! 4@������!?�0[$0h�@]5Z�ٿ� W���@��ͧ! 4@������!?�0[$0h�@]5Z�ٿ� W���@��ͧ! 4@������!?�0[$0h�@0��8�ٿk�����@�Ŝ7��3@
��s�!?Z������@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@�8g�U�ٿϑwhѢ�@VD����3@�����!?b��W��@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@_��@L�ٿ/�mq{��@�i�6 4@��,Տ!?xǌ���@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@�"���ٿ��m0��@�V:O4@t��T�!?�U�ٟ�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@Te�V�ٿ٦k�s�@|�X��3@9�x�!?�2 ��]�@FL+%ٞٿ!�ɢ�8�@�D6��3@7c�o��!?�_���@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@��-�ٿo�-�|Y�@����4@��GU��!?NZ�w��@�>vp�ٿ��X�f�@bJ�ݾ�3@�X�1��!?Go_yҜ�@-��C��ٿ�Ȧ8�@8,���3@~*㪏!?lX��S�@���E�ٿ����U��@��*��3@� �p��!?��,VI�@���E�ٿ����U��@��*��3@� �p��!?��,VI�@���E�ٿ����U��@��*��3@� �p��!?��,VI�@���E�ٿ����U��@��*��3@� �p��!?��,VI�@���E�ٿ����U��@��*��3@� �p��!?��,VI�@+=I<�ٿ~/��l�@��m]�3@��c���!?z�YSgj�@Lm ~��ٿݺ�Z�S�@���� 4@��7Џ!?�Xxͭs�@Lm ~��ٿݺ�Z�S�@���� 4@��7Џ!?�Xxͭs�@Lm ~��ٿݺ�Z�S�@���� 4@��7Џ!?�Xxͭs�@Lm ~��ٿݺ�Z�S�@���� 4@��7Џ!?�Xxͭs�@�9��ٿI����E�@��G#F4@g�eз�!?����]c�@�9��ٿI����E�@��G#F4@g�eз�!?����]c�@�9��ٿI����E�@��G#F4@g�eз�!?����]c�@�9��ٿI����E�@��G#F4@g�eз�!?����]c�@�9��ٿI����E�@��G#F4@g�eз�!?����]c�@�,�}\�ٿ��b7���@�f���3@�Gi�W�!?G�h��@�,�}\�ٿ��b7���@�f���3@�Gi�W�!?G�h��@T]nƲٿ�'7�
��@�0�x��3@��3�z�!?��:Y���@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@ɟj��ٿ����w@�@�|	 4@����`�!?�
�C]+�@���Λٿ�W����@�\���3@�u��p�!?;f�����@���Λٿ�W����@�\���3@�u��p�!?;f�����@���Λٿ�W����@�\���3@�u��p�!?;f�����@ӡ/L5�ٿ��6rc�@K�r�3@�Ӽd��!?�J���@��Vw�ٿ��p�a�@:�L��3@^0ϵڏ!?��"��@ą����ٿ��C�z��@tr��z�3@����!?JX��@ą����ٿ��C�z��@tr��z�3@����!?JX��@ą����ٿ��C�z��@tr��z�3@����!?JX��@ą����ٿ��C�z��@tr��z�3@����!?JX��@ą����ٿ��C�z��@tr��z�3@����!?JX��@͛��ޡٿr�hP�@��^g 4@�ˊ��!?�&�\d�@͛��ޡٿr�hP�@��^g 4@�ˊ��!?�&�\d�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��$Tr�ٿ6K��D�@�]]IT 4@���B׏!?ˤ~Zݹ�@��4~�ٿ��Dd��@%��� 4@C�<$�!?A�W�b~�@*,�&�ٿ�BM���@�Tob4@��t��!?5}���@ .�B��ٿ+��>M��@S�KB54@���!?��FqN��@ .�B��ٿ+��>M��@S�KB54@���!?��FqN��@�Xf��ٿ��&�k�@v�����3@w��Tя!?gC��}�@d#��ٿjl+}��@�Lge 4@����!?3�X�Ԉ�@d#��ٿjl+}��@�Lge 4@����!?3�X�Ԉ�@d#��ٿjl+}��@�Lge 4@����!?3�X�Ԉ�@d#��ٿjl+}��@�Lge 4@����!?3�X�Ԉ�@.-:nt�ٿ�:z?��@r�u���3@O�-ŏ!?(�-p�@.-:nt�ٿ�:z?��@r�u���3@O�-ŏ!?(�-p�@.-:nt�ٿ�:z?��@r�u���3@O�-ŏ!?(�-p�@.-:nt�ٿ�:z?��@r�u���3@O�-ŏ!?(�-p�@�8~���ٿ?<~���@"c���3@���0ȏ!?Ɇ��	�@�8~���ٿ?<~���@"c���3@���0ȏ!?Ɇ��	�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@g�3f��ٿI���?]�@��";~�3@e�v�!?[��+�@tC'&��ٿo�lh�@c}� ��3@�J�l��!?ߤW��"�@�sޘ��ٿX"�G2�@�m����3@��}���!?�M+��@�A�(g�ٿx��r�i�@=��˥�3@)�T6O�!?n�7��@vI�ާٿa�����@�Wi��3@w�<��!?p�N:�Q�@vI�ާٿa�����@�Wi��3@w�<��!?p�N:�Q�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@~���B�ٿ���ѧF�@�����3@�b�~�!?�3�E�^�@l6���ٿ���nJ�@]B8��3@	*����!?�!�~�d�@l6���ٿ���nJ�@]B8��3@	*����!?�!�~�d�@l6���ٿ���nJ�@]B8��3@	*����!?�!�~�d�@�먭�ٿ Oq����@7���3@����я!?BE�T�;�@��n~�ٿ���
���@��$Z� 4@mb�~�!?h' �w�@��n~�ٿ���
���@��$Z� 4@mb�~�!?h' �w�@��n~�ٿ���
���@��$Z� 4@mb�~�!?h' �w�@��n~�ٿ���
���@��$Z� 4@mb�~�!?h' �w�@��n~�ٿ���
���@��$Z� 4@mb�~�!?h' �w�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@G�T(��ٿ��Ёԝ�@:��; 4@���8�!?�Z���x�@_2�]��ٿA�J�L�@����� 4@�'�K̏!?���Fyq�@_2�]��ٿA�J�L�@����� 4@�'�K̏!?���Fyq�@_2�]��ٿA�J�L�@����� 4@�'�K̏!?���Fyq�@2�ۯНٿ�m��e��@"ʘ#�4@��Z�!?ڮ!��@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@v�a���ٿ�VhC���@�57�� 4@���l��!?A�vvΑ�@�F�ٿR�n$��@�E��4@�̫�s�!?��)���@�F�ٿR�n$��@�E��4@�̫�s�!?��)���@�F�ٿR�n$��@�E��4@�̫�s�!?��)���@A.�3�ٿ�CDľ]�@����J 4@IJ���!?hᨨl�@�/3���ٿY���1h�@c���w 4@�l*[�!?��|�o�@�/3���ٿY���1h�@c���w 4@�l*[�!?��|�o�@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@C��1��ٿ��B�c�@Eэ 4@��W6�!?�#P����@b���ٿ��M ��@��� 4@���E�!?-tf����@b���ٿ��M ��@��� 4@���E�!?-tf����@����ٿ9�c��@�F�?�3@�o�&{�!?�g���@����ٿ9�c��@�F�?�3@�o�&{�!?�g���@����ٿ9�c��@�F�?�3@�o�&{�!?�g���@;j�-��ٿ��Q5��@iz�lP�3@��xxp�!?�M�#3�@;j�-��ٿ��Q5��@iz�lP�3@��xxp�!?�M�#3�@8�*�i�ٿ�'v�� �@���~��3@s�HkP�!?��f^�@8�*�i�ٿ�'v�� �@���~��3@s�HkP�!?��f^�@8�*�i�ٿ�'v�� �@���~��3@s�HkP�!?��f^�@���3�ٿ��%���@�X�y��3@H�)��!?r�6e#�@���3�ٿ��%���@�X�y��3@H�)��!?r�6e#�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@Ofwf�ٿ�3�V��@B˕# 4@lˍ_��!?��LY�j�@s�>3i�ٿJ�4`��@�%1�4@CR�I��!?`q=���@s�>3i�ٿJ�4`��@�%1�4@CR�I��!?`q=���@s�>3i�ٿJ�4`��@�%1�4@CR�I��!?`q=���@s�>3i�ٿJ�4`��@�%1�4@CR�I��!?`q=���@���ٿQv�r�@"��4@7��!?Z㣶o��@���ٿQv�r�@"��4@7��!?Z㣶o��@���ٿQv�r�@"��4@7��!?Z㣶o��@7dAEW�ٿ����[X�@=�n�4@��Jϸ�!?�Ug�\�@7dAEW�ٿ����[X�@=�n�4@��Jϸ�!?�Ug�\�@7dAEW�ٿ����[X�@=�n�4@��Jϸ�!?�Ug�\�@7dAEW�ٿ����[X�@=�n�4@��Jϸ�!?�Ug�\�@Q��=΢ٿ/3���@���%� 4@��(:�!?@�W���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@<�
<H�ٿ~�V����@�� 4@2�/��!?�P���@�����ٿ��[���@VeZ/ 4@��Rw�!?�쟮�3�@�����ٿ��[���@VeZ/ 4@��Rw�!?�쟮�3�@v����ٿ�O��@Yu 4@���T��!?$7��_��@v����ٿ�O��@Yu 4@���T��!?$7��_��@v����ٿ�O��@Yu 4@���T��!?$7��_��@v����ٿ�O��@Yu 4@���T��!?$7��_��@v����ٿ�O��@Yu 4@���T��!?$7��_��@m'?�:�ٿ~������@��WR� 4@�y7J͏!?P>n����@�Q���ٿ�tժ��@�E8�� 4@�;�$��!?��H1��@�Q���ٿ�tժ��@�E8�� 4@�;�$��!?��H1��@�Q���ٿ�tժ��@�E8�� 4@�;�$��!?��H1��@�Q���ٿ�tժ��@�E8�� 4@�;�$��!?��H1��@��$��ٿ����@�@qIN���3@hZ���!?`0��/��@��$��ٿ����@�@qIN���3@hZ���!?`0��/��@����ٿ��d;Ĥ�@�ԡP 4@g#��̏!?��[��@����ٿ��d;Ĥ�@�ԡP 4@g#��̏!?��[��@����ٿ��d;Ĥ�@�ԡP 4@g#��̏!?��[��@����ٿ��d;Ĥ�@�ԡP 4@g#��̏!?��[��@����ٿ��d;Ĥ�@�ԡP 4@g#��̏!?��[��@*��b�ٿH�_]v�@ga����3@���� �!?��e����@*��b�ٿH�_]v�@ga����3@���� �!?��e����@*��b�ٿH�_]v�@ga����3@���� �!?��e����@�,Xb�ٿ7o� -��@�8e.�4@�����!?33^�f�@�,Xb�ٿ7o� -��@�8e.�4@�����!?33^�f�@�,Xb�ٿ7o� -��@�8e.�4@�����!?33^�f�@�,Xb�ٿ7o� -��@�8e.�4@�����!?33^�f�@�,Xb�ٿ7o� -��@�8e.�4@�����!?33^�f�@��E�o�ٿ�H\{�@ Ƣ��4@ k �!?�g�#v�@��E�o�ٿ�H\{�@ Ƣ��4@ k �!?�g�#v�@��E�o�ٿ�H\{�@ Ƣ��4@ k �!?�g�#v�@��E�o�ٿ�H\{�@ Ƣ��4@ k �!?�g�#v�@��E�o�ٿ�H\{�@ Ƣ��4@ k �!?�g�#v�@�&N�ٿ�y ����@������3@�����!?����@����Чٿ�o+g�@�0�� 4@"�֥��!?�M�礃�@����Чٿ�o+g�@�0�� 4@"�֥��!?�M�礃�@����Чٿ�o+g�@�0�� 4@"�֥��!?�M�礃�@��Z6�ٿo
���@�`1nU4@�B䩾�!?�ɭ��_�@��Z6�ٿo
���@�`1nU4@�B䩾�!?�ɭ��_�@��Z6�ٿo
���@�`1nU4@�B䩾�!?�ɭ��_�@����ٿ�c�����@`��4@�w]kZ�!?!�`*�@����ٿ�c�����@`��4@�w]kZ�!?!�`*�@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@~�4G�ٿz�%k�@�~�� 4@��b�ˏ!?�[q%��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@I�z�ٿ&H�
���@F�.�}4@�i���!?]2��V��@B��Hӱٿe����@��A�3 4@��
jҏ!?�rk�>R�@B��Hӱٿe����@��A�3 4@��
jҏ!?�rk�>R�@B��Hӱٿe����@��A�3 4@��
jҏ!?�rk�>R�@B��Hӱٿe����@��A�3 4@��
jҏ!?�rk�>R�@a\o��ٿ�e|����@��=e� 4@���=��!?�A��I�@a\o��ٿ�e|����@��=e� 4@���=��!?�A��I�@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@A|M�I�ٿ�2\�s��@Hf�s)4@4��}�!?9��s��@{��
�ٿ�<�^���@�pM4@�a�p��!?�����@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@=�{���ٿE<|� ��@+�{�4@1�0g��!?.mHƬ��@�bFGV�ٿ�V�=��@�e�"�4@���:�!?!��{��@�bFGV�ٿ�V�=��@�e�"�4@���:�!?!��{��@�FNiA�ٿB�]���@c�<8�4@�<�}V�!?��!��[�@.��y�ٿ�u�zu\�@�̠x�4@;ȾDU�!?swR�P��@.��y�ٿ�u�zu\�@�̠x�4@;ȾDU�!?swR�P��@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@l����ٿ��E�|�@,4�9 4@O��y�!?ױ���i�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@)��ٿH	�Tr|�@�?���3@�!<G��!?$� sp,�@T�2�ٿ7�����@I�5� 4@����!?���cK�@8��QΟٿ�X���@�r�&�4@2o�ݏ!?���h]�@8��QΟٿ�X���@�r�&�4@2o�ݏ!?���h]�@8��QΟٿ�X���@�r�&�4@2o�ݏ!?���h]�@8��QΟٿ�X���@�r�&�4@2o�ݏ!?���h]�@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�fFP�ٿL�g���@�7]�4@��ڻӏ!?uId~��@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@�H)īٿ���'9��@+��dk4@-Y�z��!?(��
���@���e4�ٿEhr�!&�@����d4@NvȊ��!?��h'�t�@���e4�ٿEhr�!&�@����d4@NvȊ��!?��h'�t�@���e4�ٿEhr�!&�@����d4@NvȊ��!?��h'�t�@���e4�ٿEhr�!&�@����d4@NvȊ��!?��h'�t�@�Ͳ�C�ٿ7���=Y�@��� 4@qn#��!?��LB���@�Ͳ�C�ٿ7���=Y�@��� 4@qn#��!?��LB���@�Ͳ�C�ٿ7���=Y�@��� 4@qn#��!?��LB���@�Ͳ�C�ٿ7���=Y�@��� 4@qn#��!?��LB���@�Ͳ�C�ٿ7���=Y�@��� 4@qn#��!?��LB���@��
�e�ٿ#$)��@o2}C��3@�푺��!?mן��@��R��ٿ���=�'�@rKֶt4@�;���!?b��i��@��R��ٿ���=�'�@rKֶt4@�;���!?b��i��@��R��ٿ���=�'�@rKֶt4@�;���!?b��i��@��R��ٿ���=�'�@rKֶt4@�;���!?b��i��@���ٿ>�6+�@Blp�;4@�,��!?h�ed��@���ٿ>�6+�@Blp�;4@�,��!?h�ed��@���ٿ>�6+�@Blp�;4@�,��!?h�ed��@���ٿ>�6+�@Blp�;4@�,��!?h�ed��@�[b�ʥٿ��,q�@͡�KW4@
�м�!?M�=JP�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@x�y���ٿ�!����@p"%{��3@B�!)7�!?i���S�@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@gsWg�ٿy�(-ޜ�@���� 4@�3����!?����@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@W�*Ry�ٿY!j@hl�@'�q��4@�Y��!? !da��@��[���ٿ(����@��B4@�:E�y�!?FP�gs��@��[���ٿ(����@��B4@�:E�y�!?FP�gs��@��[���ٿ(����@��B4@�:E�y�!?FP�gs��@�(�A�ٿo�p��.�@#yKW4@�+R-V�!?�k�r-��@�(�A�ٿo�p��.�@#yKW4@�+R-V�!?�k�r-��@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@o
��ٿ��s6�@� �Ph4@]\#�_�!?^EB�FX�@'���ٿ�vDy��@���	�4@��f)��!?�3؏G�@Z��.�ٿ�?���Q�@��{�4@��osT�!?T`����@Z��.�ٿ�?���Q�@��{�4@��osT�!?T`����@�~(嚬ٿY�~#��@.�G�F4@��f�'�!?D�u��@�_��ٿ>kQY��@�uۦ4@!v�Z��!?����x-�@�_��ٿ>kQY��@�uۦ4@!v�Z��!?����x-�@j�v!�ٿ��7�_��@���8�4@r��@��!?�����9�@j�v!�ٿ��7�_��@���8�4@r��@��!?�����9�@/خ<�ٿȑ>�Q8�@%�d�3@��U{v�!?���L�u�@/خ<�ٿȑ>�Q8�@%�d�3@��U{v�!?���L�u�@/خ<�ٿȑ>�Q8�@%�d�3@��U{v�!?���L�u�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@<�)R;�ٿ�����@�,z���3@��cNt�!?��J^]1�@
5=�ğٿ5δ���@
P�m� 4@��z�c�!?��?�UG�@
5=�ğٿ5δ���@
P�m� 4@��z�c�!?��?�UG�@
5=�ğٿ5δ���@
P�m� 4@��z�c�!?��?�UG�@
5=�ğٿ5δ���@
P�m� 4@��z�c�!?��?�UG�@
5=�ğٿ5δ���@
P�m� 4@��z�c�!?��?�UG�@1;6��ٿ[�!����@<�c�s4@��w���!?O	��@�߾{�ٿ�Hń���@s�
�\�3@�Ճ�[�!?4}p^v�@�߾{�ٿ�Hń���@s�
�\�3@�Ճ�[�!?4}p^v�@�/�A��ٿ�T��@�ԏ��3@����w�!?�R��@��@�/�A��ٿ�T��@�ԏ��3@����w�!?�R��@��@�+�p�ٿݫ}}��@���.>�3@�`��_�!?ex����@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@؏��2�ٿ�Ķ���@L+�'�3@z�^+j�!?�B	�n�@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@=H����ٿ�9���@�h��� 4@<��E�!?K`8���@�L���ٿ�+ƺb��@؛��s 4@��rO��!?	#<����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@'9����ٿa$��U�@�}h�� 4@i���!?��W����@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@(w�Ճ�ٿws(����@�_R��4@L
����!?n�6�k�@�yv,o�ٿ���&��@N.R+�4@�o��!?�����X�@�yv,o�ٿ���&��@N.R+�4@�o��!?�����X�@�yv,o�ٿ���&��@N.R+�4@�o��!?�����X�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@ ��卫ٿ#q���@z*���4@(���!?�(D6�\�@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@/a0q�ٿE�s.��@x����4@k��n��!?����@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@��Ê�ٿ1BRw�@����4@F��f��!?�A<{�]�@S$P'�ٿ������@�� z�3@��3]��!?�gm_���@O8e��ٿ6��r���@�pM��3@��U��!?�]E\��@O8e��ٿ6��r���@�pM��3@��U��!?�]E\��@O8e��ٿ6��r���@�pM��3@��U��!?�]E\��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@�BơٿT�kE��@����3@�7Ļ�!?�M�8)��@6�у��ٿ���Z��@�r2�3@������!?c�O)#�@6�у��ٿ���Z��@�r2�3@������!?c�O)#�@゜-�ٿ�NIIGo�@�B` 4@ݿJJ��!?�6 �h�@゜-�ٿ�NIIGo�@�B` 4@ݿJJ��!?�6 �h�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@A���ٿ�����@�Zî� 4@L(�P��!?�5���^�@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@�j�ٿ,eE#�r�@˪k7b 4@�U팏!?dG3#���@��a�,�ٿ5}k�u�@����;�3@�btȋ�!?qd= q�@��a�,�ٿ5}k�u�@����;�3@�btȋ�!?qd= q�@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�!ͫ��ٿ�~.��@lR!n��3@z�b��!?������@�CAN��ٿ�����@�pr\�4@��K��!?��C���@�CAN��ٿ�����@�pr\�4@��K��!?��C���@�CAN��ٿ�����@�pr\�4@��K��!?��C���@�7��Ԩٿx��o��@8C_�4@5���L�!?4I8/���@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@����ٿ0Q_��@�Ĝ 4@B��}�!?������@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@�z U�ٿse�?�@Ah��4@w��R��!?T�ie��@ �g�*�ٿ�G�����@��Po� 4@h,�!?\����@*��*�ٿ�A� �@�
���4@ G�X��!?�X����@*��*�ٿ�A� �@�
���4@ G�X��!?�X����@*��*�ٿ�A� �@�
���4@ G�X��!?�X����@�阚ٿ���@�7G��4@���·�!?H󠄴�@2��7�ٿ���Sx��@K{8� 4@T%�cZ�!?�>n�c�@2��7�ٿ���Sx��@K{8� 4@T%�cZ�!?�>n�c�@2��7�ٿ���Sx��@K{8� 4@T%�cZ�!?�>n�c�@2��7�ٿ���Sx��@K{8� 4@T%�cZ�!?�>n�c�@2��7�ٿ���Sx��@K{8� 4@T%�cZ�!?�>n�c�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@�/2�{�ٿ��x$���@]��<4@{c��ڏ!?P���^�@1��Ţٿ�É�=�@.E�� 4@�Z�Ʉ�!?Ynfc^�@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@x����ٿ6��+��@s}m�d4@8	6N��!?�*���@����ٿK�^����@��[2�4@ ���!?;?QsQ�@pR.-�ٿ�{��@r�/z 4@�
���!?P�:��@pR.-�ٿ�{��@r�/z 4@�
���!?P�:��@pR.-�ٿ�{��@r�/z 4@�
���!?P�:��@�DzܥٿqC�����@���E4@��Vа�!?�oLm��@�DzܥٿqC�����@���E4@��Vа�!?�oLm��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@P�7���ٿ�M���@�h�5P 4@�A��u�!?X4n�y��@��+�I�ٿu�s�^�@ ��� 4@�8T���!?�'��\��@�=�W)�ٿ���O�*�@駓�3@Տ��Ϗ!?O�*���@�=�W)�ٿ���O�*�@駓�3@Տ��Ϗ!?O�*���@t���s�ٿ9K'L��@���y�3@�z�Ə!?�3�z��@Y��f��ٿ��p����@]�t��4@�eP�Ï!?�"B�_�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@u=-$�ٿt"��@�$� 4@S;�ɡ�!?��E��|�@kw=x�ٿ��3kp�@�#��m�3@S����!?�0��]�@kw=x�ٿ��3kp�@�#��m�3@S����!?�0��]�@kw=x�ٿ��3kp�@�#��m�3@S����!?�0��]�@�0��Ġٿ�Կ��@��.�.�3@���۵�!?
��E�@�0��Ġٿ�Կ��@��.�.�3@���۵�!?
��E�@�0��Ġٿ�Կ��@��.�.�3@���۵�!?
��E�@�0��Ġٿ�Կ��@��.�.�3@���۵�!?
��E�@_
��0�ٿ~�G�*l�@�{�\��3@�W���!?�`mƧL�@SJw�ٿ����%��@�J 4@��t��!?�����@SJw�ٿ����%��@�J 4@��t��!?�����@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@���0E�ٿ�#O���@��a� 4@���Y��!?�-q^���@]Ja��ٿ߽�Yt�@����4@���v�!?XC���@]Ja��ٿ߽�Yt�@����4@���v�!?XC���@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@ѻm�ٿ7�7lBX�@��ns 4@@��w�!?k����P�@_��$�ٿT~'�G��@�e3^ 4@:m�ԟ�!?ddF�"�@_��$�ٿT~'�G��@�e3^ 4@:m�ԟ�!?ddF�"�@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@,|���ٿ�;��~�@�`^�E 4@�����!?=�e���@�'r��ٿÅ�N(��@��%��3@�,Q(��!?j�Y0^#�@�'r��ٿÅ�N(��@��%��3@�,Q(��!?j�Y0^#�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@��.RU�ٿ��?�v�@qWlaK�3@J�w���!?�pK�_�@QcU)�ٿ���AOq�@l��Q 4@�\鳏!?�5�����@QcU)�ٿ���AOq�@l��Q 4@�\鳏!?�5�����@QcU)�ٿ���AOq�@l��Q 4@�\鳏!?�5�����@QcU)�ٿ���AOq�@l��Q 4@�\鳏!?�5�����@w���̢ٿ^:��c��@؜�� 4@��ۏ!?P���8��@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@)�?;��ٿ�mBA�X�@6�a� 4@�􏥏!?Ri� �@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@g�~�¬ٿ5�@�}�@��f]� 4@�ȩ.��!??+�j�	�@W�ɹ��ٿ&�C}���@�����4@��;t�!?�Mڣ �@�E��B�ٿ�""S��@D�}r�4@�	���!?���3��@�E��B�ٿ�""S��@D�}r�4@�	���!?���3��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@_��)m�ٿ���s�@�L�q 4@R�T�J�!?/`��2��@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@mћs�ٿrc�Br�@�"P4@�1i�!?�
n�O�@��mhC�ٿ~j)� ��@D�d�s 4@G�`\�!?td����@)`��֯ٿ1IT2,�@!�{�r�3@����\�!?�,]�/��@)`��֯ٿ1IT2,�@!�{�r�3@����\�!?�,]�/��@)`��֯ٿ1IT2,�@!�{�r�3@����\�!?�,]�/��@)`��֯ٿ1IT2,�@!�{�r�3@����\�!?�,]�/��@�(g�V�ٿ�+g�,�@P-�a�3@�|V�y�!?���X���@�(g�V�ٿ�+g�,�@P-�a�3@�|V�y�!?���X���@��TB�ٿ�>y�O�@�����3@'3���!?)q�TE�@��TB�ٿ�>y�O�@�����3@'3���!?)q�TE�@��TB�ٿ�>y�O�@�����3@'3���!?)q�TE�@��TB�ٿ�>y�O�@�����3@'3���!?)q�TE�@Ƣ('[�ٿ��ٶ>��@S�
)u 4@����z�!?.j.���@���`[�ٿq��>�@ꍏA� 4@Hlr���!?R�� ?�@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@ۑ�"-�ٿ�筠�B�@�Z#�3@c>��]�!?�fC�Z��@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@���e�ٿ��,�K�@�0@T� 4@SL��!?���Y���@{*���ٿoT�Z�}�@�( ��3@�~t�!?�D ���@{*���ٿoT�Z�}�@�( ��3@�~t�!?�D ���@{*���ٿoT�Z�}�@�( ��3@�~t�!?�D ���@{*���ٿoT�Z�}�@�( ��3@�~t�!?�D ���@��x�t�ٿ��Q z�@��;?� 4@���Ξ�!?&��1�@��x�t�ٿ��Q z�@��;?� 4@���Ξ�!?&��1�@��x�t�ٿ��Q z�@��;?� 4@���Ξ�!?&��1�@\��q��ٿ!l����@5z��� 4@�A��!?UF�m���@\��q��ٿ!l����@5z��� 4@�A��!?UF�m���@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��0Ԝ�ٿ��
��@���� 4@w��T��!?�bqUˁ�@��9��ٿ $����@o� �4@�C��!?N"\*��@��9��ٿ $����@o� �4@�C��!?N"\*��@��9��ٿ $����@o� �4@�C��!?N"\*��@A���ٿ�Ŋ���@�2��4@p8�Hڏ!?U2o\ �@A���ٿ�Ŋ���@�2��4@p8�Hڏ!?U2o\ �@�|8 ��ٿ����/�@z���4@�P��!?�!���@�|8 ��ٿ����/�@z���4@�P��!?�!���@�|8 ��ٿ����/�@z���4@�P��!?�!���@����ٿh����@���4@��wĻ�!?[��ǋ(�@����ٿh����@���4@��wĻ�!?[��ǋ(�@����ٿh����@���4@��wĻ�!?[��ǋ(�@y��M>�ٿ�}�c���@���4@��ф��!?����@y��M>�ٿ�}�c���@���4@��ф��!?����@y��M>�ٿ�}�c���@���4@��ф��!?����@	 ��K�ٿ�t�W���@eC�.��3@�f)���!?����@	 ��K�ٿ�t�W���@eC�.��3@�f)���!?����@1�r.��ٿLҋ���@EU��H 4@�o3�!?b�AL�g�@1�r.��ٿLҋ���@EU��H 4@�o3�!?b�AL�g�@
��8ȯٿ0�Τ��@�R���3@���ߏ!?��3Ɖ��@W��D��ٿ	U%�`G�@�bXa 4@��؏!?ƚ��D]�@W��D��ٿ	U%�`G�@�bXa 4@��؏!?ƚ��D]�@W��D��ٿ	U%�`G�@�bXa 4@��؏!?ƚ��D]�@Ӵg��ٿ#5�(�K�@�eMo�3@f�P�!?�"�Z,�@���#�ٿ60��cm�@](��4@��3:ɏ!?���+`��@���#�ٿ60��cm�@](��4@��3:ɏ!?���+`��@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�n��X�ٿ����)�@�)�  4@F�����!?�#`�}�@�V����ٿ�,x[+��@�@tfN 4@#u�n��!?ۻp���@�I>t�ٿ�<�"��@�ˑ ��3@��x�!?^F܁��@�I>t�ٿ�<�"��@�ˑ ��3@��x�!?^F܁��@�I>t�ٿ�<�"��@�ˑ ��3@��x�!?^F܁��@�!���ٿ��x���@�HR7� 4@��i�!?�r|�U�@(ZF�ٿðz[��@�F�� 4@}�㼜�!?�ǧ��P�@(ZF�ٿðz[��@�F�� 4@}�㼜�!?�ǧ��P�@(ZF�ٿðz[��@�F�� 4@}�㼜�!?�ǧ��P�@	�z�P�ٿŖ9�Uy�@g��fi4@f"�s`�!?!�`H;�@	�z�P�ٿŖ9�Uy�@g��fi4@f"�s`�!?!�`H;�@}�3���ٿ󑜠"��@d��4@�z{���!?��.�@}�3���ٿ󑜠"��@d��4@�z{���!?��.�@}�3���ٿ󑜠"��@d��4@�z{���!?��.�@}�3���ٿ󑜠"��@d��4@�z{���!?��.�@��k��ٿ,g-%�a�@hU��_4@Y!���!?���g��@��k��ٿ,g-%�a�@hU��_4@Y!���!?���g��@��k��ٿ,g-%�a�@hU��_4@Y!���!?���g��@X�קٿ���F|�@L�8�J4@�KG�A�!?m�N@��@X�קٿ���F|�@L�8�J4@�KG�A�!?m�N@��@X�קٿ���F|�@L�8�J4@�KG�A�!?m�N@��@X�קٿ���F|�@L�8�J4@�KG�A�!?m�N@��@�5���ٿG�j.���@V/�G4@r#""H�!?�W��E�@�5���ٿG�j.���@V/�G4@r#""H�!?�W��E�@�zúz�ٿ�|���@����� 4@"?eft�!?�@b�p�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@!�񂚤ٿ�<]k��@q*@6�4@ax)���!?��c�7�@�ȴE��ٿ}��&G��@�[�4@�f+؏!?T�u����@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�S��O�ٿX�A�/�@5k�#D 4@�@�@*�!?%	���@�%᠊�ٿV���bG�@+U�K 4@���ߏ!?眀?}t�@�%᠊�ٿV���bG�@+U�K 4@���ߏ!?眀?}t�@gZ��ѰٿQ����p�@W�vX4@�9׼��!?���k���@gZ��ѰٿQ����p�@W�vX4@�9׼��!?���k���@pt�"G�ٿz��[�@;���4@�z�n�!?<W�ݲ��@��a҅�ٿ�����@�
+� 4@����!?�d��G�@��a҅�ٿ�����@�
+� 4@����!?�d��G�@�� V[�ٿy>/��L�@��U�4@�r���!?J�I��@'3fX�ٿ���{ah�@��$v<4@#���!?a�ϢZi�@'3fX�ٿ���{ah�@��$v<4@#���!?a�ϢZi�@'3fX�ٿ���{ah�@��$v<4@#���!?a�ϢZi�@'3fX�ٿ���{ah�@��$v<4@#���!?a�ϢZi�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�Tz�U�ٿϭJb� �@�Ғ� 4@���<�!?ǉ�c�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@�&��ٿ��nڲ�@Sz��� 4@đ�E�!?�!�:�g�@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@.?hb2�ٿ����@�?�U4@��
ӏ!?Ts��\��@ꯪ�עٿbx��0�@'��7:4@��W�Ï!?�]�{=��@�rz�!�ٿ��)S��@T��Z 4@����!?7�S����@�rz�!�ٿ��)S��@T��Z 4@����!?7�S����@�rz�!�ٿ��)S��@T��Z 4@����!?7�S����@;V���ٿ��ā�@�a*C 4@�s���!?p
��9�@!���ٿ9������@��.t�3@�p�ߓ�!?YCyv��@!���ٿ9������@��.t�3@�p�ߓ�!?YCyv��@!���ٿ9������@��.t�3@�p�ߓ�!?YCyv��@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@��G��ٿJ���@[�UȬ 4@�|:T|�!?�T����@�"�|�ٿڬ�N�(�@E+��3@w\޽��!?������@�	Dªٿ��_����@��l��3@Ј���!?��eZ��@߳hO~�ٿȏ�/�}�@�e�E� 4@�0Qv�!?��C����@߳hO~�ٿȏ�/�}�@�e�E� 4@�0Qv�!?��C����@߳hO~�ٿȏ�/�}�@�e�E� 4@�0Qv�!?��C����@߳hO~�ٿȏ�/�}�@�e�E� 4@�0Qv�!?��C����@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@bܝ�ٿ��-P�>�@�:d�7 4@ߵ���!?Ip5���@$a�%��ٿ m���-�@��O1��3@�aЏ!?gJgX��@$a�%��ٿ m���-�@��O1��3@�aЏ!?gJgX��@�^L	�ٿ�ֶ x�@�{���3@$�=��!?7�R���@���O�ٿ�n&� ��@0��&5�3@�6`�!?�G�{���@���O�ٿ�n&� ��@0��&5�3@�6`�!?�G�{���@���O�ٿ�n&� ��@0��&5�3@�6`�!?�G�{���@���O�ٿ�n&� ��@0��&5�3@�6`�!?�G�{���@���O�ٿ�n&� ��@0��&5�3@�6`�!?�G�{���@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��!l��ٿ������@���  4@@�,�4�!? �w��a�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@��q��ٿ������@�h+�4@�꣨��!?e蹫SW�@m��ٿ�Y�4��@?�-\4@QVF���!?y[����@ҡ���ٿ�>��@4T�&4@x�s��!?R�A��!�@ҡ���ٿ�>��@4T�&4@x�s��!?R�A��!�@ҡ���ٿ�>��@4T�&4@x�s��!?R�A��!�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@���ٿ!*� ���@�?Ng94@�=2�!?���^-�@.��W�ٿ +3�\"�@��\)4@{�f��!?C��o���@.��W�ٿ +3�\"�@��\)4@{�f��!?C��o���@.��W�ٿ +3�\"�@��\)4@{�f��!?C��o���@�oN��ٿp@�ug��@p��T�4@�F����!?p�{����@$����ٿ��%S	�@`nw,�4@ߡR�ӏ!?���x��@)��ɬٿm"}�,�@D"_�k4@f'tu��!?��k��@י�=��ٿ�h�F�@�⨟�4@�7_���!?#'׼��@�M���ٿ�$��\�@��{��4@�՞���!?r�!�1�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@����~�ٿ�a���u�@����4@���K̏!?r��,�b�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@�dU[�ٿ��0����@�И�y 4@�x�x؏!?]��^x�@���1ȡٿIY�LV�@�ay���3@&d���!?̔Ak��@���1ȡٿIY�LV�@�ay���3@&d���!?̔Ak��@���1ȡٿIY�LV�@�ay���3@&d���!?̔Ak��@t�Z��ٿXkxj�f�@��W	��3@]���!?���&�@t�Z��ٿXkxj�f�@��W	��3@]���!?���&�@t�Z��ٿXkxj�f�@��W	��3@]���!?���&�@t�Z��ٿXkxj�f�@��W	��3@]���!?���&�@t�Z��ٿXkxj�f�@��W	��3@]���!?���&�@�Y0���ٿ;HU����@}k��� 4@{�p�F�!?�T� ��@b��nl�ٿ�cd׎��@;��4@�
L�~�!?�S�y��@b��nl�ٿ�cd׎��@;��4@�
L�~�!?�S�y��@b��nl�ٿ�cd׎��@;��4@�
L�~�!?�S�y��@b��nl�ٿ�cd׎��@;��4@�
L�~�!?�S�y��@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@ѾOm�ٿ9>��JV�@�L��4@���[��!?!�T���@1��a�ٿ�F2ɺD�@��) �4@�I4��!?sAqU���@��5�H�ٿG�ڜ��@O��}�4@ 4h���!?If����@`3	�S�ٿ}���t��@����4@�d}�O�!?��(t<��@`3	�S�ٿ}���t��@����4@�d}�O�!?��(t<��@���*�ٿÔ�E�p�@���� 4@M?�S��!?s�,�@D�ri.�ٿxj�nP��@��K?p�3@�j����!?�=��@D�ri.�ٿxj�nP��@��K?p�3@�j����!?�=��@D�ri.�ٿxj�nP��@��K?p�3@�j����!?�=��@D�ri.�ٿxj�nP��@��K?p�3@�j����!?�=��@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@̊� Θٿܵ=���@�v�s�3@�>��!?^��X�W�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@�&q�ٿK�g�TQ�@*�$���3@�v�n�!?��u�7�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@з�˞ٿ�������@R��s4@+���l�!?��uc�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@Pg#��ٿ_�z�@�ƶ`�4@�#H=�!?�ѡ�Z	�@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@��tZ�ٿ�%EͰ��@y�x�4@3�Lj��!? ;�N���@�fW-��ٿ��غ��@o�К4@$�F�@�!?x~%� �@�fW-��ٿ��غ��@o�К4@$�F�@�!?x~%� �@�fW-��ٿ��غ��@o�К4@$�F�@�!?x~%� �@�fW-��ٿ��غ��@o�К4@$�F�@�!?x~%� �@�fW-��ٿ��غ��@o�К4@$�F�@�!?x~%� �@��~�!�ٿ��S�@��Ҿw�3@�Ed�̏!?���1�@��~�!�ٿ��S�@��Ҿw�3@�Ed�̏!?���1�@Z�)`�ٿ��KX�@�J�I	 4@8�J��!?}V�A�?�@Z�)`�ٿ��KX�@�J�I	 4@8�J��!?}V�A�?�@Z�)`�ٿ��KX�@�J�I	 4@8�J��!?}V�A�?�@Z�)`�ٿ��KX�@�J�I	 4@8�J��!?}V�A�?�@��y�2�ٿ��x�]�@-��|C�3@/U���!?����W��@��y�2�ٿ��x�]�@-��|C�3@/U���!?����W��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@Li��ٿ�g[�|�@�i�ԗ4@�A�l��!?ٱ7:��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@�	�C��ٿ�e�]gJ�@׋�K$4@y����!?�#r�=��@��bY�ٿG?p��1�@轌��4@	0���!?�uF��@��bY�ٿG?p��1�@轌��4@	0���!?�uF��@~S�/��ٿa@A<�@��\�4@N�S�!?���if1�@~S�/��ٿa@A<�@��\�4@N�S�!?���if1�@~S�/��ٿa@A<�@��\�4@N�S�!?���if1�@~S�/��ٿa@A<�@��\�4@N�S�!?���if1�@~S�/��ٿa@A<�@��\�4@N�S�!?���if1�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@s��P�ٿ���K���@���l 4@��Ґ(�!?�h��[�@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@V��`�ٿ+0	����@��P\ 4@�y",��!?�����@R�a�ٿ��H����@�)���3@�T�}�!?�|=eLP�@�:�|x�ٿ/Bݏ|��@���.4@'폠��!?�@�?�b�@�:�|x�ٿ/Bݏ|��@���.4@'폠��!?�@�?�b�@�:�|x�ٿ/Bݏ|��@���.4@'폠��!?�@�?�b�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@s�81�ٿT���T�@h|3/�4@�$�~�!?��=*;)�@[�gol�ٿ��7b�@�b�f4@!�րI�!?�z�F1&�@���C�ٿݨ/m�@��&�X�3@M},XR�!?gV���s�@���C�ٿݨ/m�@��&�X�3@M},XR�!?gV���s�@���C�ٿݨ/m�@��&�X�3@M},XR�!?gV���s�@���C�ٿݨ/m�@��&�X�3@M},XR�!?gV���s�@���C�ٿݨ/m�@��&�X�3@M},XR�!?gV���s�@�'��p�ٿYx�襍�@���h4@���%��!?� ���@�'��p�ٿYx�襍�@���h4@���%��!?� ���@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�W;�ٿ���s���@}�˚Y4@J��i�!?yf`i�@�{i'`�ٿ���l��@��X_4@�j�TÏ!?� �Q���@�{i'`�ٿ���l��@��X_4@�j�TÏ!?� �Q���@�{i'`�ٿ���l��@��X_4@�j�TÏ!?� �Q���@�{i'`�ٿ���l��@��X_4@�j�TÏ!?� �Q���@cF��ٿ�'⚝s�@��k� 4@Q#Cש�!?�K��\��@cF��ٿ�'⚝s�@��k� 4@Q#Cש�!?�K��\��@cF��ٿ�'⚝s�@��k� 4@Q#Cש�!?�K��\��@cF��ٿ�'⚝s�@��k� 4@Q#Cש�!?�K��\��@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@*vJ�l�ٿ��9<�@8�,� 4@�_��ʏ!?�3�+�@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@��E��ٿ��dYM�@U��\� 4@i���!?,�#���@�縋��ٿ:��/p�@�&3�4@!bƴ�!?#��U��@�縋��ٿ:��/p�@�&3�4@!bƴ�!?#��U��@�縋��ٿ:��/p�@�&3�4@!bƴ�!?#��U��@���B��ٿ�	'\���@��i�l4@=�/�!?��2)��@V����ٿT<����@��15A 4@g1���!?������@V����ٿT<����@��15A 4@g1���!?������@V����ٿT<����@��15A 4@g1���!?������@_ri�t�ٿ������@�n����3@<�T��!? y�o��@ޯ�q��ٿ��M�$��@��[� 4@�m()�!?��F<�@ޯ�q��ٿ��M�$��@��[� 4@�m()�!?��F<�@ޯ�q��ٿ��M�$��@��[� 4@�m()�!?��F<�@ޯ�q��ٿ��M�$��@��[� 4@�m()�!?��F<�@��oR�ٿ��V��@'�Ҿ04@+�^��!?c\$�P�@���j�ٿ��'ܷ��@��� �3@�'��z�!?CqȞ�D�@���j�ٿ��'ܷ��@��� �3@�'��z�!?CqȞ�D�@���j�ٿ��'ܷ��@��� �3@�'��z�!?CqȞ�D�@���j�ٿ��'ܷ��@��� �3@�'��z�!?CqȞ�D�@ �v���ٿ��a#��@�(�#@ 4@����!?��.�d��@e�~!��ٿ��;����@�AK�4@b����!?-ZE7H��@e�~!��ٿ��;����@�AK�4@b����!?-ZE7H��@e�~!��ٿ��;����@�AK�4@b����!?-ZE7H��@e�~!��ٿ��;����@�AK�4@b����!?-ZE7H��@e�~!��ٿ��;����@�AK�4@b����!?-ZE7H��@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@���g5�ٿ#�Y���@���4@!�7ԏ!?�� +�S�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�E*w�ٿ�� ����@��'�4@��V讏!?�{���>�@�-Ct)�ٿ��~\���@֕,�4@5>��!?�U�@�-Ct)�ٿ��~\���@֕,�4@5>��!?�U�@�-Ct)�ٿ��~\���@֕,�4@5>��!?�U�@�-Ct)�ٿ��~\���@֕,�4@5>��!?�U�@�
��'�ٿ��B� _�@Y��4@��wG��!?E��io5�@�
��'�ٿ��B� _�@Y��4@��wG��!?E��io5�@d�PZ�ٿVXL7�8�@+sI� 4@������!?��N����@��!��ٿO@M(��@�HN�� 4@_{��!?��23�Y�@��!��ٿO@M(��@�HN�� 4@_{��!?��23�Y�@��!��ٿO@M(��@�HN�� 4@_{��!?��23�Y�@���0�ٿ�K����@��� 4@�R��!?S�Գ{�@�h=!�ٿ꬯�m�@6�T�.4@+n76ŏ!?(�z؛�@�h=!�ٿ꬯�m�@6�T�.4@+n76ŏ!?(�z؛�@�.�+2�ٿ���e�@G� -4@�oڏ!?�f�w���@?6�ٿ�K����@g� 4�4@h<@6��!?+�n����@?6�ٿ�K����@g� 4�4@h<@6��!?+�n����@c?U���ٿ24��J�@�Z��� 4@�U��!?��{�@c?U���ٿ24��J�@�Z��� 4@�U��!?��{�@c?U���ٿ24��J�@�Z��� 4@�U��!?��{�@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�abգٿP�gz!=�@�r��3@t�0�Ǐ!?���Ţ��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@�+�ˢٿ��q�d=�@�I K� 4@��)4g�!?��o�0��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@2��ٿ��_�z��@��6��4@����u�!?�S�o5��@�ⲽf�ٿ�Sa�$1�@��-�Y4@�1��?�!?�����@�ⲽf�ٿ�Sa�$1�@��-�Y4@�1��?�!?�����@�ⲽf�ٿ�Sa�$1�@��-�Y4@�1��?�!?�����@�ⲽf�ٿ�Sa�$1�@��-�Y4@�1��?�!?�����@�ⲽf�ٿ�Sa�$1�@��-�Y4@�1��?�!?�����@�Q�D��ٿD������@x��Q�4@����N�!?#&z���@�Q�D��ٿD������@x��Q�4@����N�!?#&z���@�Q�D��ٿD������@x��Q�4@����N�!?#&z���@�Q�D��ٿD������@x��Q�4@����N�!?#&z���@���1��ٿ7w�����@2�<;��3@%��@��!?]�1���@O��b!�ٿ6�B�))�@����� 4@λ���!?"��W���@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@7	�{$�ٿ4V*��@m�L84@����L�!?5,����@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@��ki�ٿ��k"��@�@kČ 4@�IH?X�!?���7#n�@���r�ٿ�6���@�����3@�|<Y�!?���m��@Ǉ�Z��ٿ:Q&��6�@�QÐ�4@[���!?As�l֜�@Ǉ�Z��ٿ:Q&��6�@�QÐ�4@[���!?As�l֜�@�@X
�ٿ�Y�&N�@)��H�4@)/�!?�B�
��@�@X
�ٿ�Y�&N�@)��H�4@)/�!?�B�
��@s(pQ?�ٿK�tы]�@�T�>4@�5�c��!?K@��F��@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@@��<�ٿ��u��@��c�� 4@��wʏ!??8���@��K�'�ٿ,ʯ�l�@˔�4@��j���!?�{>q�@��K�'�ٿ,ʯ�l�@˔�4@��j���!?�{>q�@��K�'�ٿ,ʯ�l�@˔�4@��j���!?�{>q�@��K�'�ٿ,ʯ�l�@˔�4@��j���!?�{>q�@��K�'�ٿ,ʯ�l�@˔�4@��j���!?�{>q�@ �����ٿo�����@f���q 4@8&�yR�!?fԝ���@ �����ٿo�����@f���q 4@8&�yR�!?fԝ���@����ٿ�X���?�@��G4@hn�%ˏ!?N��Q*Q�@����ٿ�X���?�@��G4@hn�%ˏ!?N��Q*Q�@����ٿ�X���?�@��G4@hn�%ˏ!?N��Q*Q�@����ٿ�X���?�@��G4@hn�%ˏ!?N��Q*Q�@���V�ٿ�%d�[��@�x2�4@��ξ��!?���]�@r��[p�ٿ�
����@6��s� 4@8��_��!?�^�؃�@r��[p�ٿ�
����@6��s� 4@8��_��!?�^�؃�@r��[p�ٿ�
����@6��s� 4@8��_��!?�^�؃�@�aٿڳٿ9Ѐ�.�@�d;^4@ ~��!?<�7
��@D��^�ٿҴ]���@T�,W 4@�)��!?�҂�*�@6��ʬٿS�HF�7�@�@T� 4@j�}�!?�p]R?��@�>�ϫٿ�|jnkJ�@?���� 4@�T9���!?��y�#�@�>�ϫٿ�|jnkJ�@?���� 4@�T9���!?��y�#�@�>�ϫٿ�|jnkJ�@?���� 4@�T9���!?��y�#�@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@��9X��ٿ��ZƓ�@�J(DG4@n����!?&1{{V��@�B�[�ٿv�T)���@a�vz 4@uL��r�!?u�m��<�@�B�[�ٿv�T)���@a�vz 4@uL��r�!?u�m��<�@�B�[�ٿv�T)���@a�vz 4@uL��r�!?u�m��<�@�B�[�ٿv�T)���@a�vz 4@uL��r�!?u�m��<�@�`�?�ٿ�"�`��@7͵h� 4@<Ɛu�!?��B��|�@�`�?�ٿ�"�`��@7͵h� 4@<Ɛu�!?��B��|�@��'���ٿ��Z���@�=�#o 4@��썏!?�j��p`�@��'���ٿ��Z���@�=�#o 4@��썏!?�j��p`�@��'���ٿ��Z���@�=�#o 4@��썏!?�j��p`�@��'���ٿ��Z���@�=�#o 4@��썏!?�j��p`�@�;�r��ٿ��q���@ ��6� 4@����!?���c���@�;�r��ٿ��q���@ ��6� 4@����!?���c���@�;�r��ٿ��q���@ ��6� 4@����!?���c���@��+���ٿw{�	��@���^��3@b����!?ʬFS��@�ĥp�ٿceE�5�@�����3@����S�!?�8�:*�@�ĥp�ٿceE�5�@�����3@����S�!?�8�:*�@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@��!&�ٿ�k�c<�@?�� n�3@�sr�z�!?;���u��@���ٌ�ٿ~퇂9�@dɲG��3@m����!?�h�#��@(��RE�ٿ�Ç���@b��9�4@S��t��!?�>\1P�@(��RE�ٿ�Ç���@b��9�4@S��t��!?�>\1P�@(��RE�ٿ�Ç���@b��9�4@S��t��!?�>\1P�@(��RE�ٿ�Ç���@b��9�4@S��t��!?�>\1P�@(��RE�ٿ�Ç���@b��9�4@S��t��!?�>\1P�@��kad�ٿ������@�8��4@*�Fߏ!?{c�k�l�@��kad�ٿ������@�8��4@*�Fߏ!?{c�k�l�@��kad�ٿ������@�8��4@*�Fߏ!?{c�k�l�@��kad�ٿ������@�8��4@*�Fߏ!?{c�k�l�@�Cdο�ٿd� Va�@�X�4@���Ѽ�!?��!�u�@��=�,�ٿ�����@N�Js4@;��,G�!?�R�#5�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@���]Y�ٿ��-ޗ.�@��� 4@��!?�WV�ص�@�D�1��ٿ�7)l��@L ��3@5Y� Տ!?;��D��@�D�1��ٿ�7)l��@L ��3@5Y� Տ!?;��D��@�D�1��ٿ�7)l��@L ��3@5Y� Տ!?;��D��@�D�1��ٿ�7)l��@L ��3@5Y� Տ!?;��D��@�D�1��ٿ�7)l��@L ��3@5Y� Տ!?;��D��@/��j�ٿ)	>�S��@G���W4@��'�ݏ!?����7��@/��j�ٿ)	>�S��@G���W4@��'�ݏ!?����7��@/��j�ٿ)	>�S��@G���W4@��'�ݏ!?����7��@/��j�ٿ)	>�S��@G���W4@��'�ݏ!?����7��@$m`D��ٿJ �u6�@�X���3@�w^��!?��t��?�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@�6�Y��ٿ>���4��@��Ě� 4@�I��!?Jl`�g�@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@���</�ٿ=�հ#R�@[�{* 4@�3���!?*����@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@�e�/�ٿ�(���@���J�3@[Dlڏ!?h�q�,��@T�<3$�ٿ�Z~	C��@&�ux 4@U�o!?{3'F#��@T�<3$�ٿ�Z~	C��@&�ux 4@U�o!?{3'F#��@sd��ٿ���D�-�@p���3@����ݏ!?�����@{�3�l�ٿ�fΙ�d�@��_,�3@0_v�!? L���@{�3�l�ٿ�fΙ�d�@��_,�3@0_v�!? L���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@� �A�ٿ�]�P)�@�X��3@M�Wc�!?R9�i���@�u,:�ٿ<��F�\�@=��� 4@�E�u.�!?��>W��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@8a�yR�ٿ�.>!G�@��z�� 4@d=�!?=�Le��@���	�ٿ�����@j�� 4@��j�>�!?_W4F��@���	�ٿ�����@j�� 4@��j�>�!?_W4F��@���	�ٿ�����@j�� 4@��j�>�!?_W4F��@�:Ţٿ~��* ��@��Q!� 4@,z9hb�!?��C	@}�@�:Ţٿ~��* ��@��Q!� 4@,z9hb�!?��C	@}�@�:Ţٿ~��* ��@��Q!� 4@,z9hb�!?��C	@}�@�:Ţٿ~��* ��@��Q!� 4@,z9hb�!?��C	@}�@�:Ţٿ~��* ��@��Q!� 4@,z9hb�!?��C	@}�@�[l�ٿ���A��@)��	4@�N���!?uf���@q�9�ٿ-+���@��><� 4@[WC;��!?_�"��|�@q�9�ٿ-+���@��><� 4@[WC;��!?_�"��|�@q�9�ٿ-+���@��><� 4@[WC;��!?_�"��|�@q�9�ٿ-+���@��><� 4@[WC;��!?_�"��|�@�ԫQ�ٿ�d�E�X�@vn�#� 4@�>G}w�!?�|�6�@�ԫQ�ٿ�d�E�X�@vn�#� 4@�>G}w�!?�|�6�@u��{�ٿ۴gΗ%�@QW��w4@Sw~,��!?�[��8�@u��{�ٿ۴gΗ%�@QW��w4@Sw~,��!?�[��8�@u��{�ٿ۴gΗ%�@QW��w4@Sw~,��!?�[��8�@u��{�ٿ۴gΗ%�@QW��w4@Sw~,��!?�[��8�@��0��ٿ|;�O��@�_� 4@R^;��!?ԛ�b��@��0��ٿ|;�O��@�_� 4@R^;��!?ԛ�b��@��0��ٿ|;�O��@�_� 4@R^;��!?ԛ�b��@��0��ٿ|;�O��@�_� 4@R^;��!?ԛ�b��@��k١ٿ\2+���@w�!�C 4@-Á�!?PJs�@��k١ٿ\2+���@w�!�C 4@-Á�!?PJs�@��k١ٿ\2+���@w�!�C 4@-Á�!?PJs�@��k١ٿ\2+���@w�!�C 4@-Á�!?PJs�@��k١ٿ\2+���@w�!�C 4@-Á�!?PJs�@w��
9�ٿ�� ���@q$Idv 4@x�[��!?�tvl�	�@w��
9�ٿ�� ���@q$Idv 4@x�[��!?�tvl�	�@w��
9�ٿ�� ���@q$Idv 4@x�[��!?�tvl�	�@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���+M�ٿvf\8$�@�0��4@N�O�܏!?�k�����@���3��ٿ"��9V��@nKҀ�4@��^���!?U���y��@���3��ٿ"��9V��@nKҀ�4@��^���!?U���y��@���3��ٿ"��9V��@nKҀ�4@��^���!?U���y��@A���ٿ��0�n�@�J0� 4@��fv�!?�+� m�@A���ٿ��0�n�@�J0� 4@��fv�!?�+� m�@A���ٿ��0�n�@�J0� 4@��fv�!?�+� m�@A���ٿ��0�n�@�J0� 4@��fv�!?�+� m�@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@VnD
��ٿ�~. �E�@\Nݩ��3@"sT�`�!?�YM���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@� �,��ٿWzʫ�p�@�"����3@̠�ˏ!?��q���@) !�ʩٿ0���@�^W��3@T}�x�!?������@) !�ʩٿ0���@�^W��3@T}�x�!?������@�pKạٿ��I��@D��: 4@޷�;�!?�oV���@M&��ĥٿH�V��@���Z4@N�Z�I�!?MU���@M&��ĥٿH�V��@���Z4@N�Z�I�!?MU���@M&��ĥٿH�V��@���Z4@N�Z�I�!?MU���@M&��ĥٿH�V��@���Z4@N�Z�I�!?MU���@M&��ĥٿH�V��@���Z4@N�Z�I�!?MU���@$�4�ҭٿ&�+	���@���9�4@y;VM��!?�B,���@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@��e �ٿRdJ,S�@"񗔰�3@�@���!?�濿�_�@|��hקٿM�緙�@��y�� 4@��Q��!?ղAR �@|��hקٿM�緙�@��y�� 4@��Q��!?ղAR �@|��hקٿM�緙�@��y�� 4@��Q��!?ղAR �@|��hקٿM�緙�@��y�� 4@��Q��!?ղAR �@|��hקٿM�緙�@��y�� 4@��Q��!?ղAR �@����r�ٿ>�ќ2�@�_�;% 4@#�●!?v�p>�@����r�ٿ>�ќ2�@�_�;% 4@#�●!?v�p>�@����r�ٿ>�ќ2�@�_�;% 4@#�●!?v�p>�@�W�|��ٿ��9�Y.�@P��
4@=���C�!?����$m�@�W�|��ٿ��9�Y.�@P��
4@=���C�!?����$m�@��`Ϩٿbo��)m�@Q�� 4@��֏!?c�����@��`Ϩٿbo��)m�@Q�� 4@��֏!?c�����@��`Ϩٿbo��)m�@Q�� 4@��֏!?c�����@��`Ϩٿbo��)m�@Q�� 4@��֏!?c�����@��`Ϩٿbo��)m�@Q�� 4@��֏!?c�����@�8%3�ٿ����v�@PA�c�3@q	̏!?EV�G��@�8%3�ٿ����v�@PA�c�3@q	̏!?EV�G��@;�L1�ٿ4�H|��@�J߭O�3@ 콌��!?��K�3�@���j�ٿ\����@���y� 4@<ƥ�!?�	�f�_�@���j�ٿ\����@���y� 4@<ƥ�!?�	�f�_�@���j�ٿ\����@���y� 4@<ƥ�!?�	�f�_�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@|�0��ٿ$i;<���@�F&6�4@�ek��!?5�=�kw�@9�NxH�ٿR; ̘��@�w%es4@>J���!?��G�n�@9�NxH�ٿR; ̘��@�w%es4@>J���!?��G�n�@�V�ٿ�;n��:�@@��~�4@�{0P��!?bLV�M��@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@8��Ĭٿ���b��@+LA�4@'�$��!?�9�j���@0&`�j�ٿJ��s3��@����4@/���[�!?A^��b�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@��{�|�ٿ�Da��@_�(q 4@0�I7Z�!?�JXÕ�@s��fR�ٿhp�a��@ھX�U 4@,�w��!?��F"��@s��fR�ٿhp�a��@ھX�U 4@,�w��!?��F"��@s��fR�ٿhp�a��@ھX�U 4@,�w��!?��F"��@s��fR�ٿhp�a��@ھX�U 4@,�w��!?��F"��@��&Q�ٿ]n5���@��ˀr 4@�p�2�!?�jt�_T�@��&Q�ٿ]n5���@��ˀr 4@�p�2�!?�jt�_T�@��&Q�ٿ]n5���@��ˀr 4@�p�2�!?�jt�_T�@[�.1�ٿ�uo�+J�@�ӂos 4@R�q���!?HWO� 	�@[�.1�ٿ�uo�+J�@�ӂos 4@R�q���!?HWO� 	�@[�.1�ٿ�uo�+J�@�ӂos 4@R�q���!?HWO� 	�@[�.1�ٿ�uo�+J�@�ӂos 4@R�q���!?HWO� 	�@[�.1�ٿ�uo�+J�@�ӂos 4@R�q���!?HWO� 	�@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@#�����ٿs
W9�@S��O�3@W"v���!?7Ͻ�� �@}����ٿ�Z���@��\Ĉ4@�,>6�!?vO/O�@�J	�Ġٿ�4yrFe�@��� 4@���\y�!?9��Q,��@�J	�Ġٿ�4yrFe�@��� 4@���\y�!?9��Q,��@�J	�Ġٿ�4yrFe�@��� 4@���\y�!?9��Q,��@����ٿ�����(�@Έ�M 4@��YcO�!?|�$"�@����ٿ�����(�@Έ�M 4@��YcO�!?|�$"�@����ٿ�����(�@Έ�M 4@��YcO�!?|�$"�@����ٿ�����(�@Έ�M 4@��YcO�!?|�$"�@��LR�ٿ�<c~#�@w�~e�3@�7�M�!?��^�]^�@��LR�ٿ�<c~#�@w�~e�3@�7�M�!?��^�]^�@��LR�ٿ�<c~#�@w�~e�3@�7�M�!?��^�]^�@nbQƝ�ٿ�D*&r�@f�m�4@�y���!?L��wC��@k��&ĥٿ�,x��@(�4@���'��!?6u��-�@k��&ĥٿ�,x��@(�4@���'��!?6u��-�@adV6>�ٿ�r��Ï�@�~a,��3@O��Iݏ!?G����@!�y�Q�ٿ&�y	��@l&�T�3@&�}U��!? �
�@!�y�Q�ٿ&�y	��@l&�T�3@&�}U��!? �
�@�#:�ٿ�������@�tg�3@��㐃�!?����n��@�#:�ٿ�������@�tg�3@��㐃�!?����n��@�#:�ٿ�������@�tg�3@��㐃�!?����n��@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@C�4�ٿ܏ـb�@a����3@��>���!?�_�|�@K��(�ٿG�қ ��@�
t*4@&<���!?���Й}�@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@I��.��ٿ\͡����@�p��4@�|IXȏ!?ⶆ���@�:�|��ٿŃ����@hH9� 4@��q�]�!?��QpA�@�:�|��ٿŃ����@hH9� 4@��q�]�!?��QpA�@{��2��ٿ��߅��@�K<	 4@��p]r�!?W,�+EH�@{��2��ٿ��߅��@�K<	 4@��p]r�!?W,�+EH�@{��2��ٿ��߅��@�K<	 4@��p]r�!?W,�+EH�@{��2��ٿ��߅��@�K<	 4@��p]r�!?W,�+EH�@{��2��ٿ��߅��@�K<	 4@��p]r�!?W,�+EH�@����ٿ���$���@�r�+A 4@�9� ��!?H���l�@����ٿ���$���@�r�+A 4@�9� ��!?H���l�@����ٿ���$���@�r�+A 4@�9� ��!?H���l�@����ٿ���$���@�r�+A 4@�9� ��!?H���l�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@J�/
��ٿ�6�R�@�~����3@���[�!?�W+�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@ߜv��ٿ�����S�@o�өI�3@5��ݏ!?���9�@lʊ�͚ٿ�F>�{��@鸂?��3@����֏!?��|�l��@lʊ�͚ٿ�F>�{��@鸂?��3@����֏!?��|�l��@lʊ�͚ٿ�F>�{��@鸂?��3@����֏!?��|�l��@1;�S�ٿ<����@����3@d�֐�!?�� ��@�Zc6]�ٿX��'�>�@�4���3@��M%n�!?����@
�_U2�ٿ6�\X!��@��YZI�3@�zXZ�!?�AG�x�@s&X��ٿ������@�]Ҵ��3@:ًU^�!?x 7�s��@��UD�ٿ9L��@dB�4@SOo�m�!?�k�%:�@�e΁��ٿ	�'\|�@�C�ʶ�3@S����!?l��-��@�e΁��ٿ	�'\|�@�C�ʶ�3@S����!?l��-��@�e΁��ٿ	�'\|�@�C�ʶ�3@S����!?l��-��@�bx�ٿj���t�@.\��G�3@����w�!?N���@�bx�ٿj���t�@.\��G�3@����w�!?N���@L�r�k�ٿ��Be�z�@����% 4@T	u��!?���?��@L�r�k�ٿ��Be�z�@����% 4@T	u��!?���?��@L�r�k�ٿ��Be�z�@����% 4@T	u��!?���?��@eDEիٿ���|��@c3<_4@�i����!?uLS_�F�@eDEիٿ���|��@c3<_4@�i����!?uLS_�F�@���I�ٿq�2ۛf�@]i3�, 4@�Y$iݏ!?S�� ��@���I�ٿq�2ۛf�@]i3�, 4@�Y$iݏ!?S�� ��@���I�ٿq�2ۛf�@]i3�, 4@�Y$iݏ!?S�� ��@���I�ٿq�2ۛf�@]i3�, 4@�Y$iݏ!?S�� ��@���I�ٿq�2ۛf�@]i3�, 4@�Y$iݏ!?S�� ��@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@��Y�ٿ�y:��@xa�Z� 4@q8>��!?%*��B�@L��c�ٿ�X��@�@I� 
4@XޭЏ!?�v3��@L��c�ٿ�X��@�@I� 
4@XޭЏ!?�v3��@L��c�ٿ�X��@�@I� 
4@XޭЏ!?�v3��@L��c�ٿ�X��@�@I� 
4@XޭЏ!?�v3��@L��c�ٿ�X��@�@I� 
4@XޭЏ!?�v3��@�u�eT�ٿw*�M�A�@� A� 4@O��폏!?��0}�[�@xW�a�ٿ]�q����@| 4@�(҄��!?��J���@xW�a�ٿ]�q����@| 4@�(҄��!?��J���@xW�a�ٿ]�q����@| 4@�(҄��!?��J���@xW�a�ٿ]�q����@| 4@�(҄��!?��J���@xW�a�ٿ]�q����@| 4@�(҄��!?��J���@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@�*Z�U�ٿ�i��@ߘg��3@�w���!?�t8U�p�@X/���ٿz���'�@�ȭ��3@�h�Rŏ!?r�~�@X/���ٿz���'�@�ȭ��3@�h�Rŏ!?r�~�@X/���ٿz���'�@�ȭ��3@�h�Rŏ!?r�~�@�.���ٿ�i��@t{vB��3@Q<���!?��K�@�.���ٿ�i��@t{vB��3@Q<���!?��K�@�.���ٿ�i��@t{vB��3@Q<���!?��K�@�C��ٿ3%#���@ŚJ�< 4@�'��Տ!?1.���5�@�y�$7�ٿ�[�]��@5i�&R4@PE���!?s���J9�@���囜ٿZ��T�g�@�vU�4@+h�Mۏ!?S�
}�~�@���囜ٿZ��T�g�@�vU�4@+h�Mۏ!?S�
}�~�@���囜ٿZ��T�g�@�vU�4@+h�Mۏ!?S�
}�~�@���囜ٿZ��T�g�@�vU�4@+h�Mۏ!?S�
}�~�@���囜ٿZ��T�g�@�vU�4@+h�Mۏ!?S�
}�~�@1)�*��ٿ�,�Lʖ�@����4@Z�'H͏!?��[�;��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@P�$���ٿn�7��@�KشL4@S,)���!?��ç��@h���
�ٿ����~�@<�% 4@qz
�l�!?�/[\�{�@O�\�ٿX@�&G�@���t 4@��5]G�!?��C�%�@O�\�ٿX@�&G�@���t 4@��5]G�!?��C�%�@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@=�9Ý�ٿ^�e�ѻ�@�=7#84@��tV�!?��i��@��2�Ӡٿ�������@d��8� 4@�0f�!?IMi'��@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@�����ٿ��o�@ת�!� 4@(��L��!?́���g�@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@��� ��ٿ�}ar�@�&����3@�14���!?3�*���@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@t� �ٿ���%���@�]�x,4@gC��!?�B���<�@b��{�ٿ�<��1E�@lX�� 4@��Eݞ�!?�b�ܜ*�@b��{�ٿ�<��1E�@lX�� 4@��Eݞ�!?�b�ܜ*�@b��{�ٿ�<��1E�@lX�� 4@��Eݞ�!?�b�ܜ*�@b��{�ٿ�<��1E�@lX�� 4@��Eݞ�!?�b�ܜ*�@b��{�ٿ�<��1E�@lX�� 4@��Eݞ�!?�b�ܜ*�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��+6�ٿۻ'�[�@�e`�4@�auŏ!?���w�@��Q���ٿ�����@}�?84@�W��!?^al�,��@��Q���ٿ�����@}�?84@�W��!?^al�,��@��Q���ٿ�����@}�?84@�W��!?^al�,��@r���ٿ����Q�@��Va� 4@K#����!?Y��b��@r���ٿ����Q�@��Va� 4@K#����!?Y��b��@!U2�ٿų��#��@�<0U4@��协!?�;8��H�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@�p��ٿ����c��@\S0W� 4@'�r~��!?�ǩ�@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@ ���ٿ�ȬAs��@�2�v$4@�x�-o�!?�.ң��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@�D(�ٿ��*[L�@�d���3@������!?_N}�@��@w,����ٿ����@��Åw 4@��ҏ!?k.���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@X��¥ٿ !�0�D�@K�	4 4@@hӏ!?���@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@q���Q�ٿ�gJ.[�@Լ[]��3@�TW̏!?��,�@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@����ٿ�Z��7N�@֙�UB 4@�tQ�ӏ!?�������@�K�]�ٿ4:�b���@��5+� 4@�֩��!?���a$��@V�CՑ�ٿW�u�@���`)�3@X��U�!?htTT�2�@V�CՑ�ٿW�u�@���`)�3@X��U�!?htTT�2�@S�_�W�ٿh�]�d��@�	=��3@&"r�!?-wP�e��@Y�L�ٿ��(�D��@�u�k6 4@���9�!?�>���@Y�L�ٿ��(�D��@�u�k6 4@���9�!?�>���@Y�L�ٿ��(�D��@�u�k6 4@���9�!?�>���@��0F�ٿ��l�K�@�I�^. 4@[�8���!?2��E��@��4E�ٿ�\"��@���� 4@.�fqf�!?��R	��@��\�צٿ�y�ܶ�@�!� 4@��:���!?�7�����@��\�צٿ�y�ܶ�@�!� 4@��:���!?�7�����@��\�צٿ�y�ܶ�@�!� 4@��:���!?�7�����@���(8�ٿ����G}�@дy�4@YJ���!?�)�`��@���(8�ٿ����G}�@дy�4@YJ���!?�)�`��@���(8�ٿ����G}�@дy�4@YJ���!?�)�`��@��Y���ٿ oزg�@:%�k 4@�5;��!?�[����@��Y���ٿ oزg�@:%�k 4@�5;��!?�[����@��Y���ٿ oزg�@:%�k 4@�5;��!?�[����@��Y���ٿ oزg�@:%�k 4@�5;��!?�[����@h�mc�ٿY�w ��@냦� 4@�wC���!?�K^�+�@h�mc�ٿY�w ��@냦� 4@�wC���!?�K^�+�@h�mc�ٿY�w ��@냦� 4@�wC���!?�K^�+�@h�mc�ٿY�w ��@냦� 4@�wC���!?�K^�+�@h�mc�ٿY�w ��@냦� 4@�wC���!?�K^�+�@���%�ٿW�%)o��@��D�F 4@�ܰ�!?��Z��@���%�ٿW�%)o��@��D�F 4@�ܰ�!?��Z��@���%�ٿW�%)o��@��D�F 4@�ܰ�!?��Z��@��zed�ٿ���@� 4@��s|��!?K��v���@��zed�ٿ���@� 4@��s|��!?K��v���@��zed�ٿ���@� 4@��s|��!?K��v���@��zed�ٿ���@� 4@��s|��!?K��v���@��zed�ٿ���@� 4@��s|��!?K��v���@��8dg�ٿ����'��@���|4@ ���̏!?��X���@��8dg�ٿ����'��@���|4@ ���̏!?��X���@�\'�/�ٿu�š��@C�!�$4@�Di��!?\����-�@�\'�/�ٿu�š��@C�!�$4@�Di��!?\����-�@E�*S��ٿ5�����@���%4@�2�ҝ�!?���A&�@�ׄ��ٿ�#����@�߮)c 4@اf���!?O��p��@�ׄ��ٿ�#����@�߮)c 4@اf���!?O��p��@`Ҷ�ٿt�%�@��b{4@��qҏ!?��t�!�@`Ҷ�ٿt�%�@��b{4@��qҏ!?��t�!�@`Ҷ�ٿt�%�@��b{4@��qҏ!?��t�!�@`Ҷ�ٿt�%�@��b{4@��qҏ!?��t�!�@Y�b�ٿ�N�ǜ	�@ʐ�b14@V?��!?�V	ӵ��@�ʔvx�ٿ���
��@����3 4@�8Y�!?����@�<�.#�ٿb�0U��@��T\ 4@�>,�ʏ!?������@�<�.#�ٿb�0U��@��T\ 4@�>,�ʏ!?������@Ck-ڣٿ��*��@6)���3@^�#�ɏ!?��m���@Ck-ڣٿ��*��@6)���3@^�#�ɏ!?��m���@��B��ٿF��b]�@���?I 4@��в�!?�]2�s:�@��B��ٿF��b]�@���?I 4@��в�!?�]2�s:�@��B��ٿF��b]�@���?I 4@��в�!?�]2�s:�@N��ٿ{/���N�@�B^� 4@�pr���!?>�3�n��@k�bs�ٿ�m_�7�@��ȾG�3@���1��!?X������@k�bs�ٿ�m_�7�@��ȾG�3@���1��!?X������@k�bs�ٿ�m_�7�@��ȾG�3@���1��!?X������@k�bs�ٿ�m_�7�@��ȾG�3@���1��!?X������@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@"�hi��ٿצ�o�@�ۤ�3@9���B�!?M��O6�@��=�ٿY�W���@MU^W4@�W��S�!?Uf�fy�@��=�ٿY�W���@MU^W4@�W��S�!?Uf�fy�@��=�ٿY�W���@MU^W4@�W��S�!?Uf�fy�@���<j�ٿ�.��6L�@�
�َ4@9�� `�!?�4�,�R�@���<j�ٿ�.��6L�@�
�َ4@9�� `�!?�4�,�R�@�V[\Z�ٿr�&�>�@���f�4@/sg�=�!?�:x��x�@�V[\Z�ٿr�&�>�@���f�4@/sg�=�!?�:x��x�@�V[\Z�ٿr�&�>�@���f�4@/sg�=�!?�:x��x�@��A-�ٿk�ɹpi�@�>��4@<��g�!?@'��A��@��A-�ٿk�ɹpi�@�>��4@<��g�!?@'��A��@��A-�ٿk�ɹpi�@�>��4@<��g�!?@'��A��@��D���ٿWL^��@�38�D4@͂�|�!?��ED@�@{�[U��ٿ�6&x0=�@ju�4@{OG�w�!?DՁJ��@{�[U��ٿ�6&x0=�@ju�4@{OG�w�!?DՁJ��@rğ�ٿ@��4S�@����4@�_S���!?�î���@rğ�ٿ@��4S�@����4@�_S���!?�î���@ЋX���ٿ�ܡp��@��4@�̩:��!?�vz��@�ޗ�i�ٿ���Z��@U��� 4@�QЭ�!?�k�id��@�cS���ٿ�6(Nn	�@~��#l�3@�W��!?�Khv���@�cS���ٿ�6(Nn	�@~��#l�3@�W��!?�Khv���@=d���ٿ�w�?K�@��U��3@t-���!?����|�@p��9C�ٿ�����@1���4@��c���!?;g��\�@p��9C�ٿ�����@1���4@��c���!?;g��\�@p��9C�ٿ�����@1���4@��c���!?;g��\�@�p*Ò�ٿ�J���@&
� 4@D�q� �!?�b#�8�@�p*Ò�ٿ�J���@&
� 4@D�q� �!?�b#�8�@�uu�ٿ�v4�%r�@>�5�� 4@�h+�+�!?�����@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@�"i)͘ٿ�f���@@G}�) 4@�ک���!?s��@��u�ٿ����v�@�_:� �3@�^��!?��ꙵf�@��u�ٿ����v�@�_:� �3@�^��!?��ꙵf�@��k���ٿ|�p /�@�y>p�3@[m:�q�!?kEN*���@j$){y�ٿa*Lԙ�@\e��7�3@;F�V/�!?'�wd�u�@j$){y�ٿa*Lԙ�@\e��7�3@;F�V/�!?'�wd�u�@�6r�:�ٿ�'r+��@8 P�-�3@���ZA�!?� *���@�6r�:�ٿ�'r+��@8 P�-�3@���ZA�!?� *���@�6r�:�ٿ�'r+��@8 P�-�3@���ZA�!?� *���@�6r�:�ٿ�'r+��@8 P�-�3@���ZA�!?� *���@�6r�:�ٿ�'r+��@8 P�-�3@���ZA�!?� *���@w&�酚ٿZl���H�@��:�	4@�,��J�!?荽T�@w&�酚ٿZl���H�@��:�	4@�,��J�!?荽T�@��͙�ٿ/!�{�@���� 4@nr����!?��ۗ&��@�E��h�ٿܻ3����@+��Q 4@8��g�!?�|LU1.�@�C��V�ٿ(�9��2�@"i'�� 4@��J-|�!?�"�a=g�@�C��V�ٿ(�9��2�@"i'�� 4@��J-|�!?�"�a=g�@�C��V�ٿ(�9��2�@"i'�� 4@��J-|�!?�"�a=g�@�C��V�ٿ(�9��2�@"i'�� 4@��J-|�!?�"�a=g�@FV���ٿ��m�S�@�n�n�3@�J����!?���-�@FV���ٿ��m�S�@�n�n�3@�J����!?���-�@���ٿ$$�}a�@�����3@��J���!?*����@�@�KF�ٿ2�T3���@�к��3@���ӏ!?����3v�@�~��ٿ�4����@jq�� 4@��[�!?�1\���@�~��ٿ�4����@jq�� 4@��[�!?�1\���@�'�j��ٿ����@x� �4@���!?V0�J���@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@X���E�ٿ�Ē���@�|]��4@w��{܏!?�y��w�@(e��6�ٿtv/�Q�@���z?4@f����!?ğ>r;�@(e��6�ٿtv/�Q�@���z?4@f����!?ğ>r;�@,�(�ٿd�ͨ���@6�Lޟ4@5�
�!?��9��@,�(�ٿd�ͨ���@6�Lޟ4@5�
�!?��9��@(���ٿybn���@��w�� 4@N՗ ��!?���d�1�@N"@�S�ٿ.bq�� �@�f�#� 4@�hԂZ�!?>�/�pG�@N"@�S�ٿ.bq�� �@�f�#� 4@�hԂZ�!?>�/�pG�@N"@�S�ٿ.bq�� �@�f�#� 4@�hԂZ�!?>�/�pG�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@znh��ٿ�#�'��@j#�d`�3@־=��!?�ZX�X�@/�Mͨٿ��f�B��@%%%o�4@p��d�!?��+9̳�@/�Mͨٿ��f�B��@%%%o�4@p��d�!?��+9̳�@/�Mͨٿ��f�B��@%%%o�4@p��d�!?��+9̳�@��P9�ٿ]7`�:
�@&m68 4@o�W���!?y��ʥ-�@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@s	�@�ٿ-oUnP��@D�`q4@kW^��!?Y���E��@�]��'�ٿxR��2��@C��o4@;���!?e�����@�]��'�ٿxR��2��@C��o4@;���!?e�����@�]��'�ٿxR��2��@C��o4@;���!?e�����@Lt`EB�ٿ����]"�@Тd��4@����ď!?Y�S���@Lt`EB�ٿ����]"�@Тd��4@����ď!?Y�S���@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@�HW+�ٿo�誔��@���0� 4@�r3�ԏ!?W� ��@.�+�ٿF�����@�����3@����!?@��=���@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ)�����@:3���3@�t���!?*����z�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@����ٿ���M?�@�)�x 4@��#\��!?�0��+�@E�}�b�ٿ����S�@$�?54@�=���!?�3D*�@E�}�b�ٿ����S�@$�?54@�=���!?�3D*�@E�}�b�ٿ����S�@$�?54@�=���!?�3D*�@E�}�b�ٿ����S�@$�?54@�=���!?�3D*�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@��#ݨٿ�C5��z�@F*P�(4@	�Gr~�!?��*ź�@����ٿCE����@���4@� KL�!?+��Q;k�@����ٿCE����@���4@� KL�!?+��Q;k�@����ٿCE����@���4@� KL�!?+��Q;k�@����ٿCE����@���4@� KL�!?+��Q;k�@����ٿCE����@���4@� KL�!?+��Q;k�@C��hG�ٿy�i�+��@V��ef4@�拏!?*���Z�@C��hG�ٿy�i�+��@V��ef4@�拏!?*���Z�@C��hG�ٿy�i�+��@V��ef4@�拏!?*���Z�@C��hG�ٿy�i�+��@V��ef4@�拏!?*���Z�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@zE}��ٿJ�ki���@ ���S4@J8�Bj�!?,���y�@�%+̩ٿQ3%���@����4@���ُ!?�}���@�%+̩ٿQ3%���@����4@���ُ!?�}���@�%+̩ٿQ3%���@����4@���ُ!?�}���@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@�Q�j%�ٿ+Y��~��@0s�94@�myw�!?�R����@=�Ey�ٿmt�#t�@;0����3@��꘏!?�	^�@=�Ey�ٿmt�#t�@;0����3@��꘏!?�	^�@=�Ey�ٿmt�#t�@;0����3@��꘏!?�	^�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@�Ɋ�ٿ��ν���@����3@A���ˏ!?
��{�4�@����,�ٿ��	{�@��uV� 4@�x��!?�ꝑ��@����,�ٿ��	{�@��uV� 4@�x��!?�ꝑ��@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@���ٿ���T��@�HJ4@~z��!?`�����@�@#��ٿ�=��(}�@G0��� 4@OeI�!?�n��w	�@�@#��ٿ�=��(}�@G0��� 4@OeI�!?�n��w	�@�@#��ٿ�=��(}�@G0��� 4@OeI�!?�n��w	�@$XX_��ٿ����@�UC��3@m #k�!?,&����@$XX_��ٿ����@�UC��3@m #k�!?,&����@k�sɬٿ�+g=�@�v�|54@�1\_��!?����g��@k�sɬٿ�+g=�@�v�|54@�1\_��!?����g��@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@F`n�y�ٿ��BtH��@�K�4@d~綏!?N�����@[�a�1�ٿ�[�f��@�W$�4@�m�u�!?����w�@[�a�1�ٿ�[�f��@�W$�4@�m�u�!?����w�@[�a�1�ٿ�[�f��@�W$�4@�m�u�!?����w�@[�a�1�ٿ�[�f��@�W$�4@�m�u�!?����w�@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@cy��X�ٿ0^�]���@"�yk��3@Y���!?��7�[��@�'@�ٿu���\�@P��F��3@�PY{�!?PN��*��@U��3�ٿA�(�'�@B �f��3@m��R�!?��<x_�@�Ȟ_��ٿlD6m?|�@$n9Η�3@�N_���!?�w�� �@��f�}�ٿ��!�;��@�0�q�4@8�
�!?"�B���@��f�}�ٿ��!�;��@�0�q�4@8�
�!?"�B���@��f�}�ٿ��!�;��@�0�q�4@8�
�!?"�B���@m9��ˤٿ��ˁ�@ք�� 4@mZ��!?,L,q.�@m9��ˤٿ��ˁ�@ք�� 4@mZ��!?,L,q.�@m9��ˤٿ��ˁ�@ք�� 4@mZ��!?,L,q.�@]�Q�ٿ]�_����@~��8�4@����!?|�b���@]�Q�ٿ]�_����@~��8�4@����!?|�b���@gB����ٿ/�@����@ ��0 4@���!?h��!$�@��6�ٿd�(I�+�@H��"4@�<C���!?�G$A��@��6�ٿd�(I�+�@H��"4@�<C���!?�G$A��@�e&Κٿ�מ�Y��@<�����3@DQd'��!?K��d�@�e&Κٿ�מ�Y��@<�����3@DQd'��!?K��d�@�e&Κٿ�מ�Y��@<�����3@DQd'��!?K��d�@�e&Κٿ�מ�Y��@<�����3@DQd'��!?K��d�@��&B��ٿ�20Lm��@֓����3@l��Ս�!?j�j���@��&B��ٿ�20Lm��@֓����3@l��Ս�!?j�j���@��&B��ٿ�20Lm��@֓����3@l��Ս�!?j�j���@�ཌ��ٿ8 g^���@���E�3@��c��!?k%˞�B�@�ཌ��ٿ8 g^���@���E�3@��c��!?k%˞�B�@�ཌ��ٿ8 g^���@���E�3@��c��!?k%˞�B�@�ཌ��ٿ8 g^���@���E�3@��c��!?k%˞�B�@�ཌ��ٿ8 g^���@���E�3@��c��!?k%˞�B�@�𝧕ٿE�K��@6Bt� 4@���C��!?��t���@�𝧕ٿE�K��@6Bt� 4@���C��!?��t���@�𝧕ٿE�K��@6Bt� 4@���C��!?��t���@�𝧕ٿE�K��@6Bt� 4@���C��!?��t���@�ȕ�ٿ��6��@ɘ���4@Vv�x�!?n�L	�D�@�ȕ�ٿ��6��@ɘ���4@Vv�x�!?n�L	�D�@��a��ٿOi�:��@��@� 4@� �;��!?�d���@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@?H�ll�ٿ��$�3��@�`L�e�3@��s/��!?8����g�@��k��ٿG����@��#[P�3@�߅7�!?I4䀌-�@��k��ٿG����@��#[P�3@�߅7�!?I4䀌-�@��k��ٿG����@��#[P�3@�߅7�!?I4䀌-�@���H�ٿ�YNf�@�)��3@��٣ݏ!?�+���@���H�ٿ�YNf�@�)��3@��٣ݏ!?�+���@AH���ٿGu��@@�Y@4@3��O�!?��s�d�@AH���ٿGu��@@�Y@4@3��O�!?��s�d�@AH���ٿGu��@@�Y@4@3��O�!?��s�d�@�}���ٿ�G��@��@n����3@f�y��!?���Q�@�}���ٿ�G��@��@n����3@f�y��!?���Q�@�}���ٿ�G��@��@n����3@f�y��!?���Q�@�}���ٿ�G��@��@n����3@f�y��!?���Q�@��i�1�ٿ�E�Ƽ�@�H����3@��f|��!?[��/�@��i�1�ٿ�E�Ƽ�@�H����3@��f|��!?[��/�@��i�1�ٿ�E�Ƽ�@�H����3@��f|��!?[��/�@S'��U�ٿ������@�pA�4@Bu�G�!?斐wjY�@S'��U�ٿ������@�pA�4@Bu�G�!?斐wjY�@S'��U�ٿ������@�pA�4@Bu�G�!?斐wjY�@NU��Ģٿ�����@g[H�4@���ٮ�!?��η�6�@�jf�ٿ؇�b�@(��Sy4@��K)*�!?��.?u-�@욛q6�ٿ�كE4"�@��X 4@� ��R�!?�ō
��@욛q6�ٿ�كE4"�@��X 4@� ��R�!?�ō
��@"U ��ٿ��Ni��@��Tg�3@kw#�!?R�1�p`�@"U ��ٿ��Ni��@��Tg�3@kw#�!?R�1�p`�@"U ��ٿ��Ni��@��Tg�3@kw#�!?R�1�p`�@"U ��ٿ��Ni��@��Tg�3@kw#�!?R�1�p`�@"U ��ٿ��Ni��@��Tg�3@kw#�!?R�1�p`�@%�s�ٿ��>��@Qi�2�3@"婂"�!?�z�RE�@%�s�ٿ��>��@Qi�2�3@"婂"�!?�z�RE�@%�s�ٿ��>��@Qi�2�3@"婂"�!?�z�RE�@%�s�ٿ��>��@Qi�2�3@"婂"�!?�z�RE�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@��!�ٿT�����@��*d� 4@�\)��!?�9ڶZF�@�fT/�ٿ^�ޘU�@� ��3@�r鵏!?�����%�@�fT/�ٿ^�ޘU�@� ��3@�r鵏!?�����%�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@�]ʰٿ��YY=��@��� 4@�
ņ��!?'
��6e�@��s0�ٿ�l�6���@���=} 4@I�0��!?����T,�@��s0�ٿ�l�6���@���=} 4@I�0��!?����T,�@��s0�ٿ�l�6���@���=} 4@I�0��!?����T,�@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@�%��ٿ����"��@�uKƨ 4@�=6uY�!?�Wnc/��@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@`���s�ٿ���h�@��a��4@�kkCW�!?c��WU[�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@��tf�ٿv�R/���@ʚ^�\ 4@��y�!?�X��.�@�[�R��ٿ�k����@�a|�4@4�)�{�!?���k��@jo�ٿ�k_���@"�q�4@6�a�3�!?el��*�@jo�ٿ�k_���@"�q�4@6�a�3�!?el��*�@jo�ٿ�k_���@"�q�4@6�a�3�!?el��*�@jo�ٿ�k_���@"�q�4@6�a�3�!?el��*�@jo�ٿ�k_���@"�q�4@6�a�3�!?el��*�@��j.�ٿ�<��f��@I"&4@W����!?�䂫5��@��j.�ٿ�<��f��@I"&4@W����!?�䂫5��@��j.�ٿ�<��f��@I"&4@W����!?�䂫5��@��j.�ٿ�<��f��@I"&4@W����!?�䂫5��@��j.�ٿ�<��f��@I"&4@W����!?�䂫5��@����ٿ?2+�@��Xz��3@x�$�!?���U�<�@����ٿ?2+�@��Xz��3@x�$�!?���U�<�@�bi�ٿ�;t���@�w�w 4@�?2��!?��"�Ȃ�@�bi�ٿ�;t���@�w�w 4@�?2��!?��"�Ȃ�@�bi�ٿ�;t���@�w�w 4@�?2��!?��"�Ȃ�@�bi�ٿ�;t���@�w�w 4@�?2��!?��"�Ȃ�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@�]u��ٿ�=Ki)��@ÜKw�4@L�^��!?��m�L�@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@^�~�ٿ�/�x�w�@��"�� 4@<��Ώ!?A6����@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@�#�?��ٿw�4��t�@�^��� 4@c�V\�!??�/f��@T�{&�ٿ�8C����@�S��j4@��e��!?3�ɤ�{�@T�{&�ٿ�8C����@�S��j4@��e��!?3�ɤ�{�@Z�âٿ�A'�z�@9�� 4@������!?���T,\�@Z�âٿ�A'�z�@9�� 4@������!?���T,\�@Z�âٿ�A'�z�@9�� 4@������!?���T,\�@Z�âٿ�A'�z�@9�� 4@������!?���T,\�@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@hU�i��ٿ�l�4B�@�@�4 4@+�����!?J�y���@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@IޞԟٿI8z��@ �wR( 4@�"k�!?'��R��@� /2ҥٿ8ߏ�h��@a���3@�[l
��!?��J8�@� /2ҥٿ8ߏ�h��@a���3@�[l
��!?��J8�@� /2ҥٿ8ߏ�h��@a���3@�[l
��!?��J8�@� /2ҥٿ8ߏ�h��@a���3@�[l
��!?��J8�@MP����ٿ4�m�ݪ�@h��C��3@?A�!?�0*��{�@MP����ٿ4�m�ݪ�@h��C��3@?A�!?�0*��{�@MP����ٿ4�m�ݪ�@h��C��3@?A�!?�0*��{�@MP����ٿ4�m�ݪ�@h��C��3@?A�!?�0*��{�@MP����ٿ4�m�ݪ�@h��C��3@?A�!?�0*��{�@�Q�[�ٿo����z�@�<� 4@���c��!?k<�?���@�Q�[�ٿo����z�@�<� 4@���c��!?k<�?���@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@���ٿ��ـ���@ 2� 4@��alv�!?,.ף:��@�!=�#�ٿ����v|�@�D��q 4@%`���!?�A�]f��@�!=�#�ٿ����v|�@�D��q 4@%`���!?�A�]f��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@;b*��ٿ��*�T��@;��I4@]s��h�!?�T;FC��@�b�`��ٿC�����@�5�Q4@oO?��!?�w����@�b�`��ٿC�����@�5�Q4@oO?��!?�w����@�b�`��ٿC�����@�5�Q4@oO?��!?�w����@�b�`��ٿC�����@�5�Q4@oO?��!?�w����@Cb� �ٿ!)��9��@��CM4@����K�!?��q]��@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@y��Rܣٿiٹ����@i
۵ 4@����b�!?h����@�%a�0�ٿOפ3o�@4m�]p 4@ᯋ�ȏ!?�6w�L.�@�%a�0�ٿOפ3o�@4m�]p 4@ᯋ�ȏ!?�6w�L.�@�%a�0�ٿOפ3o�@4m�]p 4@ᯋ�ȏ!?�6w�L.�@�%a�0�ٿOפ3o�@4m�]p 4@ᯋ�ȏ!?�6w�L.�@�%a�0�ٿOפ3o�@4m�]p 4@ᯋ�ȏ!?�6w�L.�@�Q�)��ٿN2r��B�@d	FX�3@@�n��!?6eto#��@�Q�)��ٿN2r��B�@d	FX�3@@�n��!?6eto#��@���i�ٿzݻ's��@�"�y 4@�>��n�!?U��!Q�@���i�ٿzݻ's��@�"�y 4@�>��n�!?U��!Q�@���i�ٿzݻ's��@�"�y 4@�>��n�!?U��!Q�@���i�ٿzݻ's��@�"�y 4@�>��n�!?U��!Q�@���i�ٿzݻ's��@�"�y 4@�>��n�!?U��!Q�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@9�=�ٿ7;�n.b�@��v4@��� ��!?��L0�@ѻ}�ٿv��,��@j�5l�4@�a����!?�ŭ+�@ѻ}�ٿv��,��@j�5l�4@�a����!?�ŭ+�@ѻ}�ٿv��,��@j�5l�4@�a����!?�ŭ+�@ѻ}�ٿv��,��@j�5l�4@�a����!?�ŭ+�@����l�ٿ������@�%�+4@o��T�!?����'�@����l�ٿ������@�%�+4@o��T�!?����'�@����l�ٿ������@�%�+4@o��T�!?����'�@����l�ٿ������@�%�+4@o��T�!?����'�@����l�ٿ������@�%�+4@o��T�!?����'�@����l�ٿ������@�%�+4@o��T�!?����'�@QȲ�ٿ�FZC��@���4@LN'͏!?zZ�nU��@QȲ�ٿ�FZC��@���4@LN'͏!?zZ�nU��@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�rbȫٿ������@�Im4@�/Hԏ!?��6i�@�^����ٿm�h����@�2̱4@=����!?�>�I���@�^����ٿm�h����@�2̱4@=����!?�>�I���@�^����ٿm�h����@�2̱4@=����!?�>�I���@��59��ٿRq�<&��@�u=,�4@
)���!?�We�V��@��59��ٿRq�<&��@�u=,�4@
)���!?�We�V��@��59��ٿRq�<&��@�u=,�4@
)���!?�We�V��@��59��ٿRq�<&��@�u=,�4@
)���!?�We�V��@��59��ٿRq�<&��@�u=,�4@
)���!?�We�V��@�f�:H�ٿ]�\���@���#/4@?��x�!?97��~��@�f�:H�ٿ]�\���@���#/4@?��x�!?97��~��@�an�)�ٿký����@	�hv4@J{%ď!??�rJ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@�E��\�ٿ7���l��@�l��Z4@�h�Ѯ�!?Iw�ҭ�@���P�ٿ�2Np���@��j4@j�ieď!?���a��@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@����ٿ:@U�f�@HILi�3@9�v��!?�G�����@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@T3,�{�ٿW&|�C;�@*�I���3@�x�J��!?F�+ɀ�@&0Z�x�ٿ������@6�� 4@�0�s��!?�[�����@&0Z�x�ٿ������@6�� 4@�0�s��!?�[�����@&0Z�x�ٿ������@6�� 4@�0�s��!?�[�����@&0Z�x�ٿ������@6�� 4@�0�s��!?�[�����@�&>˥ٿ�`7���@4L�0y 4@O0���!?�R�Y��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�%2�ٿ�I�l��@h��~ 4@��_�u�!?�cH�{��@�#vsϚٿ��8����@�P��r 4@R��؜�!?sOjm�v�@�#vsϚٿ��8����@�P��r 4@R��؜�!?sOjm�v�@�#vsϚٿ��8����@�P��r 4@R��؜�!?sOjm�v�@��w��ٿ0m�����@#�}4@v�r��!?Y�Y2�@��w��ٿ0m�����@#�}4@v�r��!?Y�Y2�@��w��ٿ0m�����@#�}4@v�r��!?Y�Y2�@��w��ٿ0m�����@#�}4@v�r��!?Y�Y2�@'G�f�ٿ&��Z���@�e�� 4@�׸��!?`�&`e�@'G�f�ٿ&��Z���@�e�� 4@�׸��!?`�&`e�@'G�f�ٿ&��Z���@�e�� 4@�׸��!?`�&`e�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@�'�O�ٿ�����4�@����Y 4@a=d��!?�����x�@��{ëٿ���6��@.B27� 4@�!F�l�!?r��=�@��{ëٿ���6��@.B27� 4@�!F�l�!?r��=�@��{ëٿ���6��@.B27� 4@�!F�l�!?r��=�@��{ëٿ���6��@.B27� 4@�!F�l�!?r��=�@*�H��ٿ[�]TK�@��D�� 4@��<p�!?~ND�v�@*�H��ٿ[�]TK�@��D�� 4@��<p�!?~ND�v�@/�Ѱ�ٿ0�v���@2c� 4@m�oΗ�!?>5D;��@/�Ѱ�ٿ0�v���@2c� 4@m�oΗ�!?>5D;��@/�Ѱ�ٿ0�v���@2c� 4@m�oΗ�!?>5D;��@/�Ѱ�ٿ0�v���@2c� 4@m�oΗ�!?>5D;��@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@9��3�ٿ?i�Zz��@rRo� 4@t)[��!?�J�r���@>��O�ٿmI�����@��c�4@� z���!?}i��u�@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�4{&Q�ٿ��vc��@`�'�64@�T��!?I�:"���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@�A}�ٿ�`�W��@�t~4@�XɆ��!?��k)���@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@$W*$�ٿ�7!^���@"&��S4@���!?���ߢ�@��>���ٿ��06��@�e��4@ENݒ&�!?��1� �@��>���ٿ��06��@�e��4@ENݒ&�!?��1� �@��>���ٿ��06��@�e��4@ENݒ&�!?��1� �@��>���ٿ��06��@�e��4@ENݒ&�!?��1� �@��>���ٿ��06��@�e��4@ENݒ&�!?��1� �@5s\汩ٿB���ң�@0C�%4@�q���!?|��[��@o��z�ٿ���*�4�@:/5���3@!�%`�!?��m����@o��z�ٿ���*�4�@:/5���3@!�%`�!?��m����@��~Ù�ٿ�6A0�G�@k��� 4@�g;��!?ݔ���@��m�ٿR� �d��@����4@t܏!?�!ju���@��m�ٿR� �d��@����4@t܏!?�!ju���@��m�ٿR� �d��@����4@t܏!?�!ju���@��m�ٿR� �d��@����4@t܏!?�!ju���@��m�ٿR� �d��@����4@t܏!?�!ju���@R�մ�ٿ�߉Wq��@u���4@�(��Ϗ!?����1�@R�մ�ٿ�߉Wq��@u���4@�(��Ϗ!?����1�@R�մ�ٿ�߉Wq��@u���4@�(��Ϗ!?����1�@R�մ�ٿ�߉Wq��@u���4@�(��Ϗ!?����1�@�f�B{�ٿ�2���@\jb5k4@c����!?��W��@�f�B{�ٿ�2���@\jb5k4@c����!?��W��@�f�B{�ٿ�2���@\jb5k4@c����!?��W��@�f�B{�ٿ�2���@\jb5k4@c����!?��W��@�f�B{�ٿ�2���@\jb5k4@c����!?��W��@2�f�ٿ`-����@0�6�� 4@��M�ӏ!?�� �T�@2�f�ٿ`-����@0�6�� 4@��M�ӏ!?�� �T�@��Ԑ�ٿ\Zo|�@�үw� 4@B���܏!?�Qo���@��Ԑ�ٿ\Zo|�@�үw� 4@B���܏!?�Qo���@��:��ٿ�r�T��@����4@����!?���O۸�@��:��ٿ�r�T��@����4@����!?���O۸�@��:��ٿ�r�T��@����4@����!?���O۸�@)P���ٿ@U`���@ )Vz04@���8�!?��H�]�@)P���ٿ@U`���@ )Vz04@���8�!?��H�]�@m=�F�ٿ���:��@_�?A� 4@o X�!?������@m=�F�ٿ���:��@_�?A� 4@o X�!?������@`���ٿ��Y����@oUd�� 4@@l���!?]9��V �@`���ٿ��Y����@oUd�� 4@@l���!?]9��V �@T�<��ٿ��t���@$Ձ�g4@b|�`��!?q\�rI�@T�<��ٿ��t���@$Ձ�g4@b|�`��!?q\�rI�@T�<��ٿ��t���@$Ձ�g4@b|�`��!?q\�rI�@T�<��ٿ��t���@$Ձ�g4@b|�`��!?q\�rI�@�e��ٿ��kR���@��R"� 4@�@�,�!?�%����@.�Լ��ٿc8�x\�@�q7jP4@�ۆ�!?˾�T�@.�Լ��ٿc8�x\�@�q7jP4@�ۆ�!?˾�T�@.�Լ��ٿc8�x\�@�q7jP4@�ۆ�!?˾�T�@R�j�q�ٿ��*D0H�@zޒ(74@,W��я!?�������@R�j�q�ٿ��*D0H�@zޒ(74@,W��я!?�������@R�j�q�ٿ��*D0H�@zޒ(74@,W��я!?�������@R�j�q�ٿ��*D0H�@zޒ(74@,W��я!?�������@� G���ٿ�n�g�=�@
��4@/@G��!?�\��@)`�H�ٿ����}`�@|��4@�,�Y�!?�-!fj�@��)ӦٿH=��O��@�Sۖ�4@�;�dD�!?�V��"��@��)ӦٿH=��O��@�Sۖ�4@�;�dD�!?�V��"��@��)ӦٿH=��O��@�Sۖ�4@�;�dD�!?�V��"��@��)ӦٿH=��O��@�Sۖ�4@�;�dD�!?�V��"��@��)ӦٿH=��O��@�Sۖ�4@�;�dD�!?�V��"��@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@7w/K�ٿ�d�3���@����4@������!?7[q	?-�@�a2p�ٿ������@ˏW��4@9���!?��@��@�a2p�ٿ������@ˏW��4@9���!?��@��@�a2p�ٿ������@ˏW��4@9���!?��@��@�a2p�ٿ������@ˏW��4@9���!?��@��@�a2p�ٿ������@ˏW��4@9���!?��@��@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@(b?�\�ٿx�3p���@����� 4@����ُ!?�/��P�@c_\p��ٿw�a�S��@^�0��4@��mĵ�!?��=��@c_\p��ٿw�a�S��@^�0��4@��mĵ�!?��=��@c_\p��ٿw�a�S��@^�0��4@��mĵ�!?��=��@c_\p��ٿw�a�S��@^�0��4@��mĵ�!?��=��@�U����ٿ�QĘ��@*�ߟ4@�y+2�!?^s�b�@�U����ٿ�QĘ��@*�ߟ4@�y+2�!?^s�b�@�U����ٿ�QĘ��@*�ߟ4@�y+2�!?^s�b�@SS�X֤ٿ��H0���@rP4�( 4@t19�[�!?����:x�@�n�ݦٿte��@h�T��4@'G�z��!?�t�%��@�n�ݦٿte��@h�T��4@'G�z��!?�t�%��@�n�ݦٿte��@h�T��4@'G�z��!?�t�%��@Qz��ٿ����@Ds��4@��s��!?��e��@Qz��ٿ����@Ds��4@��s��!?��e��@Qz��ٿ����@Ds��4@��s��!?��e��@��z��ٿ.}����@H�|�^ 4@����F�!?��!P��@��z��ٿ.}����@H�|�^ 4@����F�!?��!P��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@BSњٿ�
�m��@oh%��3@��ܲ��!?�24LR��@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@�QI,�ٿ������@�ݮj��3@.qj���!?[�S��]�@s�'&R�ٿ�=���@�h�3��3@51Q�p�!?��j���@s�'&R�ٿ�=���@�h�3��3@51Q�p�!?��j���@s�'&R�ٿ�=���@�h�3��3@51Q�p�!?��j���@s�'&R�ٿ�=���@�h�3��3@51Q�p�!?��j���@s�'&R�ٿ�=���@�h�3��3@51Q�p�!?��j���@-+�ާٿu�ڗ�@�C�4@$}(�D�!?/�����@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@i,#\�ٿa�.�f�@:�b���3@g6�Y�!?�������@n�!�{�ٿ8P�<�Z�@R�e�A 4@��=~�!?���5�@�m�ٿ_���@�)@��4@�FaҤ�!?�J�/0�@�m�ٿ_���@�)@��4@�FaҤ�!?�J�/0�@�m�ٿ_���@�)@��4@�FaҤ�!?�J�/0�@�m�ٿ_���@�)@��4@�FaҤ�!?�J�/0�@�m�ٿ_���@�)@��4@�FaҤ�!?�J�/0�@�5&�ٿ������@��q4@)����!?�^��@�5&�ٿ������@��q4@)����!?�^��@�5&�ٿ������@��q4@)����!?�^��@�5&�ٿ������@��q4@)����!?�^��@�5&�ٿ������@��q4@)����!?�^��@3���ٿYs�?���@܄M��3@�+L�Y�!?��p��U�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�5<J�ٿ�偬�x�@�\	`��3@�ܼS��!?;�K�r�@�*ү�ٿ��@�R�@���e� 4@�F���!?��Ȭxk�@�*ү�ٿ��@�R�@���e� 4@�F���!?��Ȭxk�@�*ү�ٿ��@�R�@���e� 4@�F���!?��Ȭxk�@�*ү�ٿ��@�R�@���e� 4@�F���!?��Ȭxk�@�*ү�ٿ��@�R�@���e� 4@�F���!?��Ȭxk�@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@tk' ۝ٿ�༰YC�@��{4@��j���!?��L����@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@����9�ٿ��S$���@��r�H4@bikø�!? �D��`�@�!ü��ٿF�?��@�E4@�J��!?4X���@�B-=�ٿ�}�����@7z:(14@�D���!?O�?3���@�B-=�ٿ�}�����@7z:(14@�D���!?O�?3���@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@��.B*�ٿ+�	z��@~��q� 4@��.o��!?J�|L�@g �%g�ٿ�t��mr�@<m+4@#�_��!?܇�jF�@g �%g�ٿ�t��mr�@<m+4@#�_��!?܇�jF�@8��]�ٿ����{�@�mp� 4@�;rn�!?��,�)M�@8��]�ٿ����{�@�mp� 4@�;rn�!?��,�)M�@8��]�ٿ����{�@�mp� 4@�;rn�!?��,�)M�@8��]�ٿ����{�@�mp� 4@�;rn�!?��,�)M�@�ϊ�x�ٿ�J�w�@W�b4@{�m���!?�C�˟�@�ϊ�x�ٿ�J�w�@W�b4@{�m���!?�C�˟�@�ϊ�x�ٿ�J�w�@W�b4@{�m���!?�C�˟�@�ϊ�x�ٿ�J�w�@W�b4@{�m���!?�C�˟�@4o��ٿ@�!A���@]�wf^ 4@��֏!?�o&Q�U�@4o��ٿ@�!A���@]�wf^ 4@��֏!?�o&Q�U�@FP幂�ٿ��?0>��@L�l�U�3@���Џ!?O�U��H�@FP幂�ٿ��?0>��@L�l�U�3@���Џ!?O�U��H�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@��0��ٿ��ԋ��@�s 4@�����!?רr4x�@t�Fk�ٿ���Ѕ�@�Y��a�3@�ƇI��!?3#tO��@t�Fk�ٿ���Ѕ�@�Y��a�3@�ƇI��!?3#tO��@t�Fk�ٿ���Ѕ�@�Y��a�3@�ƇI��!?3#tO��@t�Fk�ٿ���Ѕ�@�Y��a�3@�ƇI��!?3#tO��@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@_B���ٿt�����@������3@MC�%��!?c���t�@��؅C�ٿ��U���@�� 4@�����!?j���@��؅C�ٿ��U���@�� 4@�����!?j���@ ԥC�ٿ�br
a��@S��Z� 4@�;7���!?B_>����@ ԥC�ٿ�br
a��@S��Z� 4@�;7���!?B_>����@ ԥC�ٿ�br
a��@S��Z� 4@�;7���!?B_>����@+ci��ٿE�W���@~��
�4@{J��ԏ!?�0���@+ci��ٿE�W���@~��
�4@{J��ԏ!?�0���@+ci��ٿE�W���@~��
�4@{J��ԏ!?�0���@+ci��ٿE�W���@~��
�4@{J��ԏ!?�0���@+ci��ٿE�W���@~��
�4@{J��ԏ!?�0���@�؄9u�ٿD�XL5u�@���4@���ѯ�!?�qל��@��5zr�ٿ��l^��@`�L�i4@Ҳ���!?5��8�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@n6N$�ٿ��4���@�X�q4@@hq���!?ة�b0�@^�v;�ٿҹk���@>�t�^4@�&pf�!?��]���@^�v;�ٿҹk���@>�t�^4@�&pf�!?��]���@^�v;�ٿҹk���@>�t�^4@�&pf�!?��]���@^�v;�ٿҹk���@>�t�^4@�&pf�!?��]���@^�v;�ٿҹk���@>�t�^4@�&pf�!?��]���@����ٿ!7�$��@���$4@�y�㡏!?��K���@-oq+�ٿ_� O	��@a~��54@D��zǏ!?�q6I�q�@l�y,�ٿ�_q[�~�@��'�4@2����!?k����=�@l�y,�ٿ�_q[�~�@��'�4@2����!?k����=�@l�y,�ٿ�_q[�~�@��'�4@2����!?k����=�@wf��c�ٿO�_���@����4@T1v��!?� �����@wf��c�ٿO�_���@����4@T1v��!?� �����@wf��c�ٿO�_���@����4@T1v��!?� �����@+:]��ٿ�l�z-��@��|�64@���!?��Z}T:�@+:]��ٿ�l�z-��@��|�64@���!?��Z}T:�@+:]��ٿ�l�z-��@��|�64@���!?��Z}T:�@+:]��ٿ�l�z-��@��|�64@���!?��Z}T:�@+:]��ٿ�l�z-��@��|�64@���!?��Z}T:�@
L~��ٿ�T�w+�@n$�e4@w ���!?������@
L~��ٿ�T�w+�@n$�e4@w ���!?������@
L~��ٿ�T�w+�@n$�e4@w ���!?������@
L~��ٿ�T�w+�@n$�e4@w ���!?������@
L~��ٿ�T�w+�@n$�e4@w ���!?������@m蠜ٿڍ�׳��@���Y 4@=�wp��!?�J���@��Cs١ٿ�p�^K��@��O��4@�D�dȏ!?�nq��@�򯩐�ٿW�h ���@�i��/4@xAT�|�!?�l�Hc�@�򯩐�ٿW�h ���@�i��/4@xAT�|�!?�l�Hc�@��C���ٿx������@��5��4@�Es�h�!?��
˵�@��b@��ٿ[�����@��%P�4@����:�!?�����@��b@��ٿ[�����@��%P�4@����:�!?�����@���aџٿ���d6��@ę8�4@d9dˏ!?��+R�@���aџٿ���d6��@ę8�4@d9dˏ!?��+R�@���aџٿ���d6��@ę8�4@d9dˏ!?��+R�@���aџٿ���d6��@ę8�4@d9dˏ!?��+R�@��:rĝٿ��R&4��@�W� 4@ˈ{��!?ZI��8�@��:rĝٿ��R&4��@�W� 4@ˈ{��!?ZI��8�@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@,��:/�ٿh�j�A��@>�]x4@
t箏�!?/74��@Y�����ٿd0Pnq�@.p]? 4@F 2�̏!?�'�>]*�@Y�����ٿd0Pnq�@.p]? 4@F 2�̏!?�'�>]*�@Y�����ٿd0Pnq�@.p]? 4@F 2�̏!?�'�>]*�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@�钋ϡٿǘ��Ń�@֏��� 4@w|�?��!?E	��($�@4�/�ٿ� /�	�@WH��3@s<6�!? ���U�@=����ٿx�� �@�uv�R�3@�S�!?.�e*p�@=����ٿx�� �@�uv�R�3@�S�!?.�e*p�@=����ٿx�� �@�uv�R�3@�S�!?.�e*p�@=����ٿx�� �@�uv�R�3@�S�!?.�e*p�@=����ٿx�� �@�uv�R�3@�S�!?.�e*p�@HR:,�ٿ+4~�-�@%�w4�3@f(I�+�!?�����@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@�k���ٿ%�����@��Z/) 4@M���!?����y�@.��b�ٿ}❩P��@���W4@�a�zh�!?@$��2��@.��b�ٿ}❩P��@���W4@�a�zh�!?@$��2��@.��b�ٿ}❩P��@���W4@�a�zh�!?@$��2��@.��b�ٿ}❩P��@���W4@�a�zh�!?@$��2��@.��b�ٿ}❩P��@���W4@�a�zh�!?@$��2��@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@G�5q�ٿL)�U���@��~I4@���eO�!?���Gܰ�@��dq�ٿ�k8��\�@�{��O�3@�q�F�!?r�i���@��dq�ٿ�k8��\�@�{��O�3@�q�F�!?r�i���@��dq�ٿ�k8��\�@�{��O�3@�q�F�!?r�i���@���ХٿS�.O�@P��� 4@RCҝY�!?ڡ��U�@���ХٿS�.O�@P��� 4@RCҝY�!?ڡ��U�@���ХٿS�.O�@P��� 4@RCҝY�!?ڡ��U�@^�d�ٿ�͙��F�@4�\�� 4@�W����!?��5��=�@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@k��`�ٿYvZd0�@��� 4@���}֏!?�����@Rڽ2��ٿ������@F�{,4@]�`z��!?ۀ�$���@Rڽ2��ٿ������@F�{,4@]�`z��!?ۀ�$���@Rڽ2��ٿ������@F�{,4@]�`z��!?ۀ�$���@Rڽ2��ٿ������@F�{,4@]�`z��!?ۀ�$���@��G��ٿ�fVS+��@ȍ/���3@����!?-��Z�@��G��ٿ�fVS+��@ȍ/���3@����!?-��Z�@��G��ٿ�fVS+��@ȍ/���3@����!?-��Z�@4O�l�ٿ �$z�@3���H4@t��Q��!?e��*A�@4O�l�ٿ �$z�@3���H4@t��Q��!?e��*A�@�q���ٿ�Y���@֋<�y4@������!?%�T&:�@G%��ٿ��TU_��@\"��f�3@�,j�p�!?�\�2>�@G%��ٿ��TU_��@\"��f�3@�,j�p�!?�\�2>�@G%��ٿ��TU_��@\"��f�3@�,j�p�!?�\�2>�@G%��ٿ��TU_��@\"��f�3@�,j�p�!?�\�2>�@G%��ٿ��TU_��@\"��f�3@�,j�p�!?�\�2>�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@�j���ٿ�{�l�@�ӄX)4@�&����!?�J��ڝ�@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@S�!r�ٿ|4�j��@b�9!� 4@�TO���!?��3!���@+Dq/�ٿ�}��&x�@�\�,� 4@�c��!? ���7��@+Dq/�ٿ�}��&x�@�\�,� 4@�c��!? ���7��@+Dq/�ٿ�}��&x�@�\�,� 4@�c��!? ���7��@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@�2�T�ٿ��/����@�nJ�4@W���!?(6��<�@m��9��ٿ��A����@���<�4@~Ru��!?���s���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@"d����ٿ�S��f��@��(W4@(`�V��!?�y���@�/1�r�ٿ	�|��@D��4@�1�p��!?ǒ�����@�/1�r�ٿ	�|��@D��4@�1�p��!?ǒ�����@�/1�r�ٿ	�|��@D��4@�1�p��!?ǒ�����@v�K��ٿ)���R��@��n�4@)���~�!?��/bn��@v�K��ٿ)���R��@��n�4@)���~�!?��/bn��@v�K��ٿ)���R��@��n�4@)���~�!?��/bn��@v�K��ٿ)���R��@��n�4@)���~�!?��/bn��@v�K��ٿ)���R��@��n�4@)���~�!?��/bn��@#��s�ٿf
E���@��5�4@Lp�}�!?[�Qw�@#��s�ٿf
E���@��5�4@Lp�}�!?[�Qw�@#��s�ٿf
E���@��5�4@Lp�}�!?[�Qw�@#��s�ٿf
E���@��5�4@Lp�}�!?[�Qw�@�[	ɰ�ٿ3g;J���@�w���3@��u�!?�&�L�2�@�[	ɰ�ٿ3g;J���@�w���3@��u�!?�&�L�2�@�[	ɰ�ٿ3g;J���@�w���3@��u�!?�&�L�2�@�[	ɰ�ٿ3g;J���@�w���3@��u�!?�&�L�2�@�[	ɰ�ٿ3g;J���@�w���3@��u�!?�&�L�2�@��r@��ٿ�>��G��@lٌ^��3@>+��p�!?ݝȅ���@��r@��ٿ�>��G��@lٌ^��3@>+��p�!?ݝȅ���@J����ٿ�{m�@磃�!4@X��@��!?)��T��@J����ٿ�{m�@磃�!4@X��@��!?)��T��@�\N�ٿ��cdg�@��9�; 4@t�����!?U�3����@�\N�ٿ��cdg�@��9�; 4@t�����!?U�3����@d��J��ٿS����@��
i 4@O�ܬ�!?8�4p�E�@d��J��ٿS����@��
i 4@O�ܬ�!?8�4p�E�@d��J��ٿS����@��
i 4@O�ܬ�!?8�4p�E�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@�L�ՠٿG��8��@� �4@�]ք̏!?NY�Ĳ�@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@v!�ٿO���k�@p_R�3@5��ݧ�!?�s�l���@�6�ٿ7���@SG ���3@x��f�!?X���%��@�6�ٿ7���@SG ���3@x��f�!?X���%��@�6�ٿ7���@SG ���3@x��f�!?X���%��@�6�ٿ7���@SG ���3@x��f�!?X���%��@�6�ٿ7���@SG ���3@x��f�!?X���%��@ч�AG�ٿ]?�1n��@�y��4@��� �!?!޸�<\�@ч�AG�ٿ]?�1n��@�y��4@��� �!?!޸�<\�@,4Cd�ٿ�U�C��@ǧڋJ4@3U���!?5�.�%�@,4Cd�ٿ�U�C��@ǧڋJ4@3U���!?5�.�%�@)�Y�J�ٿ������@�"�	%4@"i6Ï!?�oTA��@�`�V�ٿ�/"���@n�BL�4@p�+���!?	�O����@��&y�ٿl u1	v�@p!� 4@fJ��X�!?�#z͍�@��&y�ٿl u1	v�@p!� 4@fJ��X�!?�#z͍�@��&y�ٿl u1	v�@p!� 4@fJ��X�!?�#z͍�@łO��ٿ��O����@<�S��4@u�w�J�!?�:����@łO��ٿ��O����@<�S��4@u�w�J�!?�:����@łO��ٿ��O����@<�S��4@u�w�J�!?�:����@łO��ٿ��O����@<�S��4@u�w�J�!?�:����@łO��ٿ��O����@<�S��4@u�w�J�!?�:����@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@G>�hx�ٿ�I0�vX�@��{+ 4@5ܢ���!?�<��V�@j��
��ٿ�;:���@����04@{�&��!?��+F�@��ŧ�ٿ�q�����@3źO 4@��s֏!?��9t�@6^��ٿ��.k��@�G��} 4@�N���!?�27%w��@6^��ٿ��.k��@�G��} 4@�N���!?�27%w��@6^��ٿ��.k��@�G��} 4@�N���!?�27%w��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@���ky�ٿ��,����@���(� 4@�<�vR�!?��ٓ��@7,S/�ٿ��^���@i��С�3@:�%O�!?{𩢝z�@7,S/�ٿ��^���@i��С�3@:�%O�!?{𩢝z�@7,S/�ٿ��^���@i��С�3@:�%O�!?{𩢝z�@7,S/�ٿ��^���@i��С�3@:�%O�!?{𩢝z�@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@W��J��ٿY��}g��@gH���3@�:�M�!?e9�1��@q/�V�ٿ�M/�J�@������3@��;��!?��ǯ��@q/�V�ٿ�M/�J�@������3@��;��!?��ǯ��@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@�5�zS�ٿ��~�t�@AD�o��3@�t(2Ώ!?8��ּ�@-�# �ٿa��'.��@aB�ER�3@,ю�e�!?�Y�@�@-�# �ٿa��'.��@aB�ER�3@,ю�e�!?�Y�@�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@&+�/�ٿhN?�z�@ {:lw�3@�?�*_�!?\�>Hܘ�@��tçٿ��J�v��@}�;��3@�J��z�!?� �C>[�@��tçٿ��J�v��@}�;��3@�J��z�!?� �C>[�@�B����ٿ(b�?9�@�T����3@Y�X��!?��8�8�@��9N��ٿie����@�{�0;�3@m�4nS�!?��U�,��@��9N��ٿie����@�{�0;�3@m�4nS�!?��U�,��@��9N��ٿie����@�{�0;�3@m�4nS�!?��U�,��@}Fb֜ٿ��Z�@�0�3@h1s�v�!?��ċN�@}Fb֜ٿ��Z�@�0�3@h1s�v�!?��ċN�@}Fb֜ٿ��Z�@�0�3@h1s�v�!?��ċN�@}Fb֜ٿ��Z�@�0�3@h1s�v�!?��ċN�@}Fb֜ٿ��Z�@�0�3@h1s�v�!?��ċN�@z+XV��ٿ�wJm�@o���3@��O��!?�W4[��@z+XV��ٿ�wJm�@o���3@��O��!?�W4[��@i����ٿh�͔�Z�@>�]�3@�H��!?ÿ�>Y��@i����ٿh�͔�Z�@>�]�3@�H��!?ÿ�>Y��@�'�R�ٿ �U�.{�@T�M��3@�=�!?Rl���@�'�R�ٿ �U�.{�@T�M��3@�=�!?Rl���@k<�e�ٿ�qϙ�I�@�����3@ts�!?M!fPA�@k<�e�ٿ�qϙ�I�@�����3@ts�!?M!fPA�@k<�e�ٿ�qϙ�I�@�����3@ts�!?M!fPA�@k<�e�ٿ�qϙ�I�@�����3@ts�!?M!fPA�@k<�e�ٿ�qϙ�I�@�����3@ts�!?M!fPA�@���r��ٿ*VtV`��@�}���3@6]��4�!?D�6���@C�r�έٿͲ&O��@L��k�3@.��o׏!?��
o�@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@��|6��ٿѶ�]���@�rY�+ 4@d�C�!?n��ޏ��@�I�?m�ٿ�/m����@�Ѝ��3@�i���!?R�h_��@�I�?m�ٿ�/m����@�Ѝ��3@�i���!?R�h_��@R�yKk�ٿ��)���@���\U 4@�(t���!?-�⤺�@R�yKk�ٿ��)���@���\U 4@�(t���!?-�⤺�@R�yKk�ٿ��)���@���\U 4@�(t���!?-�⤺�@���H�ٿg�IM��@�H����3@M�dY>�!?A�~�<�@���܍�ٿK.�D|h�@�l
���3@�U����!?vn�1��@���܍�ٿK.�D|h�@�l
���3@�U����!?vn�1��@���܍�ٿK.�D|h�@�l
���3@�U����!?vn�1��@���܍�ٿK.�D|h�@�l
���3@�U����!?vn�1��@z�Z5v�ٿh
�����@=�����3@��W��!?���W �@ҩe�ٿ�3����@�����3@�V�)؏!?�.�MH �@ҩe�ٿ�3����@�����3@�V�)؏!?�.�MH �@K rݢٿ	5c_��@�d�)4@�YƏ!?�EY���@��"u0�ٿ#�?I���@����u�3@���R��!?m{Oc��@jn�H�ٿ�r���N�@��Ҵ6�3@G�mv�!?6;��;��@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@\����ٿ���m=��@�NtT4@A�����!?�#ItO�@�G�ٿN�M��@Ǯ��� 4@�@r�!?N �=S�@�G�ٿN�M��@Ǯ��� 4@�@r�!?N �=S�@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�"���ٿW�&�a@�@AV|[~ 4@g�=xe�!?��y�B��@�\Ģ�ٿ!���G��@���4@��%�W�!?�x��v2�@�\Ģ�ٿ!���G��@���4@��%�W�!?�x��v2�@%�E�M�ٿ�`@8v�@h1�4@o��]�!?\A�1G<�@��ϳ�ٿ��o:��@
8�Y4@/8�&z�!?�`���@��ϳ�ٿ��o:��@
8�Y4@/8�&z�!?�`���@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@���+n�ٿIU����@:�]k� 4@�c�`ԏ!?�����@��a�ЭٿL������@h���3@<ڡΏ!?Xb�%=�@��a�ЭٿL������@h���3@<ڡΏ!?Xb�%=�@	�
��ٿK@���@�jt4<�3@v�aߏ!?�ҁ(��@	�
��ٿK@���@�jt4<�3@v�aߏ!?�ҁ(��@	�
��ٿK@���@�jt4<�3@v�aߏ!?�ҁ(��@	�
��ٿK@���@�jt4<�3@v�aߏ!?�ҁ(��@��I��ٿ�-RW�t�@��^��3@������!?��`��@Fk���ٿ�?�NW��@�I�_4 4@�yp�!?lV�U���@Fk���ٿ�?�NW��@�I�_4 4@�yp�!?lV�U���@Fk���ٿ�?�NW��@�I�_4 4@�yp�!?lV�U���@Fk���ٿ�?�NW��@�I�_4 4@�yp�!?lV�U���@Fk���ٿ�?�NW��@�I�_4 4@�yp�!?lV�U���@VN�灧ٿ��7��&�@K-�]Y 4@:?P�ď!?��hr���@VN�灧ٿ��7��&�@K-�]Y 4@:?P�ď!?��hr���@VN�灧ٿ��7��&�@K-�]Y 4@:?P�ď!?��hr���@n=h�ٿ���rn��@΍i\G�3@F����!?�*�EB&�@n=h�ٿ���rn��@΍i\G�3@F����!?�*�EB&�@n=h�ٿ���rn��@΍i\G�3@F����!?�*�EB&�@!BC���ٿ�	�m���@���B 4@S�!я!?݉���Y�@!BC���ٿ�	�m���@���B 4@S�!я!?݉���Y�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@�'�6]�ٿ�X3z��@�4�W�4@�v��!?~���t�@���x�ٿ�9�*�@;��� 4@�W๏!?�k��fC�@���x�ٿ�9�*�@;��� 4@�W๏!?�k��fC�@���x�ٿ�9�*�@;��� 4@�W๏!?�k��fC�@���x�ٿ�9�*�@;��� 4@�W๏!?�k��fC�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@2e��x�ٿ6M���w�@�}�& 4@�DEg��!?8 ���u�@��r>��ٿ��<]��@��&V� 4@��	x�!?�����@��r>��ٿ��<]��@��&V� 4@��	x�!?�����@��r>��ٿ��<]��@��&V� 4@��	x�!?�����@��r>��ٿ��<]��@��&V� 4@��	x�!?�����@�W�{��ٿq
�0��@�j��) 4@YN�Gm�!?/��a�@�W�{��ٿq
�0��@�j��) 4@YN�Gm�!?/��a�@�W�{��ٿq
�0��@�j��) 4@YN�Gm�!?/��a�@#�өٿ��5�V�@h�� ��3@���!?wU�`�@#�өٿ��5�V�@h�� ��3@���!?wU�`�@(���U�ٿ&V��$�@���� 4@a�Wُ!?���k���@(���U�ٿ&V��$�@���� 4@a�Wُ!?���k���@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@��j�ٟٿ�(N�$�@���_4@�rd�ߏ!?�������@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@T���^�ٿBJ{0�#�@����N 4@�g�G��!?4����@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@��<녚ٿp��+&�@.v4@��_��!?X�w�ž�@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@;̊���ٿ4�2�'�@yC��4@�a��!?}eYq��@@[�¢ٿ>��S�@O�|��4@�po�ɏ!?�^Dp���@@[�¢ٿ>��S�@O�|��4@�po�ɏ!?�^Dp���@@[�¢ٿ>��S�@O�|��4@�po�ɏ!?�^Dp���@@[�¢ٿ>��S�@O�|��4@�po�ɏ!?�^Dp���@_Y�;��ٿ��0����@��и_ 4@v��%��!?^V��Z��@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���d1�ٿ��F�*��@�UZ�9�3@M�ܢ�!?8k�A�@���e�ٿ���c�@u�p��3@�T)3��!?�0��9��@���e�ٿ���c�@u�p��3@�T)3��!?�0��9��@f�O�l�ٿ�~1��g�@M�n�3@��G�!?���(B
�@�
Ք�ٿ��Ǫ*�@����3@t���m�!?�\��@�
Ք�ٿ��Ǫ*�@����3@t���m�!?�\��@�
Ք�ٿ��Ǫ*�@����3@t���m�!?�\��@�
Ք�ٿ��Ǫ*�@����3@t���m�!?�\��@�
Ք�ٿ��Ǫ*�@����3@t���m�!?�\��@�Ň��ٿ.8��%�@\�R4@��gj�!?wm�S�/�@�Ň��ٿ.8��%�@\�R4@��gj�!?wm�S�/�@�Ň��ٿ.8��%�@\�R4@��gj�!?wm�S�/�@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@q �X?�ٿ1�f���@��.|� 4@�&g���!?�RX���@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@������ٿ����m��@|q�E4@+� ڜ�!?�#�y��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@
�F�]�ٿ�*����@F�<)� 4@��͏!?]��]��@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@���!�ٿ�IQ���@$��ڰ4@PʌӜ�!?}$H���@�[��ɤٿ�wV�u�@�*.��3@z=��e�!?�e}��`�@�[��ɤٿ�wV�u�@�*.��3@z=��e�!?�e}��`�@�[��ɤٿ�wV�u�@�*.��3@z=��e�!?�e}��`�@�[��ɤٿ�wV�u�@�*.��3@z=��e�!?�e}��`�@�[��ɤٿ�wV�u�@�*.��3@z=��e�!?�e}��`�@5$�Gd�ٿ1���Z��@�����3@���*��!?Ql�o�y�@	}����ٿ�i闷�@���N<4@U�����!?a����@	}����ٿ�i闷�@���N<4@U�����!?a����@	}����ٿ�i闷�@���N<4@U�����!?a����@	}����ٿ�i闷�@���N<4@U�����!?a����@	}����ٿ�i闷�@���N<4@U�����!?a����@&t7e�ٿU��۸|�@U.3� 4@�WϏ!?������@/��6>�ٿ֙���@���y��3@���!?���ll�@/��6>�ٿ֙���@���y��3@���!?���ll�@4`�=��ٿޒ��<�@ӽ�0��3@R{-�!?��Q��@4`�=��ٿޒ��<�@ӽ�0��3@R{-�!?��Q��@�R}�ٿ5<�`���@��M۴�3@�T���!?�g Ni@�@�R}�ٿ5<�`���@��M۴�3@�T���!?�g Ni@�@�R}�ٿ5<�`���@��M۴�3@�T���!?�g Ni@�@�R}�ٿ5<�`���@��M۴�3@�T���!?�g Ni@�@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@u,�"2�ٿ���
�@���f��3@6F.�!?W9Jt��@9AXl��ٿ�D �*��@����3@�M�E�!?�X�+ w�@9AXl��ٿ�D �*��@����3@�M�E�!?�X�+ w�@9AXl��ٿ�D �*��@����3@�M�E�!?�X�+ w�@9AXl��ٿ�D �*��@����3@�M�E�!?�X�+ w�@~��D��ٿE���7�@�~u� 4@S����!?֖wT���@~��D��ٿE���7�@�~u� 4@S����!?֖wT���@~��D��ٿE���7�@�~u� 4@S����!?֖wT���@~��D��ٿE���7�@�~u� 4@S����!?֖wT���@��ci!�ٿ�hg�z�@����4@��TX�!?� (���@U$?~�ٿ���;���@��r14@���Ώ!?��"���@U$?~�ٿ���;���@��r14@���Ώ!?��"���@U$?~�ٿ���;���@��r14@���Ώ!?��"���@U$?~�ٿ���;���@��r14@���Ώ!?��"���@�y�Xo�ٿ�ku�&��@�Y4@�8qߏ!?Q�uPΔ�@�y�Xo�ٿ�ku�&��@�Y4@�8qߏ!?Q�uPΔ�@ ��_��ٿP>\��-�@0�� Q 4@B�J.��!?���涐�@ ��_��ٿP>\��-�@0�� Q 4@B�J.��!?���涐�@g��BC�ٿX�若�@�P�o$4@����I�!?؛.���@g��BC�ٿX�若�@�P�o$4@����I�!?؛.���@g��BC�ٿX�若�@�P�o$4@����I�!?؛.���@g��BC�ٿX�若�@�P�o$4@����I�!?؛.���@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@�*׷�ٿ�;Uz�r�@��%W4@kt����!?�$��y�@0�,H�ٿ���)���@�j��4@�m���!?�{�r��@0�,H�ٿ���)���@�j��4@�m���!?�{�r��@0�,H�ٿ���)���@�j��4@�m���!?�{�r��@0�,H�ٿ���)���@�j��4@�m���!?�{�r��@�Ҋ�B�ٿ���b���@4��|�4@O�uя!?�_��u�@���!�ٿ�Lv]��@H~�$�4@��>(ŏ!?W݉G;��@���!�ٿ�Lv]��@H~�$�4@��>(ŏ!?W݉G;��@���!�ٿ�Lv]��@H~�$�4@��>(ŏ!?W݉G;��@�M��ٿ����?��@�x���3@����!?-O�8hg�@�M��ٿ����?��@�x���3@����!?-O�8hg�@�V�Hg�ٿf+T����@N�3���3@V۫Ҕ�!?r��-r�@�V�Hg�ٿf+T����@N�3���3@V۫Ҕ�!?r��-r�@�V�Hg�ٿf+T����@N�3���3@V۫Ҕ�!?r��-r�@�V�Hg�ٿf+T����@N�3���3@V۫Ҕ�!?r��-r�@�V�Hg�ٿf+T����@N�3���3@V۫Ҕ�!?r��-r�@am�ԃ�ٿm�.K�@���4@��I�!?@�8	��@am�ԃ�ٿm�.K�@���4@��I�!?@�8	��@am�ԃ�ٿm�.K�@���4@��I�!?@�8	��@am�ԃ�ٿm�.K�@���4@��I�!?@�8	��@am�ԃ�ٿm�.K�@���4@��I�!?@�8	��@�t��	�ٿ��>�O��@\���s4@�]�(�!?5�)�b��@�t��	�ٿ��>�O��@\���s4@�]�(�!?5�)�b��@�t��	�ٿ��>�O��@\���s4@�]�(�!?5�)�b��@�t��	�ٿ��>�O��@\���s4@�]�(�!?5�)�b��@� ��ٿEɘh�@?�fB� 4@ۗ�_G�!?�0��Ŕ�@� ��ٿEɘh�@?�fB� 4@ۗ�_G�!?�0��Ŕ�@UqI+Ѥٿ��d�=�@�vc�  4@<��G�!?�v����@UqI+Ѥٿ��d�=�@�vc�  4@<��G�!?�v����@UqI+Ѥٿ��d�=�@�vc�  4@<��G�!?�v����@UqI+Ѥٿ��d�=�@�vc�  4@<��G�!?�v����@��Q_¦ٿzH�Z�@$�64@i>�z�!?Chۓ��@��q�ʝٿJ4����@aM��; 4@��J\�!?X���@�@��q�ʝٿJ4����@aM��; 4@��J\�!?X���@�@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�j���ٿꕫ&�w�@*)�� 4@V�fg��!?c0��{��@�-�~c�ٿ�8G�x�@T���n�3@P��5�!?���,O�@�-�~c�ٿ�8G�x�@T���n�3@P��5�!?���,O�@�˹dיٿu��Ѻ�@�X�r4@Q�Zߏ!?�d,\���@�˹dיٿu��Ѻ�@�X�r4@Q�Zߏ!?�d,\���@�˹dיٿu��Ѻ�@�X�r4@Q�Zߏ!?�d,\���@�˹dיٿu��Ѻ�@�X�r4@Q�Zߏ!?�d,\���@�˹dיٿu��Ѻ�@�X�r4@Q�Zߏ!?�d,\���@0z��%�ٿb�:Ui�@$����3@�m��!?���!�%�@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@FVz�4�ٿ��K�]�@��~���3@�:m��!?D�c��@7��'4�ٿ�P�[<��@긒O�4@{�C��!?��	��@7��'4�ٿ�P�[<��@긒O�4@{�C��!?��	��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@�2=��ٿ5���=D�@<����4@HX��!?j8�b��@X0!���ٿ��I�@(���(4@Y^�p�!?�@��ܼ�@V4��ٿ���Z�@�o�TF4@jD��!?������@V4��ٿ���Z�@�o�TF4@jD��!?������@�R륞ٿƣ��0�@� �� 4@s�� <�!?�pnXu)�@�R륞ٿƣ��0�@� �� 4@s�� <�!?�pnXu)�@�R륞ٿƣ��0�@� �� 4@s�� <�!?�pnXu)�@�R륞ٿƣ��0�@� �� 4@s�� <�!?�pnXu)�@�[�ۡٿ�Z{���@����4@�ς/z�!?�I&�4�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@߉��R�ٿRdF���@��� 4@^�g$ߏ!?|�ԗ$�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@s��2�ٿj>���@��y� 4@Sns���!?5:K�8�@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�+�G`�ٿ���n��@� U�4@N+E��!?�he] ��@�kP���ٿ�i��Wn�@�5�j��3@չ.���!?��8}`�@�kP���ٿ�i��Wn�@�5�j��3@չ.���!?��8}`�@��	Ǡ�ٿ;��(��@��[��3@�05I��!?\�/�@�����ٿ��=fw��@ �\�| 4@Ճڤ�!?�q�a���@�����ٿ��=fw��@ �\�| 4@Ճڤ�!?�q�a���@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@ 1JP|�ٿF�Tg�x�@�o � 4@�|ǞЏ!?�Z[�?�@����ٿ�e���@mpG��4@��(!�!?���0��@B#�ٟ�ٿ N@�@��@�.Ki�4@��:Xȏ!?�� ���@B#�ٟ�ٿ N@�@��@�.Ki�4@��:Xȏ!?�� ���@B#�ٟ�ٿ N@�@��@�.Ki�4@��:Xȏ!?�� ���@B#�ٟ�ٿ N@�@��@�.Ki�4@��:Xȏ!?�� ���@�@+oЛٿP?����@�����4@E	N���!?i��4���@Ǣ�lO�ٿh�$A�@ġl�P4@��vB��!?g�+"��@Ǣ�lO�ٿh�$A�@ġl�P4@��vB��!?g�+"��@Ǣ�lO�ٿh�$A�@ġl�P4@��vB��!?g�+"��@Ǣ�lO�ٿh�$A�@ġl�P4@��vB��!?g�+"��@Ǣ�lO�ٿh�$A�@ġl�P4@��vB��!?g�+"��@����ٿ��(<�@^rHZ4@���@ď!?2�X����@����ٿ��(<�@^rHZ4@���@ď!?2�X����@{L���ٿOD�Ŷ��@�;�N\4@�p�!?���U�@{L���ٿOD�Ŷ��@�;�N\4@�p�!?���U�@��p��ٿCP����@�Me�p�3@��Vȸ�!?�C/�/*�@��p��ٿCP����@�Me�p�3@��Vȸ�!?�C/�/*�@Y�p��ٿQ*G��@y�!� 4@�K�w��!?��6���@a�L��ٿq&����@�D��H�3@ϡ� G�!?���ب��@a�L��ٿq&����@�D��H�3@ϡ� G�!?���ب��@a�L��ٿq&����@�D��H�3@ϡ� G�!?���ب��@Wp rO�ٿ�f~���@>��� 4@�+E*O�!?�6�?�@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@ϟ���ٿ�p�n���@���9 4@"h�꟏!?�ے���@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@MI��ѧٿ�R��t��@����� 4@2�w�x�!?;yb>�@�f)q�ٿr�V7�4�@2W�� 4@W2O��!?�T�#�@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@����t�ٿ�e�@��@
���4@�	�s��!?���Y��@�NZ�ٿ�V��C,�@�[��4@�<Z�!?����L�@�NZ�ٿ�V��C,�@�[��4@�<Z�!?����L�@�NZ�ٿ�V��C,�@�[��4@�<Z�!?����L�@�NZ�ٿ�V��C,�@�[��4@�<Z�!?����L�@�xN���ٿ0��e���@�%�TN�3@X��b��!?Ճh��}�@�!R��ٿ&L[K~@�@õz���3@�+gz��!?;X[���@�!R��ٿ&L[K~@�@õz���3@�+gz��!?;X[���@�*s�P�ٿm5����@�����3@��*l�!?H?x}I�@��s�ٿ�w/��-�@�p��3@F��7��!?d���Of�@���ٿ�Q����@:u��3@<A͏!?�Zt�h�@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@YxY&	�ٿЏ���@�)k��4@ԸY�Ï!?����@����ٿ��]�&j�@�W��4@�tU_��!?�@c<���@����ٿ��]�&j�@�W��4@�tU_��!?�@c<���@����ٿ��]�&j�@�W��4@�tU_��!?�@c<���@�{�!��ٿ%�`����@:��6E4@f��t�!?��?�g��@�{�!��ٿ%�`����@:��6E4@f��t�!?��?�g��@���d�ٿ���O��@��_�4@{Q�H�!?� ����@���d�ٿ���O��@��_�4@{Q�H�!?� ����@���d�ٿ���O��@��_�4@{Q�H�!?� ����@q�,.�ٿ�:�7��@���\�4@P�>�!?.�i���@��l�ٿ}:A�p�@��"4@��(c�!?��w�@�uƂg�ٿ/��Kg!�@���B�4@nZw�|�!?�u0��e�@�uƂg�ٿ/��Kg!�@���B�4@nZw�|�!?�u0��e�@�uƂg�ٿ/��Kg!�@���B�4@nZw�|�!?�u0��e�@�uƂg�ٿ/��Kg!�@���B�4@nZw�|�!?�u0��e�@qH��_�ٿWǜ;;��@ajMX�4@���$�!?^�uo��@�Ͳٿ���^e�@$���4@�#��H�!?�!�`D��@�!B�ٿ�b�C���@��.��4@0ۊUV�!?p$���@�!B�ٿ�b�C���@��.��4@0ۊUV�!?p$���@�!B�ٿ�b�C���@��.��4@0ۊUV�!?p$���@�!B�ٿ�b�C���@��.��4@0ۊUV�!?p$���@=0�ٿ�ξ��@�6B4@�[���!?<m��,�@=0�ٿ�ξ��@�6B4@�[���!?<m��,�@��m��ٿ<�fj���@x�����3@
/��L�!?ۼ��^�@��m��ٿ<�fj���@x�����3@
/��L�!?ۼ��^�@��m��ٿ<�fj���@x�����3@
/��L�!?ۼ��^�@��D�H�ٿ�x�ǁ�@��mi��3@ZX;�ʏ!?�ܸ;~�@������ٿ��[NF��@ڡ2N 4@W2=��!?�R�� ��@������ٿ��[NF��@ڡ2N 4@W2=��!?�R�� ��@������ٿ��[NF��@ڡ2N 4@W2=��!?�R�� ��@F����ٿ�����E�@"B�Ѣ 4@���5�!?�	悙A�@F����ٿ�����E�@"B�Ѣ 4@���5�!?�	悙A�@W�ma�ٿydIzF��@���e�3@!D=ey�!?.;+^ԭ�@W�ma�ٿydIzF��@���e�3@!D=ey�!?.;+^ԭ�@W�ma�ٿydIzF��@���e�3@!D=ey�!?.;+^ԭ�@W�ma�ٿydIzF��@���e�3@!D=ey�!?.;+^ԭ�@�X���ٿ�馔�&�@V��a�3@t�z�!?���d�l�@�X���ٿ�馔�&�@V��a�3@t�z�!?���d�l�@�X���ٿ�馔�&�@V��a�3@t�z�!?���d�l�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@�J�璤ٿ���Q^s�@��I���3@ў%,׏!?	e�!�@tU!�Ѥٿ��#LOD�@��Qi��3@R�LPU�!?뭾����@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�o��J�ٿ�AeT��@M��-��3@��`
:�!?�o�V-�@�O�)9�ٿ�s�I�@	���� 4@Jw*�Տ!?yئ���@�O�)9�ٿ�s�I�@	���� 4@Jw*�Տ!?yئ���@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@��	d��ٿ����Z4�@�P�s� 4@rI�ß�!?*�hB �@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@���ٿg�E�z��@~`k� 4@�o.홏!?�pߚ��@�ڟ���ٿ���iޚ�@V��� 4@>��0�!?��0d��@�ڟ���ٿ���iޚ�@V��� 4@>��0�!?��0d��@�ڟ���ٿ���iޚ�@V��� 4@>��0�!?��0d��@�ڟ���ٿ���iޚ�@V��� 4@>��0�!?��0d��@�ڟ���ٿ���iޚ�@V��� 4@>��0�!?��0d��@ɹ61�ٿ�Y��(��@��z�E 4@>m�:�!?��W:���@ɹ61�ٿ�Y��(��@��z�E 4@>m�:�!?��W:���@ɹ61�ٿ�Y��(��@��z�E 4@>m�:�!?��W:���@ɹ61�ٿ�Y��(��@��z�E 4@>m�:�!?��W:���@��k�a�ٿ�q��P��@ēl� 4@{���`�!?��Y���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@C`TVפٿ۽��@	��	% 4@� �O��!?�lY���@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@�-A�ٿ����Z�@5��� 4@���G�!?l��� ��@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@	0�M��ٿɺ�@�,�@ÿ�z 4@;����!?��Q�ݸ�@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@��5���ٿ�Z>���@�2ЊF 4@�-�8��!?�̴S��@f����ٿ>G띕�@m��G��3@�,'��!?cP����@f����ٿ>G띕�@m��G��3@�,'��!?cP����@�Si)C�ٿ8��ƙ�@�U����3@��d�n�!?��]z��@�Si)C�ٿ8��ƙ�@�U����3@��d�n�!?��]z��@�Si)C�ٿ8��ƙ�@�U����3@��d�n�!?��]z��@]�]j�ٿl�'|��@�!Q�~ 4@Rq|�!?��g%���@�B���ٿ�V���@��Ir��3@���W��!?�ͬ�@wnC�Ģٿw�_��?�@�	���3@$P�f�!?���e��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@�_��	�ٿ6���c��@NqL!� 4@���}F�!?��j��@]LA-�ٿI��Q6��@��W4@��MCI�!?�;��@���i2�ٿ����*�@k$��4@�7��H�!?��MM��@���i2�ٿ����*�@k$��4@�7��H�!?��MM��@���i2�ٿ����*�@k$��4@�7��H�!?��MM��@��vWu�ٿ,�mSq��@_o5P�4@��DJ�!?�nU�|�@��vWu�ٿ,�mSq��@_o5P�4@��DJ�!?�nU�|�@�:�P��ٿ�"���y�@�!Җt4@8*#���!?l�����@�:�P��ٿ�"���y�@�!Җt4@8*#���!?l�����@�:�P��ٿ�"���y�@�!Җt4@8*#���!?l�����@�:�P��ٿ�"���y�@�!Җt4@8*#���!?l�����@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�X�z�ٿؤ�9�!�@�Tj4@>~_�!?��2_�4�@�b`��ٿ��f`���@/*�� 4@n7�I�!?�x�1�@�}��Ҡٿ��$
�@�o�� 4@ad��c�!?D���m�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@�>k��ٿ��@B��@�Կ�	 4@�8�pȏ!?�솫!�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@������ٿ��L���@@b�"B 4@����!?�`�N4�@�Y��6�ٿ
Ғ���@������3@��ؔ��!?-2�g��@�Y��6�ٿ
Ғ���@������3@��ؔ��!?-2�g��@�Y��6�ٿ
Ғ���@������3@��ؔ��!?-2�g��@f�Jir�ٿ�H'���@g�$O4@���Kl�!?��C��@��O��ٿ$6����@;ʒU� 4@7�浏!?{�����@��O��ٿ$6����@;ʒU� 4@7�浏!?{�����@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@�ł%[�ٿ.Œ����@�́� 4@}$���!?'X�r>��@��g�ٿ�TG� �@�2z�4@��ƪȏ!?������@��g�ٿ�TG� �@�2z�4@��ƪȏ!?������@��g�ٿ�TG� �@�2z�4@��ƪȏ!?������@��z�ٿ�e�{�@L;�&��3@?���ď!?Ub��w�@��z�ٿ�e�{�@L;�&��3@?���ď!?Ub��w�@��z�ٿ�e�{�@L;�&��3@?���ď!?Ub��w�@��z�ٿ�e�{�@L;�&��3@?���ď!?Ub��w�@�W��ٿ��*���@�v���4@m����!?_�-��@VT>[s�ٿ}fGP�"�@4 �4@ l�1��!?W��@VT>[s�ٿ}fGP�"�@4 �4@ l�1��!?W��@VT>[s�ٿ}fGP�"�@4 �4@ l�1��!?W��@��s�ٿ�/��Q�@�X]�I4@���!?A��N��@��s�ٿ�/��Q�@�X]�I4@���!?A��N��@��s�ٿ�/��Q�@�X]�I4@���!?A��N��@��s�ٿ�/��Q�@�X]�I4@���!?A��N��@��s�ٿ�/��Q�@�X]�I4@���!?A��N��@N0W�&�ٿ�ħ�!�@.g̨�3@�~���!?�.����@N0W�&�ٿ�ħ�!�@.g̨�3@�~���!?�.����@a� �*�ٿsP)��@5��� 4@�цa��!?�~�2���@a� �*�ٿsP)��@5��� 4@�цa��!?�~�2���@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@�p����ٿ��EH&��@?��'� 4@$Ӑ��!?zײ�E��@ /7Q��ٿ�:�&�`�@�2�a� 4@�C�Q��!?�s��D��@ /7Q��ٿ�:�&�`�@�2�a� 4@�C�Q��!?�s��D��@ /7Q��ٿ�:�&�`�@�2�a� 4@�C�Q��!?�s��D��@����ٿ��k��@"��ff 4@�_���!?N����Y�@��E�ƣٿ��λr1�@�4�[� 4@�G=*��!?�Rc~j�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@�~�&��ٿ�cO���@��խ 4@!,W���!?,r_�n�@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@���Pݤٿ8���m�@��K:�4@~���i�!?>[�3���@FZ�%�ٿ%>q�]�@Hx��$ 4@R��m��!?ܿx\�|�@FZ�%�ٿ%>q�]�@Hx��$ 4@R��m��!?ܿx\�|�@�4�N�ٿ���� �@/�v?� 4@��M�!?A�f����@�4�N�ٿ���� �@/�v?� 4@��M�!?A�f����@�4�N�ٿ���� �@/�v?� 4@��M�!?A�f����@���6РٿX��u%�@�N�L4@���!?귉",�@���6РٿX��u%�@�N�L4@���!?귉",�@���6РٿX��u%�@�N�L4@���!?귉",�@���6РٿX��u%�@�N�L4@���!?귉",�@���6РٿX��u%�@�N�L4@���!?귉",�@=���x�ٿ�|ycT�@���T4@��Hӏ!?#w@H�	�@x���A�ٿm��w|�@�{��4@�]Qa�!?r�p ��@x���A�ٿm��w|�@�{��4@�]Qa�!?r�p ��@x���A�ٿm��w|�@�{��4@�]Qa�!?r�p ��@�g����ٿ�;����@���I�4@)X0Yx�!?:��P���@���`z�ٿ2�=`d&�@��.m'4@��Q��!?���xo�@���`z�ٿ2�=`d&�@��.m'4@��Q��!?���xo�@���`z�ٿ2�=`d&�@��.m'4@��Q��!?���xo�@���`z�ٿ2�=`d&�@��.m'4@��Q��!?���xo�@}0�+t�ٿ,w����@mO�Dw4@,�(쏏!?fL�,=#�@K��1ީٿDh�����@Q�'4@U�l�W�!?�=y����@d��c�ٿ������@��7Ki4@z?L���!?�L��/�@d��c�ٿ������@��7Ki4@z?L���!?�L��/�@d��c�ٿ������@��7Ki4@z?L���!?�L��/�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@�f���ٿC��z[�@�2'lc4@���!��!??k
�	�@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@zٵ�ҟٿ;a7��d�@��Ԛ�3@u�V�֏!?�����@�Ҹ�ٿ~�T	�@O�A�� 4@���ߏ!?�S��o�@�Ҹ�ٿ~�T	�@O�A�� 4@���ߏ!?�S��o�@�Ҹ�ٿ~�T	�@O�A�� 4@���ߏ!?�S��o�@�Ҹ�ٿ~�T	�@O�A�� 4@���ߏ!?�S��o�@�Ҹ�ٿ~�T	�@O�A�� 4@���ߏ!?�S��o�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@mV�7��ٿtZr����@3���� 4@�n�q��!?IM��3�@* YV�ٿ�����@�1fp4@���֏!?F�\����@* YV�ٿ�����@�1fp4@���֏!?F�\����@* YV�ٿ�����@�1fp4@���֏!?F�\����@* YV�ٿ�����@�1fp4@���֏!?F�\����@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@���D��ٿ����T�@�%�F�4@�kƎ��!?B��ȥ�@IrW�J�ٿ�㾸���@���4@��1�9�!?����0��@IrW�J�ٿ�㾸���@���4@��1�9�!?����0��@IrW�J�ٿ�㾸���@���4@��1�9�!?����0��@�N�ٿ��3l��@n�h?4@.#l�!?�#.z���@�N�ٿ��3l��@n�h?4@.#l�!?�#.z���@�N�ٿ��3l��@n�h?4@.#l�!?�#.z���@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�x՟إٿ��<<#��@"vk�� 4@ 9ەl�!?w�
�=�@�Ք�Y�ٿ���x��@�t�A�4@��*8�!?�%�B�@�Ք�Y�ٿ���x��@�t�A�4@��*8�!?�%�B�@�Ք�Y�ٿ���x��@�t�A�4@��*8�!?�%�B�@�Ք�Y�ٿ���x��@�t�A�4@��*8�!?�%�B�@�Ք�Y�ٿ���x��@�t�A�4@��*8�!?�%�B�@�M(�I�ٿHyx�
��@<�ɨ; 4@m�*���!?%�Sn�@�M(�I�ٿHyx�
��@<�ɨ; 4@m�*���!?%�Sn�@�M(�I�ٿHyx�
��@<�ɨ; 4@m�*���!?%�Sn�@�M(�I�ٿHyx�
��@<�ɨ; 4@m�*���!?%�Sn�@�M(�I�ٿHyx�
��@<�ɨ; 4@m�*���!?%�Sn�@Y�8��ٿ��|���@F��74@��pE2�!?�&����@�Y�n�ٿVk6-��@���f4@'՜��!?����h�@�Y�n�ٿVk6-��@���f4@'՜��!?����h�@�Y�n�ٿVk6-��@���f4@'՜��!?����h�@�Y�n�ٿVk6-��@���f4@'՜��!?����h�@�Y�n�ٿVk6-��@���f4@'՜��!?����h�@V��Ƞٿ}?��@��@ꪩ��4@�Ns�!?�{�/��@V��Ƞٿ}?��@��@ꪩ��4@�Ns�!?�{�/��@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@z�?��ٿ�*S��@��� 4@�{��!?nEM��:�@FY��q�ٿzL[��@� � 4@�G���!?�h��6�@FY��q�ٿzL[��@� � 4@�G���!?�h��6�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��Q���ٿ] ��lI�@g�h���3@�&Ar�!?sz�Z*�@��LⳙٿU�g���@�x9/E�3@%��gy�!?�1�����@��LⳙٿU�g���@�x9/E�3@%��gy�!?�1�����@��LⳙٿU�g���@�x9/E�3@%��gy�!?�1�����@��̷�ٿ~��'���@p�	j 4@M
��!?�K�
{�@�x;�`�ٿ�8Es�@��q�04@�-�v�!?���U�@�x;�`�ٿ�8Es�@��q�04@�-�v�!?���U�@�x;�`�ٿ�8Es�@��q�04@�-�v�!?���U�@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�SW�C�ٿ��O4g�@Gzг� 4@�Q�h�!?�wE���@�vB�ٿ��2����@f���C4@:���R�!?Bo1�z~�@�vB�ٿ��2����@f���C4@:���R�!?Bo1�z~�@�vB�ٿ��2����@f���C4@:���R�!?Bo1�z~�@�vB�ٿ��2����@f���C4@:���R�!?Bo1�z~�@~H�g�ٿ�-�[�m�@��� 4@�Gn�M�!?��7� L�@���\:�ٿ=��+;G�@�
7Z 4@��T�x�!?c�&��@���\:�ٿ=��+;G�@�
7Z 4@��T�x�!?c�&��@���\:�ٿ=��+;G�@�
7Z 4@��T�x�!?c�&��@���\:�ٿ=��+;G�@�
7Z 4@��T�x�!?c�&��@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@��&f�ٿ�$^i��@=p�4@�n�Ϗ!?8/��+�@�0�ٿ�Y#�@T�@�`�4@:vz��!?��T09��@�a^���ٿs-$0���@��F4@�i�ɺ�!?�����@�a^���ٿs-$0���@��F4@�i�ɺ�!?�����@�a^���ٿs-$0���@��F4@�i�ɺ�!?�����@�a^���ٿs-$0���@��F4@�i�ɺ�!?�����@�a^���ٿs-$0���@��F4@�i�ɺ�!?�����@7}X<��ٿ�h)�}��@��'F4@�
�r׏!?��o:��@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@�\F؝ٿ�F�2.��@_%'� 4@a.o��!?�@����@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@c	����ٿF5�y��@�<M� 4@c۹��!?r�㠽�@�NsC�ٿ�E�[��@I�C�3@��( }�!?C��)+��@�NsC�ٿ�E�[��@I�C�3@��( }�!?C��)+��@�NsC�ٿ�E�[��@I�C�3@��( }�!?C��)+��@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@59�H�ٿU�#����@�֣�% 4@��5ԏ!?2���L�@�b_'��ٿ�X����@�ړ��3@�*z�!?�q�#g��@5Y��ٿ��/����@�����3@��*&��!?= �����@5Y��ٿ��/����@�����3@��*&��!?= �����@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@S��L�ٿ����.}�@�� (?�3@�Y����!?�MC
�@j7Gi��ٿ��S��X�@���\ 4@��^���!?[�Zf��@�}�ٿY��ܾ�@%N>� 4@2�+��!?�_t�]��@�}�ٿY��ܾ�@%N>� 4@2�+��!?�_t�]��@�}�ٿY��ܾ�@%N>� 4@2�+��!?�_t�]��@�}�ٿY��ܾ�@%N>� 4@2�+��!?�_t�]��@	z��ٿ{EW?��@��H�^4@��5�F�!?)���t�@	z��ٿ{EW?��@��H�^4@��5�F�!?)���t�@	z��ٿ{EW?��@��H�^4@��5�F�!?)���t�@��i�~�ٿ����@�[�D�4@��ٗ�!? ����@��i�~�ٿ����@�[�D�4@��ٗ�!? ����@a���ٿ.qx���@��ݵ}4@J�-͏!?������@a���ٿ.qx���@��ݵ}4@J�-͏!?������@*%�Z[�ٿc�����@Q�4@�g.Z��!?�k��A��@*%�Z[�ٿc�����@Q�4@�g.Z��!?�k��A��@*%�Z[�ٿc�����@Q�4@�g.Z��!?�k��A��@*%�Z[�ٿc�����@Q�4@�g.Z��!?�k��A��@*%�Z[�ٿc�����@Q�4@�g.Z��!?�k��A��@�wK��ٿL�~�Ȱ�@I���64@�#����!?ӏ{�O��@�wK��ٿL�~�Ȱ�@I���64@�#����!?ӏ{�O��@�wK��ٿL�~�Ȱ�@I���64@�#����!?ӏ{�O��@a��RN�ٿ�`,�@���9{4@^<��!?��F~�@a��RN�ٿ�`,�@���9{4@^<��!?��F~�@a��RN�ٿ�`,�@���9{4@^<��!?��F~�@a��RN�ٿ�`,�@���9{4@^<��!?��F~�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�%V�ٿ����@����� 4@�nƀ�!?��1`؄�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@�2�RN�ٿY�}i�@ G�]�3@[.�Ư�!?����[/�@Dj\|�ٿo�
� �@tbZ+v�3@��'���!?f`*$M�@mJ��ٿ/,�P�*�@�h��3@ҳ�!?�X�BEx�@mJ��ٿ/,�P�*�@�h��3@ҳ�!?�X�BEx�@mJ��ٿ/,�P�*�@�h��3@ҳ�!?�X�BEx�@ �Ў:�ٿ�a��`t�@��z�X�3@��ޏ!?���	��@ �Ў:�ٿ�a��`t�@��z�X�3@��ޏ!?���	��@ �Ў:�ٿ�a��`t�@��z�X�3@��ޏ!?���	��@�$ƨZ�ٿ�Y����@��C�d�3@*:O���!?W
,�m��@ݕ���ٿ��.���@ן/4@�u����!?$⼔���@�>�7�ٿ>p��cT�@b�~��3@��A�P�!?���v!�@�>�7�ٿ>p��cT�@b�~��3@��A�P�!?���v!�@�>�7�ٿ>p��cT�@b�~��3@��A�P�!?���v!�@�B�hW�ٿz��B��@+PJ'� 4@���!?�d�l�@;�K0�ٿm��+X��@u�q�4@$���!?z~����@���ٿ��U �@���4@t'%y܏!?��"�),�@���ٿ��U �@���4@t'%y܏!?��"�),�@���ٿ��U �@���4@t'%y܏!?��"�),�@���ٿ��U �@���4@t'%y܏!?��"�),�@���ٿ��U �@���4@t'%y܏!?��"�),�@���ٿ��U �@���4@t'%y܏!?��"�),�@��1d�ٿK�4��@�a��4@�#�ҏ!?{�?\��@��1d�ٿK�4��@�a��4@�#�ҏ!?{�?\��@��1d�ٿK�4��@�a��4@�#�ҏ!?{�?\��@��1d�ٿK�4��@�a��4@�#�ҏ!?{�?\��@��1d�ٿK�4��@�a��4@�#�ҏ!?{�?\��@��e�ٿ3���@���4@?9�av�!?�n��@��.K��ٿ&v �@�$=�4@o\ꀙ�!?t��_�@��.K��ٿ&v �@�$=�4@o\ꀙ�!?t��_�@��.K��ٿ&v �@�$=�4@o\ꀙ�!?t��_�@��.K��ٿ&v �@�$=�4@o\ꀙ�!?t��_�@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@x'�۠ٿ)�@����@��3	4@=h��p�!?14�շ��@�3>��ٿ+N�{��@�
o��4@�퍣ޏ!?Z�n��$�@#+��˝ٿ��L��@8��w>4@4�?��!?'`y�-�@#+��˝ٿ��L��@8��w>4@4�?��!?'`y�-�@#+��˝ٿ��L��@8��w>4@4�?��!?'`y�-�@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@�	�q�ٿ����_�@3�ƥL4@:ֳ�!?��-b���@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��5~�ٿ}6Ą�@�u8d4@z�q�ԏ!?�<G�{�@��d�ٿ�8z)�@��}0� 4@x�d�;�!?��&��@��d�ٿ�8z)�@��}0� 4@x�d�;�!?��&��@g8�Ϊٿ[��F��@�Oۣ��3@Z���:�!?x)+%��@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@�C�Y�ٿFb<?Y5�@%Ӥ�[�3@������!?��C?$q�@{�8��ٿx��pO�@7&�7%�3@��*vr�!?����Y#�@�Gw���ٿ�8u���@��F"* 4@��
��!?!�F�w��@�Gw���ٿ�8u���@��F"* 4@��
��!?!�F�w��@���ڟٿO"����@Kwm� 4@N�g6��!?Z����#�@�*Q���ٿÙf�jb�@#���u�3@>(���!?p/�t&�@�*Q���ٿÙf�jb�@#���u�3@>(���!?p/�t&�@�*Q���ٿÙf�jb�@#���u�3@>(���!?p/�t&�@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@�<�|�ٿ������@9�H�3@p�����!?ֻ��u��@0��p��ٿQ�����@�}��� 4@���4k�!?L��@0��p��ٿQ�����@�}��� 4@���4k�!?L��@0��p��ٿQ�����@�}��� 4@���4k�!?L��@0��p��ٿQ�����@�}��� 4@���4k�!?L��@����ݩٿ��*!�@�3�y� 4@�Hu���!?�zx��@����ݩٿ��*!�@�3�y� 4@�Hu���!?�zx��@����ݩٿ��*!�@�3�y� 4@�Hu���!?�zx��@<I��j�ٿ�F
8=�@9,G�_ 4@���ߴ�!?���zp�@<I��j�ٿ�F
8=�@9,G�_ 4@���ߴ�!?���zp�@<I��j�ٿ�F
8=�@9,G�_ 4@���ߴ�!?���zp�@Q>�xZ�ٿy�(�1c�@O6�4@j2╏!?�1�VC�@����ٿ#)�|M��@�.��4@���E�!?H`a�\��@����ٿ#)�|M��@�.��4@���E�!?H`a�\��@P�D�ٿ1��)�~�@���4@���=�!?#C`V��@P�D�ٿ1��)�~�@���4@���=�!?#C`V��@P�D�ٿ1��)�~�@���4@���=�!?#C`V��@m7F��ٿ�K���@�t�l4@_�1P��!?��f�@m7F��ٿ�K���@�t�l4@_�1P��!?��f�@m7F��ٿ�K���@�t�l4@_�1P��!?��f�@m7F��ٿ�K���@�t�l4@_�1P��!?��f�@�+�p2�ٿ�qڰ�@0�jp4@�n����!?�m&�ݵ�@�+�p2�ٿ�qڰ�@0�jp4@�n����!?�m&�ݵ�@�+�p2�ٿ�qڰ�@0�jp4@�n����!?�m&�ݵ�@�+�p2�ٿ�qڰ�@0�jp4@�n����!?�m&�ݵ�@r��K�ٿ�o,�}P�@o��4@����!?��|���@0�_���ٿܻgJO�@í1�g 4@����Ï!?��ɢ���@0�_���ٿܻgJO�@í1�g 4@����Ï!?��ɢ���@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@�.�Ȩٿ8Q�s��@b�mi�3@
�ҏ�!?���oV��@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@ڂ;p��ٿ�;�[��@�s���3@�Ry�!?̤]����@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@�� 5+�ٿ�;?����@�Ԥ��4@@%�z�!?XN8�O��@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@������ٿ     ��@      4@�t><K�!?�ň��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@p)����ٿ&������@cY�a 4@s���_�!?ѻ��o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�:�̙ٿ������@ڧ�� 4@|��Ɠ�!?`���o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@�[���ٿ�Ac����@�ڙ
 4@�>|?��!?0��o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@y@�Ѵ�ٿ�r����@�%h 4@�@��!?�����o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@s"�i��ٿ^�߾���@���0 4@bzlՏ!?7�,��o�@��L���ٿ?(:����@tF� 4@���!?�� ��o�@��L���ٿ?(:����@tF� 4@���!?�� ��o�@��L���ٿ?(:����@tF� 4@���!?�� ��o�@��L���ٿ?(:����@tF� 4@���!?�� ��o�@��L���ٿ?(:����@tF� 4@���!?�� ��o�@� �Ùٿ��}����@R�� 4@���1(�!?�I���o�@� �Ùٿ��}����@R�� 4@���1(�!?�I���o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@~�vJřٿ�����@~Ʋ� 4@Զ��ޏ!?�:e��o�@��șٿ[�����@:	 4@l�s�!?�����o�@ڂ�șٿm�����@� 4@��\�!?}ˑ��o�@�ɺ@̙ٿ�?H����@���s 4@N��Gx�!?�Y���o�@�ɺ@̙ٿ�?H����@���s 4@N��Gx�!?�Y���o�@��7�ƙٿtf�����@$x�r 4@��u�!?`���o�@��7�ƙٿtf�����@$x�r 4@��u�!?`���o�@��7�ƙٿtf�����@$x�r 4@��u�!?`���o�@��7�ƙٿtf�����@$x�r 4@��u�!?`���o�@��7�ƙٿtf�����@$x�r 4@��u�!?`���o�@3��ęٿ�����@�MP�
 4@}��o�!?_���o�@3��ęٿ�����@�MP�
 4@}��o�!?_���o�@�SJ���ٿ-�ӹ���@M��
 4@������!?�V���o�@�SJ���ٿ-�ӹ���@M��
 4@������!?�V���o�@�SJ���ٿ-�ӹ���@M��
 4@������!?�V���o�@�SJ���ٿ-�ӹ���@M��
 4@������!?�V���o�@G����ٿT\�����@�4%�
 4@^Ē���!?���o�@G����ٿT\�����@�4%�
 4@^Ē���!?���o�@W��q��ٿq�����@cH��
 4@����Ϗ!?8����o�@W��q��ٿq�����@cH��
 4@����Ϗ!?8����o�@���E��ٿԀS����@yL�
 4@�����!?T����o�@���W��ٿ@g�����@�J
 4@���!?qB���o�@��.ʹ�ٿ��Q����@w;�
 4@7�#}��!?~#��o�@(n�b��ٿ[�غ���@���O	 4@���^r�!?��O��o�@�C�/��ٿ�Ɩ����@H)U� 4@`���2�!?
���o�@X�����ٿ�����@۬ 4@��B�!?�1���o�@A��!��ٿ:������@�� 4@,ᰲ��!?'��o�@P�tB��ٿ������@��m 4@��i܏!?�T��o�@+պ��ٿ�/f����@ӊ�R 4@��&�!?TՏ��o�@ ��0��ٿ�r����@)��g	 4@C���!�!?mH���o�@�:�ٿ�a�����@�Ѓ� 4@ƞ��j�!?�r��o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@���ٿ�����@���k 4@&hֈO�!?�����o�@�t>Q��ٿ<�����@����	 4@�(疏!?�n���o�@X�H��ٿ
�(����@�mw	 4@ʡaϏ!?��u��o�@X�H��ٿ
�(����@�mw	 4@ʡaϏ!?��u��o�@C��ɶ�ٿ������@G� \	 4@	�+n��!?�"D��o�@�Kp��ٿu������@����	 4@#���!?�k<��o�@�Kp��ٿu������@����	 4@#���!?�k<��o�@�b ��ٿ�1����@�� 4@�\$(��!?����o�@R~�࿙ٿN������@�f 4@���!?2Z���o�@R~�࿙ٿN������@�f 4@���!?2Z���o�@��>��ٿ������@ b	 4@��[�!?�S���o�@~z�о�ٿO������@h,�� 4@�����!?/̴��o�@~z�о�ٿO������@h,�� 4@�����!?/̴��o�@�����ٿ�';����@��? 4@�l8Q�!?ͷо�o�@q�|ٿ$�Y����@]\;�
 4@�	�6�!??�߹�o�@q�|ٿ$�Y����@]\;�
 4@�	�6�!??�߹�o�@q�|ٿ$�Y����@]\;�
 4@�	�6�!??�߹�o�@���ÙٿL�����@I� 4@>!�j�!?@�й�o�@���ÙٿL�����@I� 4@>!�j�!?@�й�o�@*���řٿE*�����@��V 4@�`+��!?���o�@*���řٿE*�����@��V 4@�`+��!?���o�@�x�vřٿ��'����@_R=�
 4@�t��s�!?�K��o�@�%`ęٿ�;�����@/�4 4@���ŏ!?�땶�o�@(yeęٿ�������@�oK�
 4@�w�:��!?è6��o�@(yeęٿ�������@�oK�
 4@�w�:��!?è6��o�@n+e��ٿ/r�����@7��)
 4@�0G\�!?�bG��o�@��軙ٿJ������@���
 4@k��v�!?��t��o�@�j$��ٿ[�����@k���
 4@�4(w�!?�Q��o�@u�����ٿ������@A�0�	 4@����l�!?����o�@�J��ٿ�43����@���	 4@0��l�!?�=���o�@�J��ٿ�43����@���	 4@0��l�!?�=���o�@lA����ٿl������@TF�	 4@������!?5p���o�@g>�ݵ�ٿ�Ż����@��7�	 4@F��ȏ!?z���o�@g>�ݵ�ٿ�Ż����@��7�	 4@F��ȏ!?z���o�@g>�ݵ�ٿ�Ż����@��7�	 4@F��ȏ!?z���o�@��̵�ٿ��F����@���.	 4@�FW�|�!? 0���o�@��̵�ٿ��F����@���.	 4@�FW�|�!? 0���o�@;)=��ٿ�p�����@�Rx	 4@4����!?�Һ�o�@y���ٿ	������@/5Ee	 4@�'����!?�ϸ�o�@(�)���ٿ������@,�*	 4@U��!?Lj��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@0���ٿI i����@=;�_	 4@N����!?��:��o�@��n]��ٿ,����@@iJ�	 4@���z�!?2���o�@��n]��ٿ,����@@iJ�	 4@���z�!?2���o�@ҦP��ٿ"7�����@����	 4@Wx�]�!?k����o�@ҦP��ٿ"7�����@����	 4@Wx�]�!?k����o�@�gt��ٿ�U����@�@8/	 4@����!?� 7��o�@�gt��ٿ�U����@�@8/	 4@����!?� 7��o�@�Q�ٿ||�����@��L� 4@��f��!?�(���o�@�Q�ٿ||�����@��L� 4@��f��!?�(���o�@������ٿ<M����@h� 4@�r���!?t���o�@������ٿ<M����@h� 4@�r���!?t���o�@�y*��ٿ�!�����@�2I	 4@���!�!?V���o�@�ޕ��ٿ��
����@�$	 4@!�Pa��!?�����o�@�ޕ��ٿ��
����@�$	 4@!�Pa��!?�����o�@�Wm��ٿ-c�����@"4�e	 4@j�aC��!?Uc���o�@���K��ٿ�����@��H	 4@_�)���!?�����o�@��1���ٿ�������@�JA|	 4@2��p�!?j��o�@t�!���ٿ8J����@(�Ό	 4@�|q߶�!?��H��o�@��Z��ٿ������@PI��	 4@ �]C��!?�W��o�@���p��ٿ{�����@����	 4@Ɓ�q�!?0���o�@�����ٿ;������@ǥ'
 4@�;z��!?vg��o�@�$���ٿ�2�����@� 
 4@c�mJŏ!?Q���o�@*�Y��ٿ;,�����@�X�f	 4@�/�ُ!?����o�@ n�ٿ������@���	 4@(a��!?��o�@	�ʅ��ٿ������@�	 4@`~p��!?�4���o�@�>Hr��ٿ�������@V�>h	 4@z�I�ڏ!?�ĉ��o�@�����ٿH;k����@.�g� 4@Õ '�!?�k���o�@�����ٿH;k����@.�g� 4@Õ '�!?�k���o�@r&���ٿ�������@�=�� 4@'e���!?=����o�@(7���ٿ������@9��p 4@�7��֏!?�`���o�@(7���ٿ������@9��p 4@�7��֏!?�`���o�@ݰ|���ٿ2������@'H^ 4@ ��夏!?��o�@�-���ٿ������@�ף 4@��M��!?����o�@�-���ٿ������@�ף 4@��M��!?����o�@5�����ٿ��7����@�XzQ 4@>���!?uG���o�@�,����ٿeV����@uVF
 4@%����!?u����o�@�D����ٿ;����@��� 4@�+ی�!?Zxu��o�@�D����ٿ;����@��� 4@�+ی�!?Zxu��o�@E2�ٿ<�:����@y{�� 4@+�Ï!?����o�@��*T��ٿx�w����@�c�� 4@������!?��%��o�@��*T��ٿx�w����@�c�� 4@������!?��%��o�@(�����ٿ̯�����@��@ 4@��c�!?�ƕ��o�@c�tw��ٿ��!����@��I 4@�#��Ǐ!?�E��o�@��5���ٿ7N%����@�{: 4@e=�#��!?�����o�@}9^��ٿ2�v����@�'�� 4@��일�!?omZ��o�@B��d��ٿ�aU����@�6.M 4@D�0�ɏ!?��4��o�@Q�>���ٿi������@f�1� 4@�T��ӏ!?d�6��o�@VyY멙ٿ������@b��� 4@��,�Ǐ!?g]��o�@#�^E��ٿL<�����@��O 4@�ƄЏ!?�^���o�@��M���ٿ�F�����@��]� 4@7�%ٽ�!?��=��o�@������ٿ�o����@��V 4@$����!?O����o�@�y���ٿӹ�����@�uw 4@�5����!?Z����o�@�y���ٿӹ�����@�uw 4@�5����!?Z����o�@��֯�ٿ�,����@i�6 4@���ŏ!?����o�@$V����ٿ�������@8-( 4@�����!?h���o�@Z�!ޮ�ٿJ)����@˲� 4@
GJY
�!?%o���o�@�Юլ�ٿr.L����@��"� 4@���=�!?f����o�@Ȟ�"��ٿ'h�����@�6N� 4@�7���!?$Z��o�@Q� ���ٿ�f�����@.*hU 4@tHD��!?�3���o�@Q� ���ٿ�f�����@.*hU 4@tHD��!?�3���o�@L��y��ٿ��a����@Cu�" 4@��^���!?л���o�@n�O��ٿ������@�H 4@� 4R�!?�]e��o�@n�O��ٿ������@�H 4@� 4R�!?�]e��o�@��DŪ�ٿ{�F����@��?� 4@ċ����!?�����o�@r�NU��ٿ�]�����@���� 4@ћ���!?a���o�@����ٿ������@I�m� 4@ٹ���!?�����o�@\�2��ٿG�����@'� 4@*=I�z�!?G4��o�@\�2��ٿG�����@'� 4@*=I�z�!?G4��o�@��/q��ٿ}�E����@ؙL� 4@�-�Gp�!?��R��o�@ޱM��ٿ��\����@�l�� 4@��܅�!?�ˑ��o�@uu���ٿ.�����@��S` 4@�Q���!?��R��o�@1��/��ٿ�@�����@lh�  4@*m�c�!?�%���o�@�iy��ٿ3������@ǊP  4@��_�K�!?tf���o�@�U����ٿ�R�����@B�  4@�s���!?g���o�@�&-���ٿ��:����@�;Q���3@3�|��!?��.��o�@��r��ٿ:������@4�Ҍ 4@P��ԓ�!? ����o�@��r��ٿ:������@4�Ҍ 4@P��ԓ�!? ����o�@$�e��ٿ9D�����@��Q� 4@�w�a��!?��*��o�@,ᷙٿT�'����@���" 4@��$E��!?z����o�@/�\wǙٿ]�����@p�
 4@*D_s�!?��M��o�@� �řٿ�|����@'��\ 4@��VM�!?"0U��o�@� �řٿ�|����@'��\ 4@��VM�!?"0U��o�@EkX�Ιٿ�������@L�� 4@���X�!?K�-��o�@X���֙ٿvF�����@�)i 4@��`��!?2����o�@��%�љٿg������@��� 4@��ӫ�!?�^���o�@�i�əٿ�q8����@gތn 4@�D6���!?ޣ���o�@E�2/љٿ�������@$n4
 4@<�@i�!?����o�@$���ƙٿ�y�����@ Ɏ 4@�]|ݘ�!?l���o�@� �əٿ8=����@�"W  4@�9�s�!?�ͯ�o�@� �əٿ8=����@�"W  4@�9�s�!?�ͯ�o�@� �əٿ8=����@�"W  4@�9�s�!?�ͯ�o�@� �əٿ8=����@�"W  4@�9�s�!?�ͯ�o�@g5�}әٿ[Z����@�L� 4@_��G�!?2���o�@��B�ٿz�����@���� 4@{���=�!?Aʶ�o�@�^O�ڙٿ@�����@��4 4@'\K�g�!?G�s��o�@�^O�ڙٿ@�����@��4 4@'\K�g�!?G�s��o�@4�ٿ��S����@��y� 4@�IvZ��!?Z���o�@�P6Iיٿ�U�����@��xv 4@YiS�!?�?���o�@����ƙٿp>[����@�̛ 4@@�5��!?v�ٲ�o�@u���Йٿ������@��l� 4@I}���!?#-k��o�@u���Йٿ������@��l� 4@I}���!?#-k��o�@���,ʙٿJY����@i�d 4@�b���!?ǻͬ�o�@���,ʙٿJY����@i�d 4@�b���!?ǻͬ�o�@���,ʙٿJY����@i�d 4@�b���!?ǻͬ�o�@���.ęٿ	f"����@��[? 4@����!?����o�@�%ؙٿI �����@ІO� 4@cה1ҏ!?KL$��o�@�%ؙٿI �����@ІO� 4@cה1ҏ!?KL$��o�@�	a(�ٿI�����@���+ 4@2�I��!?�e���o�@���Nޙٿ�����@Y[89# 4@����ޏ!?�j���o�@����ޙٿƲ(����@���z# 4@�>��!?H����o�@����ޙٿƲ(����@���z# 4@�>��!?H����o�@����ޙٿƲ(����@���z# 4@�>��!?H����o�@����ޙٿƲ(����@���z# 4@�>��!?H����o�@����ޙٿƲ(����@���z# 4@�>��!?H����o�@�c֙ٿɫ�����@�F�w 4@k&�!?���o�@�:|Gљٿ�mS����@��� 4@��U�ҏ!?�Wz��o�@���͙ٿ4 u����@)C� 4@*�s��!?L�B��o�@UԻ���ٿ%Fa����@����
 4@@N�띏!?�5���o�@������ٿ������@�h 4@�斺ɏ!?�R0��o�@#/�ϙٿP7�����@�T�� 4@�} ��!?��w��o�@3����ٿK�U����@oƘk 4@�7��!?5/��o�@3����ٿK�U����@oƘk 4@�7��!?5/��o�@V֖řٿ�?p����@���
 4@�şNG�!?>`��o�@�8�]��ٿ�*G����@a�b� 4@��d�R�!?�����o�@�8�]��ٿ�*G����@a�b� 4@��d�R�!?�����o�@�
�Dәٿ�����@��7 4@�H�!?ޖ��o�@�
�Dәٿ�����@��7 4@�H�!?ޖ��o�@s�!��ٿ�u�����@���	 4@�<l�Q�!?1U*��o�@�_e\Ιٿ������@h�A% 4@�f ,4�!?/�D��o�@9����ٿ�Cg����@��Ot 4@c�?G�!?���o�@9����ٿ�Cg����@��Ot 4@c�?G�!?���o�@i�Oݙٿ�"�����@�Gr� 4@b�s0\�!?���o�@�E?���ٿ�վ���@1�]" 4@f�/p?�!?�g���o�@�¹��ٿ�;����@Z���% 4@���g�!?IR��o�@O���ٿ��l����@߉�# 4@���<�!?����o�@�W��ٿ&����@��7�* 4@ގ��ԏ!?FW�o�@!�l��ٿ������@���+6 4@���虏!?�d��o�@F�X�ٿ������@��@( 4@UQ&̑�!?�ì��o�@F�X�ٿ������@��@( 4@UQ&̑�!?�ì��o�@�A�԰�ٿ$�|����@P�_� 4@�9Oʏ!?��ܷ�o�@�A�԰�ٿ$�|����@P�_� 4@�9Oʏ!?��ܷ�o�@:����ٿ�!����@|�6 4@S��ȏ!?%>3��o�@:����ٿ�!����@|�6 4@S��ȏ!?%>3��o�@���Q��ٿ�ch����@l%i1 4@.�R���!?�oa��o�@�^k�əٿ�߼���@��( 4@�'a��!?gyh��o�@ a���ٿ�������@���	 4@�
��!?�����o�@q��㶙ٿ)�f����@KQ5 4@��d؏!?k��o�@q��㶙ٿ)�f����@KQ5 4@��d؏!?k��o�@z5�ϫ�ٿ>Y�����@nt:% 4@�=啳�!?�B��o�@O�řٿP�����@���. 4@��ke��!?����o�@����ݙٿ{[�����@��_v, 4@npc�!?B�ޣ�o�@�!ǝ��ٿA�$����@��;� 4@�@A;֏!?.j��o�@)����ٿ�������@{�V 4@}(yˏ!?uI���o�@��U�m�ٿ/Sǡ���@i	�E 4@�%5Ə!?�/��o�@*y�Dz�ٿKާ���@�&[E 4@鞥��!?�ص��o�@ٮ����ٿ������@�*f�
 4@�& Va�!?�Z7��o�@G��:�ٿ7������@/؈�. 4@LJ���!?/�'��o�@G��:�ٿ7������@/؈�. 4@LJ���!?/�'��o�@��'�ٿ��Ed���@&�lrL 4@����!?�v�k�o�@���_C�ٿ]��`���@d�ҭW 4@¹���!?�_jN�o�@���_C�ٿ]��`���@d�ҭW 4@¹���!?�_jN�o�@򷴫H�ٿ&�����@�i�O 4@��gf؏!?$dCb�o�@򷴫H�ٿ&�����@�i�O 4@��gf؏!?$dCb�o�@�]<�ٿo2n���@v��`L 4@`�����!?@�w�o�@3� �ٿ��}����@5}	/ 4@ڼ]֏!?\���o�@��L�ݙٿo\�����@���- 4@�;r��!?����o�@�gKS��ٿ��p���@�(w�5 4@#?7
{�!?l����o�@��c�ٿ	������@��o� 4@LWc��!?IJ���o�@g�#�ٿ2�cw���@+�A�7 4@�:ȟ�!?����o�@g�#�ٿ2�cw���@+�A�7 4@�:ȟ�!?����o�@_��+�ٿ�M#=���@��Q 4@	K�s�!?�
���o�@E۔p�ٿ��E���@[�Yr 4@��YЏ!?^�
��o�@�2^/x�ٿgF�����@��~ 4@> 	9�!?�����o�@�2^/x�ٿgF�����@��~ 4@> 	9�!?�����o�@���ٿ~������@�P|� 4@�� �!?;���o�@NZCO�ٿ��y$���@h,-�b 4@�Y[���!?.z���o�@u@c'�ٿ��F���@� V0 4@����!?��C�o�@u@c'�ٿ��F���@� V0 4@����!?��C�o�@u@c'�ٿ��F���@� V0 4@����!?��C�o�@-a�|�ٿ� ��@K���3@L!,�z�!?��ݙ�o�@-a�|�ٿ� ��@K���3@L!,�z�!?��ݙ�o�@A�][�ٿe~ ��@�����3@k��d��!?]����o�@|YǴv�ٿ��q���@ﳽ� 4@B���ԏ!??���o�@|YǴv�ٿ��q���@ﳽ� 4@B���ԏ!??���o�@�<|��ٿ������@��G��3@��RӅ�!?/"C�o�@��d�ٿ�;-U���@cI� 4@8��`�!?C�oZ�o�@�-D!�ٿ�潆���@c����3@p��c�!?�g�g�o�@�-D!�ٿ�潆���@c����3@p��c�!?�g�g�o�@��O�ٿCa�����@�� 4@��ݢ�!?I�5��o�@�&�!��ٿx(U~���@�)fV��3@�:�Z�!?4���o�@�&�!��ٿx(U~���@�)fV��3@�:�Z�!?4���o�@�4l��ٿ�x����@)xK�2 4@�+2q�!?��a��o�@�4l��ٿ�x����@)xK�2 4@�+2q�!?��a��o�@�4l��ٿ�x����@)xK�2 4@�+2q�!?��a��o�@�4l��ٿ�x����@)xK�2 4@�+2q�!?��a��o�@���+b�ٿI��:���@�M� 4@�Ӹ��!?.	��o�@���+b�ٿI��:���@�M� 4@�Ӹ��!?.	��o�@�`"ir�ٿWQ����@���5� 4@
\���!?���*�o�@�H��ٿ��!����@$�'�H 4@;R}�!?�:x��o�@�H��ٿ��!����@$�'�H 4@;R}�!?�:x��o�@�H��ٿ��!����@$�'�H 4@;R}�!?�:x��o�@�׿��ٿ`#�����@�"�yL 4@m�*���!?$V�8�o�@�׿��ٿ`#�����@�"�yL 4@m�*���!?$V�8�o�@����l�ٿ#Ɛ����@)=ٙP 4@��;V�!?;_4[�o�@R�ƚٿ�ǑC���@�U+.y 4@�ޱ��!?&�@r�o�@���|��ٿꯪ|���@ղ� 4@:�	6��!?�	�o�@�����ٿ�/|����@�	� 4@�>�ϐ�!?8����o�@W�~�ٿR0G���@�ؿ�j 4@
�`�e�!?v:���o�@W�~�ٿR0G���@�ؿ�j 4@
�`�e�!?v:���o�@f6Y	��ٿF�� ���@'/��S 4@r�+3��!?���i�o�@;��V�ٿl/SO���@�jn4 4@V�����!?J5�9�o�@;��V�ٿl/SO���@�jn4 4@V�����!?J5�9�o�@x�z�˘ٿ������@�2y"F 4@iq�7r�!?�� ��o�@x�z�˘ٿ������@�2y"F 4@iq�7r�!?�� ��o�@x�z�˘ٿ������@�2y"F 4@iq�7r�!?�� ��o�@���4�ٿN����@��B0� 4@�P�KЏ!? �0��o�@�<0ĩ�ٿ��JF���@�A?Kx4@E��y�!?�%w��o�@�<0ĩ�ٿ��JF���@�A?Kx4@E��y�!?�%w��o�@�
oY�ٿ#!6���@���� 4@����!?@�K��o�@��~�ٿ.P����@�gLv;4@"]WÏ!?S\L�o�@ɶ�%�ٿ��b4���@@o؈ 4@��\�Ǐ!?O��B�o�@ 09�ٿ;����@`v��� 4@��4WǏ!?.����o�@ 09�ٿ;����@`v��� 4@��4WǏ!?.����o�@��f���ٿc[���@�p� 4@��ʢ�!?�6���o�@_��8�ٿ�����@
���D 4@Yv�P��!?m݋��o�@_��8�ٿ�����@
���D 4@Yv�P��!?m݋��o�@��s^��ٿ��-���@�ܾ�  4@f�v#��!?�g�E�o�@;9ٜ��ٿA��� ��@�Z	n� 4@Ƙ���!?����o�@�QtM	�ٿh�� ��@�N�� 4@�\���!? հ��o�@:����ٿЩr����@����3@'V��!?QR̢�o�@�'�GV�ٿ������@��/ 4@���J��!?���	�o�@�'�GV�ٿ������@��/ 4@���J��!?���	�o�@�'�GV�ٿ������@��/ 4@���J��!?���	�o�@�'�GV�ٿ������@��/ 4@���J��!?���	�o�@�'�GV�ٿ������@��/ 4@���J��!?���	�o�@ڦۣ��ٿtPT����@����p 4@CnAƣ�!?#B��o�@�O�4��ٿ�ѸT���@Uk�X| 4@�{x���!?0���o�@�O�4��ٿ�ѸT���@Uk�X| 4@�{x���!?0���o�@�O�4��ٿ�ѸT���@Uk�X| 4@�{x���!?0���o�@@E��3�ٿ�N� ��@<\��4@�k��ԏ!?k�G*�o�@@E��3�ٿ�N� ��@<\��4@�k��ԏ!?k�G*�o�@@E��3�ٿ�N� ��@<\��4@�k��ԏ!?k�G*�o�@@E��3�ٿ�N� ��@<\��4@�k��ԏ!?k�G*�o�@@E��3�ٿ�N� ��@<\��4@�k��ԏ!?k�G*�o�@������ٿ�����@*t�P4@;"�z��!?$��o�@�JE�o�ٿ/",����@ (	��4@�PG���!?X
i��o�@����G�ٿ��.?���@5�;4@})�[��!?�W)��o�@��d;>�ٿz�>����@xB��� 4@]o[�\�!?g8��o�@��d;>�ٿz�>����@xB��� 4@]o[�\�!?g8��o�@��d;>�ٿz�>����@xB��� 4@]o[�\�!?g8��o�@�8�-��ٿopu����@��Ar 4@W��+`�!?J [�o�@�Ȼ��ٿ�{���@M
�[r�3@8F'��!?���p�@�Ȼ��ٿ�{���@M
�[r�3@8F'��!?���p�@�����ٿ��>����@'�*� 4@��=B�!?W��i�o�@�����ٿ��>����@'�*� 4@��=B�!?W��i�o�@�����ٿ��>����@'�*� 4@��=B�!?W��i�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@��;�/�ٿ��6q���@�+ۮ�3@A-�Џ!?B�3�o�@�	�d�ٿ��UZ��@v�=Ъ�3@J�1��!?(	Ld�o�@�	�d�ٿ��UZ��@v�=Ъ�3@J�1��!?(	Ld�o�@X&t�G�ٿTz{���@�]|c��3@u&ޏ!?t�1��o�@��͝ٿ(YR���@N��˻�3@�9����!?[�3�o�@��UN�ٿ�f�
��@+%��3@��-���!?6�|b�o�@��UN�ٿ�f�
��@+%��3@��-���!?6�|b�o�@����ٿ��RP��@�	(�e 4@B�qn��!?6���o�@� b�ٿ�ʕE��@�ja4�3@�
*r��!?yi*�o�@�k�e�ٿ�����@I.�d�3@���o�!?,��L�o�@��8֖ٿ������@���lZ�3@_�z��!?����o�@��8֖ٿ������@���lZ�3@_�z��!?����o�@��8֖ٿ������@���lZ�3@_�z��!?����o�@��8֖ٿ������@���lZ�3@_�z��!?����o�@&�3���ٿ�,}��@��I
��3@��z�!?m|c�o�@&�3���ٿ�,}��@��I
��3@��z�!?m|c�o�@SF�ٿ�{~����@���H4@9��x��!?ڵ*$�o�@�y�ٿx�����@�4@�M�ݏ!?�{��o�@�y�ٿx�����@�4@�M�ݏ!?�{��o�@;��9q�ٿ�g�
��@��
ΐ 4@��px�!?�����o�@;��9q�ٿ�g�
��@��
ΐ 4@��px�!?�����o�@;��9q�ٿ�g�
��@��
ΐ 4@��px�!?�����o�@;��9q�ٿ�g�
��@��
ΐ 4@��px�!?�����o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@�ӟ<A�ٿ�����@�˚�I4@�W9��!?��6�o�@j�-b�ٿ��U��@��� 4@��{ڨ�!?d8�o�@�Y�ٿ'$S���@�k��:4@�	<�w�!?�Iy�o�@�'^K�ٿ�R�_��@���� 4@RЏ�!?.�H_�o�@�:��ٿʰ����@��:��3@Ԇ�oޏ!?33� �o�@�:��ٿʰ����@��:��3@Ԇ�oޏ!?33� �o�@�:��ٿʰ����@��:��3@Ԇ�oޏ!?33� �o�@�:��ٿʰ����@��:��3@Ԇ�oޏ!?33� �o�@�:��ٿʰ����@��:��3@Ԇ�oޏ!?33� �o�@�*�E�ٿ��L�!��@�U8^2�3@y4r���!?��*�o�@�*�E�ٿ��L�!��@�U8^2�3@y4r���!?��*�o�@ә
�ٿ�1�x��@V��E 4@�:�!?ǅ��o�@x-�C5�ٿ�����@���_�3@B�+v!?69��o�@x-�C5�ٿ�����@���_�3@B�+v!?69��o�@x-�C5�ٿ�����@���_�3@B�+v!?69��o�@�3Ζ�ٿ��V>��@�;?��3@��֪�!?9�_$�o�@��S{�ٿ [(�&��@��N��4@�,�!?�gE��o�@��S{�ٿ [(�&��@��N��4@�,�!?�gE��o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�x`�Ԥٿ��s���@i�O��4@��+Ǐ!?7J�R�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@�=��6�ٿ�h���@.��4@ߕ+`ۏ!?v��X�o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@~���ٿlW5���@Y+w4 4@@��(̏!?I�F��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@����e�ٿ�h=��@ف�?��3@�L���!?͎��o�@!�t!��ٿ�b��@,�o'�3@H��!?�'��o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�	C4Ѩٿ��&�#��@�%l�]�3@ҫt���!?���w�o�@�NBx�ٿ�k=)��@�/`�<4@Z��؏!?�@P�o�@�NBx�ٿ�k=)��@�/`�<4@Z��؏!?�@P�o�@�NBx�ٿ�k=)��@�/`�<4@Z��؏!?�@P�o�@��?�Ӭٿ�w��@�GN�� 4@x�!?�ȸ�o�@�r�֜�ٿ�~���@G�# 4@��2�!?�G���o�@�r�֜�ٿ�~���@G�# 4@��2�!?�G���o�@:��9�ٿa���#��@�L��w4@<=���!?òĦo�@:��9�ٿa���#��@�L��w4@<=���!?òĦo�@:��9�ٿa���#��@�L��w4@<=���!?òĦo�@P����ٿ�R�P��@Q�O�%4@z�^駏!?n� ��o�@P����ٿ�R�P��@Q�O�%4@z�^駏!?n� ��o�@P����ٿ�R�P��@Q�O�%4@z�^駏!?n� ��o�@P����ٿ�R�P��@Q�O�%4@z�^駏!?n� ��o�@P����ٿ�R�P��@Q�O�%4@z�^駏!?n� ��o�@dbx��ٿ �Ӥ��@+��j4@�|�+��!?gg$��o�@dbx��ٿ �Ӥ��@+��j4@�|�+��!?gg$��o�@n��Q1�ٿ��:���@��x��4@':.֌�!?�\�o�@,:�"�ٿ�њK ��@�.�H 4@�6!?ٚ�y�o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@��b�Хٿ���	��@*V�� 4@{Ԃ���!?Ɖ���o�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@�U�E��ٿ�_�~���@�����4@�K9j�!?*�R�p�@A�;.��ٿ�l�M��@�����3@��z^�!?�ɨ p�@A�;.��ٿ�l�M��@�����3@��z^�!?�ɨ p�@A�;.��ٿ�l�M��@�����3@��z^�!?�ɨ p�@A�;.��ٿ�l�M��@�����3@��z^�!?�ɨ p�@P��Z��ٿ�I����@���N 4@q����!?�cJ)�o�@P��Z��ٿ�I����@���N 4@q����!?�cJ)�o�@��}�x�ٿ<W<���@Ru7��3@cZ����!?�i��o�@��}�x�ٿ<W<���@Ru7��3@cZ����!?�i��o�@��}�x�ٿ<W<���@Ru7��3@cZ����!?�i��o�@�1%�g�ٿ�#.�	��@�n��� 4@��[A�!?u�P&�o�@O�Y���ٿ�r�y��@��%��4@
��T�!?�ԏ<�o�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@u��-�ٿ�~n$��@���
�4@�8>�Ǐ!?�V͂Ao�@ؚ���ٿ������@��� 4@I}����!?��0�o�@ؚ���ٿ������@��� 4@I}����!?��0�o�@\o����ٿ�m��5��@���
 4@��-��!?�� go�@\o����ٿ�m��5��@���
 4@��-��!?�� go�@\o����ٿ�m��5��@���
 4@��-��!?�� go�@\o����ٿ�m��5��@���
 4@��-��!?�� go�@�`Z��ٿ�UO*��@@_ 4@sԱ�[�!?W��k5o�@�`Z��ٿ�UO*��@@_ 4@sԱ�[�!?W��k5o�@���#x�ٿ�s�T��@��Mn�3@����l�!?�����o�@���#x�ٿ�s�T��@��Mn�3@����l�!?�����o�@���#x�ٿ�s�T��@��Mn�3@����l�!?�����o�@�
��ٿ7��5��@�O�8�3@�="��!?�(W�n�@�
��ٿ7��5��@�O�8�3@�="��!?�(W�n�@�
��ٿ7��5��@�O�8�3@�="��!?�(W�n�@�
��ٿ7��5��@�O�8�3@�="��!?�(W�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@�y �ٿ)t}cZ��@�Z�O4@�F}���!?�y}�n�@fz�A�ٿ�*xt���@� �4@k%��!?��:>
l�@fz�A�ٿ�*xt���@� �4@k%��!?��:>
l�@fz�A�ٿ�*xt���@� �4@k%��!?��:>
l�@(��\��ٿ*�����@Jk�u�3@�G_V�!?$�nxl�@�VHA�ٿV�����@�/v@6�3@�ɺ�!?�_A�3k�@�VHA�ٿV�����@�/v@6�3@�ɺ�!?�_A�3k�@�VHA�ٿV�����@�/v@6�3@�ɺ�!?�_A�3k�@{��nq�ٿ�	����@H�� 4@����Տ!?p��qh�@{��nq�ٿ�	����@H�� 4@����Տ!?p��qh�@{��nq�ٿ�	����@H�� 4@����Տ!?p��qh�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@��SN:�ٿ �1*��@!8���4@�;�X��!?d���ce�@<�/_(�ٿ`*��@�F�w 4@g^Fb�!?IE��a�@<�/_(�ٿ`*��@�F�w 4@g^Fb�!?IE��a�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@)-�s�ٿ���yp��@r�%� 4@AtT]�!?�'^c�h�@b��Ξٿp8���@�F��� 4@�41��!?�D�inp�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@1��!"�ٿX$W����@_��3@� �W�!?��陵l�@>͒ࠪٿ	 ���@	In��3@*]��!?�#���z�@�1|��ٿU|�L��@�~�J� 4@`6j�d�!?�S3���@��Yy�ٿ !�D��@з�� 4@�:�Mۏ!?{ꏏ���@ZQ���ٿv|f����@�]���3@��?e��!?<��.��@k`�%�ٿ����Y��@��t{�3@Z>\��!?	O�Yn�@k`�%�ٿ����Y��@��t{�3@Z>\��!?	O�Yn�@k`�%�ٿ����Y��@��t{�3@Z>\��!?	O�Yn�@\~֒v�ٿ���e���@��� 4@��J�!?�40T/^�@�_���ٿ9�.5��@y��-4@�>�'�!?��hW�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@Ԉ?�Q�ٿ�˧�!��@�ӂ��4@��o�'�!?b�vKQ�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@���ٿF�$"���@DB4!� 4@��7u�!?.V@V�^�@B!��ٿ�ٓ]R��@�p=+�3@lV(�!?V8�K�@B!��ٿ�ٓ]R��@�p=+�3@lV(�!?V8�K�@cH�j}�ٿ��_�v��@��ϓ4@M�N��!?�,�zE�@�Sic�ٿ��ąc��@	d͇�3@[f���!?�gY�#�@�Sic�ٿ��ąc��@	d͇�3@[f���!?�gY�#�@�Sic�ٿ��ąc��@	d͇�3@[f���!?�gY�#�@�Sic�ٿ��ąc��@	d͇�3@[f���!?�gY�#�@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@0�■�ٿ�.�6D��@�����3@�6���!?�zR>��@;�PZڸٿ�(�O��@}ތ��3@w�,\�!?��<#��@��c���ٿ�� �v��@.���\4@?��L#�!?�?L����@:�G;Y�ٿT+�ۨ�@���*�3@��$Э�!?���9��@:�G;Y�ٿT+�ۨ�@���*�3@��$Э�!?���9��@:�G;Y�ٿT+�ۨ�@���*�3@��$Э�!?���9��@:�G;Y�ٿT+�ۨ�@���*�3@��$Э�!?���9��@s�Y�^�ٿ!��h��@�D/P�3@������!?u���@�@s�Y�^�ٿ!��h��@�D/P�3@������!?u���@�@s�Y�^�ٿ!��h��@�D/P�3@������!?u���@�@�	9��ٿ�1Ƹ��@1&2�24@�Ӽ�`�!?�_�v�@�%�lT�ٿ���Wa��@��Ė��3@) 0tu�!?Y�N�|'�@�%�lT�ٿ���Wa��@��Ė��3@) 0tu�!?Y�N�|'�@�%�lT�ٿ���Wa��@��Ė��3@) 0tu�!?Y�N�|'�@�%�lT�ٿ���Wa��@��Ė��3@) 0tu�!?Y�N�|'�@�%�lT�ٿ���Wa��@��Ė��3@) 0tu�!?Y�N�|'�@����ٿ�&1���@I�^ 4@'i쨍�!?:-�|�b�@����ٿ�&1���@I�^ 4@'i쨍�!?:-�|�b�@����ٿ�&1���@I�^ 4@'i쨍�!?:-�|�b�@����ٿ�&1���@I�^ 4@'i쨍�!?:-�|�b�@����ٿ�&1���@I�^ 4@'i쨍�!?:-�|�b�@��p�:�ٿ�!y���@���4�3@����܎!?ԝX�{��@��p�:�ٿ�!y���@���4�3@����܎!?ԝX�{��@�m�#��ٿZ�����@	�y 4@}0*�ʏ!?�q�����@��1:/�ٿ��r���@$� 4@-ٚ�Ə!?_�3���@��1:/�ٿ��r���@$� 4@-ٚ�Ə!?_�3���@��1:/�ٿ��r���@$� 4@-ٚ�Ə!?_�3���@��1:/�ٿ��r���@$� 4@-ٚ�Ə!?_�3���@��1:/�ٿ��r���@$� 4@-ٚ�Ə!?_�3���@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@#�gQ�ٿ�v�,J(�@��A�3@�<D�!?��J�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@Y�7 �ٿc��)��@�l�, 4@�/���!?6K�P�@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@`���ٿ:�ـ���@�I4���3@E���ȏ!?�I��k��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@�;�̩ٿ	�^�J��@�w�� 4@M��i��!?�k�v��@��-:�ٿ��"�@y0z^4@f�~��!?�v�j�@��N�,�ٿ,��x"!�@��1��3@�����!?66	�tn�@��N�,�ٿ,��x"!�@��1��3@�����!?66	�tn�@��N�,�ٿ,��x"!�@��1��3@�����!?66	�tn�@��N�,�ٿ,��x"!�@��1��3@�����!?66	�tn�@�l~P �ٿ��O����@�W�4@J[s��!?���%��@�l~P �ٿ��O����@�W�4@J[s��!?���%��@�l~P �ٿ��O����@�W�4@J[s��!?���%��@�l~P �ٿ��O����@�W�4@J[s��!?���%��@�l~P �ٿ��O����@�W�4@J[s��!?���%��@�}p�z�ٿe�����@�V�4@��'��!?���zk��@�}p�z�ٿe�����@�V�4@��'��!?���zk��@�}p�z�ٿe�����@�V�4@��'��!?���zk��@�}p�z�ٿe�����@�V�4@��'��!?���zk��@�}p�z�ٿe�����@�V�4@��'��!?���zk��@:��!��ٿ���e'�@�Y�u4@n&N�m�!?2��c
�@:��!��ٿ���e'�@�Y�u4@n&N�m�!?2��c
�@�H��	�ٿq�v���@��]�-4@�5�,�!?��-N��@�H��	�ٿq�v���@��]�-4@�5�,�!?��-N��@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@TXm׉�ٿӒ����@�I[�4@�x��!?��Xt~�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@���	�ٿPt~��@W�f�d4@�g�̏!?���7\�@\��V�ٿ��t ��@�M9\{ 4@`W�8Џ!?�əS)�@0T�Z�ٿ�}� ���@@N�q 4@�,��@�!?6��^�$�@0T�Z�ٿ�}� ���@@N�q 4@�,��@�!?6��^�$�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@zĶ+��ٿ~։����@j��� 4@;G���!?L�au4�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@������ٿ��߂���@V��"	4@����!?R�zBD�@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@G{[A��ٿt�-���@Eh��m 4@��dI��!?\=���@6K�ٿT�<���@��j���3@�̀w�!?���/�@��2�2�ٿ}�S`��@��^f|�3@�����!?ѭl��1�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@���&��ٿ�q/���@�7V���3@�\��ŏ!?��9U�)�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Bj�ٿf~����@����3@���|�!?�?��"3�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@��Ik�ٿ�F�@;^���4@���9��!?��7*�@٣����ٿ����;
�@/+� 4@wz�X�!?g=�إ��@�l�؛�ٿo�� $��@�Y��4@���d�!?߰$�}�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@՝9�ٿ��~]��@�em 4@�!�Ğ�!?���~�J�@���áٿ6y�}�@���Y��3@���we�!?�Z�s���@�y����ٿ�[�@�8p��3@�h9�!?�I�ͮ�@� nߣٿ�l%u��@`�q;��3@,��}(�!?�����@� nߣٿ�l%u��@`�q;��3@,��}(�!?�����@� nߣٿ�l%u��@`�q;��3@,��}(�!?�����@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@E���ٿW�ۨ��@y�o4@&6XJ�!?�ي �@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@ݢ'*�ٿ���]���@�+�� 4@?�5I�!?Mt�=�$�@<�f���ٿ>U2���@eh[F$4@N��zs�!?���M ��@B��ٿ��8����@'��9�4@��Ԓ�!?֎���@�=��Ϧٿ�`�l���@�h�a}4@�2�붏!?���d$��@�=��Ϧٿ�`�l���@�h�a}4@�2�붏!?���d$��@�=��Ϧٿ�`�l���@�h�a}4@�2�붏!?���d$��@�7�1t�ٿ[�gR�@�پB<4@��<�q�!?��n'#��@�7�1t�ٿ[�gR�@�پB<4@��<�q�!?��n'#��@�7�1t�ٿ[�gR�@�پB<4@��<�q�!?��n'#��@��_lY�ٿ��T���@X?� 4@�w�p��!?aң>'Q�@��_lY�ٿ��T���@X?� 4@�w�p��!?aң>'Q�@��_lY�ٿ��T���@X?� 4@�w�p��!?aң>'Q�@��_lY�ٿ��T���@X?� 4@�w�p��!?aң>'Q�@��_lY�ٿ��T���@X?� 4@�w�p��!?aң>'Q�@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@���A[�ٿ���f��@��c~D4@�-5p�!?�ӭ��@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@T��͢ٿc3�����@W*�)[4@��Ua�!?o���BG�@W��Qͧٿ4��h���@s<��4@��/W�!?<��s/�@W��Qͧٿ4��h���@s<��4@��/W�!?<��s/�@W��Qͧٿ4��h���@s<��4@��/W�!?<��s/�@W��Qͧٿ4��h���@s<��4@��/W�!?<��s/�@W��Qͧٿ4��h���@s<��4@��/W�!?<��s/�@_'ƨٿ�BO���@tF��4@�M���!?�2�]��@(��f�ٿ�۶����@��Fl4@�ތ��!?���m�@(��f�ٿ�۶����@��Fl4@�ތ��!?���m�@(��f�ٿ�۶����@��Fl4@�ތ��!?���m�@a�Vf�ٿ��2���@d�f!4@p/?��!?i+�+�\�@a�Vf�ٿ��2���@d�f!4@p/?��!?i+�+�\�@�%�\�ٿ�����@�Zs4@$��0Џ!?�W%2�P�@i��@��ٿakEr�@d�k4@58�!?���M��@i��@��ٿakEr�@d�k4@58�!?���M��@�5Q*"�ٿ���I��@d���4@�o���!?�Ӓ,��@�5Q*"�ٿ���I��@d���4@�o���!?�Ӓ,��@�5Q*"�ٿ���I��@d���4@�o���!?�Ӓ,��@v~�ٿ8᜕�
�@^���^4@�&z�!?��o)��@v~�ٿ8᜕�
�@^���^4@�&z�!?��o)��@v~�ٿ8᜕�
�@^���^4@�&z�!?��o)��@u����ٿ������@��F�4@,@�_ҏ!?����X�@u����ٿ������@��F�4@,@�_ҏ!?����X�@u����ٿ������@��F�4@,@�_ҏ!?����X�@u����ٿ������@��F�4@,@�_ҏ!?����X�@'��5�ٿ���-���@!/���3@IK���!?F4��X�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@���e{�ٿL�O���@xU�B4@��2���!?\k�*U3�@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@�����ٿ*e����@�=�I�4@/����!?�V����@[fL�9�ٿ�_�%_��@6�D4@ŭ�7��!?)���/;�@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@�S��z�ٿr�S��@�E��4@���?}�!?'W�	��@9���"�ٿU+��g��@49�\ 4@��t���!?<�㧸�@5Mf�ޚٿo3~�z��@�M&� 4@,�p�ď!?�s�&��@5Mf�ޚٿo3~�z��@�M&� 4@,�p�ď!?�s�&��@Ac�a�ٿ���!,�@Ԏ��4@���ď!?�vO�	�@Ac�a�ٿ���!,�@Ԏ��4@���ď!?�vO�	�@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@j.���ٿ��#X�@���Z 4@1�E���!?$��0��@���c�ٿ�ۿ�J��@(�dr� 4@����!?}b#�h��@���c�ٿ�ۿ�J��@(�dr� 4@����!?}b#�h��@��g<�ٿ2�v���@j���|�3@�%��x�!?�Z@���@��g<�ٿ2�v���@j���|�3@�%��x�!?�Z@���@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@ɛ��ٿ�3Lw���@�ů�n�3@E��!?��b�)�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@�R 	�ٿ>ʣ'���@��x��3@Ɩb��!?��/p�@T 'A�ٿW��t;	�@�+D%4@����!?o�����@T 'A�ٿW��t;	�@�+D%4@����!?o�����@T 'A�ٿW��t;	�@�+D%4@����!?o�����@T 'A�ٿW��t;	�@�+D%4@����!?o�����@T 'A�ٿW��t;	�@�+D%4@����!?o�����@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@� /�F�ٿ�ʄ���@#P��4@�u���!?.@RHF�@��3���ٿ/y,���@:��'� 4@qid,��!?��)���@2LA5o�ٿ��'�q��@�<Z�� 4@L�{E�!?֥�j91�@��W��ٿ��|���@.<��4@Vm(��!?�~���@����ٿ}�����@P}��x 4@��2Y��!?_�nQ�H�@����ٿ}�����@P}��x 4@��2Y��!?_�nQ�H�@�Pujߕٿ�|�YT��@:�T��3@�CNÏ!?�&+c#��@t�f��ٿ���'���@�!�"�4@�A��e�!?v�Ӝ�]�@t�f��ٿ���'���@�!�"�4@�A��e�!?v�Ӝ�]�@t�f��ٿ���'���@�!�"�4@�A��e�!?v�Ӝ�]�@t�f��ٿ���'���@�!�"�4@�A��e�!?v�Ӝ�]�@t�f��ٿ���'���@�!�"�4@�A��e�!?v�Ӝ�]�@���%5�ٿ�=(�"��@����4@R
^�!?����ԑ�@�{/�k�ٿK���_�@���И4@�Asz�!?���,��@�{/�k�ٿK���_�@���И4@�Asz�!?���,��@Un4���ٿr�ǋ���@uћ4@J�5���!?<�P�b�@Un4���ٿr�ǋ���@uћ4@J�5���!?<�P�b�@Un4���ٿr�ǋ���@uћ4@J�5���!?<�P�b�@Un4���ٿr�ǋ���@uћ4@J�5���!?<�P�b�@�A�V��ٿvCS� �@_�DX� 4@�w���!?N�!W�@�A�V��ٿvCS� �@_�DX� 4@�w���!?N�!W�@�A�V��ٿvCS� �@_�DX� 4@�w���!?N�!W�@�A�V��ٿvCS� �@_�DX� 4@�w���!?N�!W�@�A�V��ٿvCS� �@_�DX� 4@�w���!?N�!W�@> �
�ٿ豓���@
5MZ4@V0nզ�!?9�:�u�@�=��ٿ�2����@3�, 4@p�Zڏ!?�9ݳ�V�@�=��ٿ�2����@3�, 4@p�Zڏ!?�9ݳ�V�@��Q�ٿ�l����@����K�3@ ]���!?h��{G�@��Q�ٿ�l����@����K�3@ ]���!?h��{G�@��Q�ٿ�l����@����K�3@ ]���!?h��{G�@��Q�ٿ�l����@����K�3@ ]���!?h��{G�@�Y���ٿ�͎F��@4F���4@Yȓ��!?�s��_�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@��	�l�ٿ��)�9�@��2H�4@q�S��!?�N�\�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@]�>��ٿ���8��@��U4@�-��!?��_"�<�@QDZAßٿ}�~{8
�@Y���Y 4@�[f��!?7��'���@QDZAßٿ}�~{8
�@Y���Y 4@�[f��!?7��'���@QDZAßٿ}�~{8
�@Y���Y 4@�[f��!?7��'���@QDZAßٿ}�~{8
�@Y���Y 4@�[f��!?7��'���@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@bj*R�ٿk��{	 �@%I4@`�� ��!?\�3��@������ٿC
�=�@�E�� 4@��j)��!?R//���@������ٿC
�=�@�E�� 4@��j)��!?R//���@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@,��@6�ٿV��[�@�Ⱦ�4@�D���!?��`)�@!T�KY�ٿҦ�R�@x��-4@��2Z�!?b�ӡ��@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@lh=��ٿ0�A�D�@x8�4@�3�雏!?�����@tD�5��ٿ0��Q��@({%�4@x ��7�!?�:�k0$�@tD�5��ٿ0��Q��@({%�4@x ��7�!?�:�k0$�@tD�5��ٿ0��Q��@({%�4@x ��7�!?�:�k0$�@
,����ٿ��R���@.�T�4@���-�!?��O�P�@
,����ٿ��R���@.�T�4@���-�!?��O�P�@
,����ٿ��R���@.�T�4@���-�!?��O�P�@
,����ٿ��R���@.�T�4@���-�!?��O�P�@	��w�ٿ"3*Y�@�߸9�4@Ht8��!?�.tG��@	��w�ٿ"3*Y�@�߸9�4@Ht8��!?�.tG��@	��w�ٿ"3*Y�@�߸9�4@Ht8��!?�.tG��@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@�.�ц�ٿ�{R	���@�%�9��3@�a�3�!?[Ũ�e,�@[̃3^�ٿf1�t'��@�����4@�{֚��!?�����$�@[̃3^�ٿf1�t'��@�����4@�{֚��!?�����$�@�
	�b�ٿ�b�=�@��4@=�ó�!?J�Sb��@.In�?�ٿ���b��@c,x\4@KyRt�!?}EO�I�@.In�?�ٿ���b��@c,x\4@KyRt�!?}EO�I�@.In�?�ٿ���b��@c,x\4@KyRt�!?}EO�I�@.In�?�ٿ���b��@c,x\4@KyRt�!?}EO�I�@.In�?�ٿ���b��@c,x\4@KyRt�!?}EO�I�@g���ٿ~�~mO��@�!�/�4@8��ۏ!?,���3�@�$�4��ٿ	�/]��@ ?����3@?��n�!?S�f+M�@����ͫٿ�T�\��@r5��` 4@�=v͏!?leͨ��@����ͫٿ�T�\��@r5��` 4@�=v͏!?leͨ��@����ͫٿ�T�\��@r5��` 4@�=v͏!?leͨ��@����ͫٿ�T�\��@r5��` 4@�=v͏!?leͨ��@pL`H��ٿ��4���@��P���3@�/�C��!?�}HQ�@pL`H��ٿ��4���@��P���3@�/�C��!?�}HQ�@pL`H��ٿ��4���@��P���3@�/�C��!?�}HQ�@ɨ�T�ٿ��J9k��@��k��4@��1��!?�
(��J�@ɨ�T�ٿ��J9k��@��k��4@��1��!?�
(��J�@ɨ�T�ٿ��J9k��@��k��4@��1��!?�
(��J�@�Lu�ߢٿ�ھi5�@&/���3@�I�)z�!?�����@�Lu�ߢٿ�ھi5�@&/���3@�I�)z�!?�����@�Lu�ߢٿ�ھi5�@&/���3@�I�)z�!?�����@�}ĥ*�ٿ���W�@�$
#Y�3@1�*M�!?�2u��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@�����ٿ�2���@퉡l 4@2Z��!?�Ͽa��@��F胠ٿT�
{���@�+����3@0ߨ ��!?�%,�R"�@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@��
��ٿ�y��O	�@���B 4@CY⊏!?h��}��@�53�9�ٿ��h=��@y��d�4@�6��f�!?�NE���@�53�9�ٿ��h=��@y��d�4@�6��f�!?�NE���@�53�9�ٿ��h=��@y��d�4@�6��f�!?�NE���@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@K���ٿ]��1���@q��l�4@Hּym�!?$��SK�@���6�ٿCLW��@�ˮ�� 4@ג)1~�!?����@���6�ٿCLW��@�ˮ�� 4@ג)1~�!?����@�S���ٿER^��@�]6���3@��̰�!?������@�S���ٿER^��@�]6���3@��̰�!?������@H+�τ�ٿ�}7��@���~ 4@����ޏ!?i�w��@H+�τ�ٿ�}7��@���~ 4@����ޏ!?i�w��@H+�τ�ٿ�}7��@���~ 4@����ޏ!?i�w��@H+�τ�ٿ�}7��@���~ 4@����ޏ!?i�w��@H+�τ�ٿ�}7��@���~ 4@����ޏ!?i�w��@�����ٿj��g�@@���3@3�|q��!?ϐ,����@�FK7��ٿ��O���@ ���3@�38��!?�����@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@g����ٿ�?\����@�f�4@N�6�!?D(ùjX�@*i���ٿ�����@\�� 4@RG�q��!?
w:�Js�@*i���ٿ�����@\�� 4@RG�q��!?
w:�Js�@"-$]۬ٿu�.���@��~k�3@dS�!?����@"-$]۬ٿu�.���@��~k�3@dS�!?����@�4͒��ٿ��a{"�@���3��3@�#z��!?�װ�޻�@���%�ٿ)Cx��@z�C/ 4@;�a"��!?�^���@���%�ٿ)Cx��@z�C/ 4@;�a"��!?�^���@[��� �ٿ������@r=B��3@m���!?�4JhP�@[��� �ٿ������@r=B��3@m���!?�4JhP�@[��� �ٿ������@r=B��3@m���!?�4JhP�@[��� �ٿ������@r=B��3@m���!?�4JhP�@��أ�ٿ�����@�Vfg 4@z�K��!?�@���@��أ�ٿ�����@�Vfg 4@z�K��!?�@���@x�ѓ��ٿ!6�2a��@o((��3@_>󊵏!?�y{hL�@x�ѓ��ٿ!6�2a��@o((��3@_>󊵏!?�y{hL�@x�ѓ��ٿ!6�2a��@o((��3@_>󊵏!?�y{hL�@x�ѓ��ٿ!6�2a��@o((��3@_>󊵏!?�y{hL�@~�7D�ٿ���9�"�@�#
�4@ݭ�u�!?�ևs^|�@~�7D�ٿ���9�"�@�#
�4@ݭ�u�!?�ևs^|�@~�7D�ٿ���9�"�@�#
�4@ݭ�u�!?�ևs^|�@~�7D�ٿ���9�"�@�#
�4@ݭ�u�!?�ևs^|�@���ٿ�(8��@0#L�4@�@HQx�!?[��yE�@���ٿ�(8��@0#L�4@�@HQx�!?[��yE�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@`~O��ٿ}���@�u��� 4@�D��!?	_��J0�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@�����ٿ�&�%���@p��X
 4@Z�'��!?�ܺ��^�@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@$P���ٿ@"B;��@U�1�� 4@(��٧�!? ���K��@U�.�!�ٿ����[��@��� 4@�l,z��!?�';��@�H���ٿB�g �@�y��4@7�%��!?�|��+�@�H���ٿB�g �@�y��4@7�%��!?�|��+�@�H���ٿB�g �@�y��4@7�%��!?�|��+�@�H���ٿB�g �@�y��4@7�%��!?�|��+�@���[�ٿ�B=^v�@0� 4@P�o���!?&�\���@���[�ٿ�B=^v�@0� 4@P�o���!?&�\���@�I ۃ�ٿMs���@C�	� 4@�~�%x�!?�[m�|�@�I ۃ�ٿMs���@C�	� 4@�~�%x�!?�[m�|�@�I ۃ�ٿMs���@C�	� 4@�~�%x�!?�[m�|�@�I ۃ�ٿMs���@C�	� 4@�~�%x�!?�[m�|�@�&wͅ�ٿ���Pg��@��fo� 4@�]��C�!?,��'��@�&wͅ�ٿ���Pg��@��fo� 4@�]��C�!?,��'��@�&wͅ�ٿ���Pg��@��fo� 4@�]��C�!?,��'��@�&wͅ�ٿ���Pg��@��fo� 4@�]��C�!?,��'��@ߏ4��ٿ�g ��@L3����3@��vWK�!?`{�ܩ��@ߏ4��ٿ�g ��@L3����3@��vWK�!?`{�ܩ��@kn��@�ٿ�$_����@p�� 4@�p�}8�!?����@kn��@�ٿ�$_����@p�� 4@�p�}8�!?����@kn��@�ٿ�$_����@p�� 4@�p�}8�!?����@z�ǧ�ٿ�b'x��@i�ܗR4@=(�U�!?��z9"�@z�ǧ�ٿ�b'x��@i�ܗR4@=(�U�!?��z9"�@����ٿVV$�?��@ud9'��3@��r�ˏ!?��å��@����ٿVV$�?��@ud9'��3@��r�ˏ!?��å��@����ٿVV$�?��@ud9'��3@��r�ˏ!?��å��@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@�hw�ٿL\p6W�@]�@�9 4@�G��ŏ!?������@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@��?�<�ٿ�<m���@1�t��3@��@x��!?��3�4�@�,s��ٿ�1�/�@���4@����Џ!?����'��@�,s��ٿ�1�/�@���4@����Џ!?����'��@�,s��ٿ�1�/�@���4@����Џ!?����'��@�,s��ٿ�1�/�@���4@����Џ!?����'��@�,s��ٿ�1�/�@���4@����Џ!?����'��@�mS�ٿ#�{��@#3��� 4@?�
���!?E}�UlI�@�mS�ٿ#�{��@#3��� 4@?�
���!?E}�UlI�@�mS�ٿ#�{��@#3��� 4@?�
���!?E}�UlI�@�mS�ٿ#�{��@#3��� 4@?�
���!?E}�UlI�@��ZלٿI<���@�x`u=4@/	��ڏ!?#��H&�@;�b�t�ٿ�aA�P��@���� 4@=��	M�!?Oۥ���@;�b�t�ٿ�aA�P��@���� 4@=��	M�!?Oۥ���@;�b�t�ٿ�aA�P��@���� 4@=��	M�!?Oۥ���@�r�m.�ٿ0v���@oV�Q� 4@@�nt�!?Ǥ����@�r�m.�ٿ0v���@oV�Q� 4@@�nt�!?Ǥ����@�r�m.�ٿ0v���@oV�Q� 4@@�nt�!?Ǥ����@�r�m.�ٿ0v���@oV�Q� 4@@�nt�!?Ǥ����@�r�m.�ٿ0v���@oV�Q� 4@@�nt�!?Ǥ����@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@��?�J�ٿ�u��V��@��m~I�3@�����!?�F���%�@���2��ٿ��._H��@�,x 4@3ԩF�!?��Z�9�@���2��ٿ��._H��@�,x 4@3ԩF�!?��Z�9�@���2��ٿ��._H��@�,x 4@3ԩF�!?��Z�9�@���2��ٿ��._H��@�,x 4@3ԩF�!?��Z�9�@�|�R�ٿ~���@��+��4@R_ ~0�!?�����@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@IZ�ۿ�ٿ�>N�7�@#��D&4@�f�!?��ʙ�@2+&�<�ٿ�Jq��@d�
�� 4@����!?9R#eT��@U�m��ٿ�KT���@�Wp(� 4@�+��ڏ!?��� �@U�m��ٿ�KT���@�Wp(� 4@�+��ڏ!?��� �@U�m��ٿ�KT���@�Wp(� 4@�+��ڏ!?��� �@U�m��ٿ�KT���@�Wp(� 4@�+��ڏ!?��� �@�����ٿ,eUo��@��Dw 4@��q��!?��@XS��@�����ٿ,eUo��@��Dw 4@��q��!?��@XS��@�����ٿ,eUo��@��Dw 4@��q��!?��@XS��@�����ٿ,eUo��@��Dw 4@��q��!?��@XS��@�����ٿ,eUo��@��Dw 4@��q��!?��@XS��@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@���D�ٿ7v%��@=��\x4@ξ-���!?���]�@]��c>�ٿ��U)���@L��^� 4@�a]R�!?�2��e�@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@��ٿ@Ȃ,��@��W�Y4@�̥_��!?Ѽ�0��@x�_F�ٿR���^9�@^�o��4@h��ш�!?m{�>��@x�_F�ٿR���^9�@^�o��4@h��ш�!?m{�>��@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@��<��ٿ�Ĵ�@*NP�3@@�:��!?���X���@`{�ߡٿ��FF��@���Q�3@G�8��!?��W��0�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@W�����ٿ1V����@�m� 4@�;k֏!?�[	�$�@Pk���ٿ������@���4@�U��|�!? B�
�I�@Pk���ٿ������@���4@�U��|�!? B�
�I�@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@���]�ٿn�y����@�J�Vy4@�����!?���f��@�!+�e�ٿ�C]+���@F��M4@~�ޏ!?>���5�@�!+�e�ٿ�C]+���@F��M4@~�ޏ!?>���5�@,��k�ٿW������@4���4@,���!?�9�: f�@b����ٿ�8X��	�@�ح"�4@N���{�!?-�7�T�@b����ٿ�8X��	�@�ح"�4@N���{�!?-�7�T�@�&�ٿ�1���@��iG�4@_�a�<�!?� �W[E�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@܂M7��ٿs<��8�@�n�ĉ 4@`rM��!?_P^�FC�@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@��Nt��ٿ��9l� �@{b<�3@��v���!?�����@ͪ�ݚٿe�C���@�h,�3@|^7��!?��;����@ͪ�ݚٿe�C���@�h,�3@|^7��!?��;����@�C�XH�ٿK������@���8�3@������!?�}��|X�@�C�XH�ٿK������@���8�3@������!?�}��|X�@�C�XH�ٿK������@���8�3@������!?�}��|X�@���N�ٿ����ʶ�@��
�' 4@�Ab��!?�&����@���N�ٿ����ʶ�@��
�' 4@�Ab��!?�&����@t����ٿ�P�����@��n��3@.��ˏ!?�\4�g��@��˩��ٿ�G���m�@"I3x�4@Z\�.��!? �<8�@��˩��ٿ�G���m�@"I3x�4@Z\�.��!? �<8�@��i>[�ٿ���e�@����= 4@��M5�!?����@��i>[�ٿ���e�@����= 4@��M5�!?����@��i>[�ٿ���e�@����= 4@��M5�!?����@��i>[�ٿ���e�@����= 4@��M5�!?����@���2�ٿ�L2y���@x�/�3@א�E?�!?[W�hA�@���2�ٿ�L2y���@x�/�3@א�E?�!?[W�hA�@w��ٿ������@�p�Ç�3@�Ǩ�"�!?ps�C3��@w��ٿ������@�p�Ç�3@�Ǩ�"�!?ps�C3��@w��ٿ������@�p�Ç�3@�Ǩ�"�!?ps�C3��@w��ٿ������@�p�Ç�3@�Ǩ�"�!?ps�C3��@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@i��F˥ٿ2u���@�}G#2�3@����!?�0e���@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@ıN���ٿ>0 ��*�@��)�� 4@6�q-��!?/  ��@8��=�ٿ�+��e�@'q�F�4@&���ď!?���w���@8��=�ٿ�+��e�@'q�F�4@&���ď!?���w���@8��=�ٿ�+��e�@'q�F�4@&���ď!?���w���@8��=�ٿ�+��e�@'q�F�4@&���ď!?���w���@(�`�ٿ����n��@�f�4@Pg4�F�!?-mG` �@(�`�ٿ����n��@�f�4@Pg4�F�!?-mG` �@(�`�ٿ����n��@�f�4@Pg4�F�!?-mG` �@(�`�ٿ����n��@�f�4@Pg4�F�!?-mG` �@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@��	�ٿe���Hb�@�����3@�S%}�!?2v��@6@���ٿ�3�Z���@ �@�	�3@���2�!?�u�6m�@d����ٿ��]�^�@ \�Y �3@5?W&�!?�$.<��@d����ٿ��]�^�@ \�Y �3@5?W&�!?�$.<��@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@П�Zڟٿ��6Wd�@|�O,�3@G�D��!?������@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@���	�ٿc2�B��@�:� � 4@s�gh��!?����}��@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@ٝ��ٿ3ΏXf�@6����3@�}@Lm�!?�ՙ�r5�@vHIƠٿt��L9��@ICY]� 4@���5��!?8L/�H�@vHIƠٿt��L9��@ICY]� 4@���5��!?8L/�H�@vHIƠٿt��L9��@ICY]� 4@���5��!?8L/�H�@�k6E�ٿF���@�����3@'+Oڷ�!?��gn���@�k6E�ٿF���@�����3@'+Oڷ�!?��gn���@�k6E�ٿF���@�����3@'+Oڷ�!?��gn���@�k6E�ٿF���@�����3@'+Oڷ�!?��gn���@�k6E�ٿF���@�����3@'+Oڷ�!?��gn���@����ٿ2N�ib��@M�����3@ڥ}�Ώ!?�^P�	��@����ٿ2N�ib��@M�����3@ڥ}�Ώ!?�^P�	��@����ٿ2N�ib��@M�����3@ڥ}�Ώ!?�^P�	��@;��*��ٿ0J�&��@����3@ȍ򚮏!?Dn%Wm�@;��*��ٿ0J�&��@����3@ȍ򚮏!?Dn%Wm�@;��*��ٿ0J�&��@����3@ȍ򚮏!?Dn%Wm�@;��*��ٿ0J�&��@����3@ȍ򚮏!?Dn%Wm�@� �_Ğٿ������@rd�l�4@�H�2��!?�N��@� �_Ğٿ������@rd�l�4@�H�2��!?�N��@� �_Ğٿ������@rd�l�4@�H�2��!?�N��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@�	��V�ٿl��^�Q�@v�{v��3@]��z��!?7�n�l��@p=�f��ٿ:����@k�W�4@}e
G��!?t�$�C�@p=�f��ٿ:����@k�W�4@}e
G��!?t�$�C�@p �J/�ٿ%� ���@��<�V 4@f��މ�!?0]c�g��@p �J/�ٿ%� ���@��<�V 4@f��މ�!?0]c�g��@p �J/�ٿ%� ���@��<�V 4@f��މ�!?0]c�g��@p �J/�ٿ%� ���@��<�V 4@f��މ�!?0]c�g��@p �J/�ٿ%� ���@��<�V 4@f��މ�!?0]c�g��@-���E�ٿ����.�@��4@G5�^�!?c뙒UK�@-���E�ٿ����.�@��4@G5�^�!?c뙒UK�@7�>�|�ٿ��KM��@x�(�7 4@����!?�\�X��@7�>�|�ٿ��KM��@x�(�7 4@����!?�\�X��@7�>�|�ٿ��KM��@x�(�7 4@����!?�\�X��@7�>�|�ٿ��KM��@x�(�7 4@����!?�\�X��@7�>�|�ٿ��KM��@x�(�7 4@����!?�\�X��@�Y�Ɗ�ٿ*�[0D�@�H7o� 4@B�<��!?��9�4t�@�Y�Ɗ�ٿ*�[0D�@�H7o� 4@B�<��!?��9�4t�@�Y�Ɗ�ٿ*�[0D�@�H7o� 4@B�<��!?��9�4t�@�Լ�ٿH�)L��@�W�94@+��4Ï!?LEBYl�@�Լ�ٿH�)L��@�W�94@+��4Ï!?LEBYl�@�Լ�ٿH�)L��@�W�94@+��4Ï!?LEBYl�@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@ڮ<�V�ٿ�[�,s��@n7�T 4@eM"
��!?R�D@,��@��}�l�ٿ���{��@+ѽ' 4@��ɏ!?�y�jδ�@��}�l�ٿ���{��@+ѽ' 4@��ɏ!?�y�jδ�@��}�l�ٿ���{��@+ѽ' 4@��ɏ!?�y�jδ�@��}�l�ٿ���{��@+ѽ' 4@��ɏ!?�y�jδ�@єmy�ٿ���be|�@dx�4@��&_i�!?�������@єmy�ٿ���be|�@dx�4@��&_i�!?�������@єmy�ٿ���be|�@dx�4@��&_i�!?�������@,q�ߣٿ-<)!@��@{�i��3@.Zԙ��!?Çq�
�@,q�ߣٿ-<)!@��@{�i��3@.Zԙ��!?Çq�
�@,q�ߣٿ-<)!@��@{�i��3@.Zԙ��!?Çq�
�@,q�ߣٿ-<)!@��@{�i��3@.Zԙ��!?Çq�
�@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�q��ٿS�ȡgy�@>H9@ 4@��v���!?�����@�e�rT�ٿt��B\��@BN� 4@)����!?�Ծh��@�e�rT�ٿt��B\��@BN� 4@)����!?�Ծh��@�e�rT�ٿt��B\��@BN� 4@)����!?�Ծh��@�e�rT�ٿt��B\��@BN� 4@)����!?�Ծh��@�e�rT�ٿt��B\��@BN� 4@)����!?�Ծh��@Cқ�ٿ��z��@��>� 4@'q��!?�_�0eA�@Cқ�ٿ��z��@��>� 4@'q��!?�_�0eA�@Cқ�ٿ��z��@��>� 4@'q��!?�_�0eA�@Cқ�ٿ��z��@��>� 4@'q��!?�_�0eA�@Cқ�ٿ��z��@��>� 4@'q��!?�_�0eA�@���7�ٿ%3����@�`+4@�8�w��!?t���*�@���7�ٿ%3����@�`+4@�8�w��!?t���*�@=��3�ٿ	� ���@p�K4@�q윏!?f��'���@=��3�ٿ	� ���@p�K4@�q윏!?f��'���@��㑄�ٿx����@�d�.4@��	��!?���"Z��@��2�ٿ���@��/�7 4@B����!?�]s�@o�xi�ٿ����/|�@O���4@3�{��!?j�)�?L�@�f�c�ٿ��^��z�@�p�4@�����!?~xEU���@�f�c�ٿ��^��z�@�p�4@�����!?~xEU���@�f�c�ٿ��^��z�@�p�4@�����!?~xEU���@��{{6�ٿ��F��@u�>z|�3@�n���!?d%���2�@��{{6�ٿ��F��@u�>z|�3@�n���!?d%���2�@�M���ٿa�N��<�@�7��_�3@�C� ��!?�8;�i�@�M���ٿa�N��<�@�7��_�3@�C� ��!?�8;�i�@�M���ٿa�N��<�@�7��_�3@�C� ��!?�8;�i�@�M���ٿa�N��<�@�7��_�3@�C� ��!?�8;�i�@k�-%k�ٿ�`�c�@�n9���3@,��b�!?�]^��@�%)�Ɲٿ�j}��@��}��3@�Q�0��!?�_3
�@�%)�Ɲٿ�j}��@��}��3@�Q�0��!?�_3
�@�%)�Ɲٿ�j}��@��}��3@�Q�0��!?�_3
�@�%)�Ɲٿ�j}��@��}��3@�Q�0��!?�_3
�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@T����ٿxf� ��@M�A�4@��4��!?N��!5�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@c*�1�ٿ���CE��@�P����3@3.�M��!?�Ȳ�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@Q`U��ٿ��{����@�u="� 4@�r񠢏!?}ĺ�B�@"��@�ٿ��GCD�@��NV� 4@�q͚�!?ￖΞZ�@"��@�ٿ��GCD�@��NV� 4@�q͚�!?ￖΞZ�@?�alݤٿ7�ͫ��@9RZi�3@����x�!?���}�@?�alݤٿ7�ͫ��@9RZi�3@����x�!?���}�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@VhLJ�ٿD�h�P�@��Q�; 4@���lw�!?�\�a�J�@���|�ٿ�9�Ėw�@!y����3@ܸVK��!?,��5��@���|�ٿ�9�Ėw�@!y����3@ܸVK��!?,��5��@7�7��ٿܧ¶$��@�G$�E 4@���Տ!?#R���@7�7��ٿܧ¶$��@�G$�E 4@���Տ!?#R���@7�7��ٿܧ¶$��@�G$�E 4@���Տ!?#R���@7�7��ٿܧ¶$��@�G$�E 4@���Տ!?#R���@7�7��ٿܧ¶$��@�G$�E 4@���Տ!?#R���@ )Ly�ٿbsg��@�F�� 4@Ĵ��Ə!?�� �K�@�jW�ٿ��@I���@����|4@��IH��!?����@{Ӳ��ٿa����@H�h��4@}�\��!?U���P��@{Ӳ��ٿa����@H�h��4@}�\��!?U���P��@{Ӳ��ٿa����@H�h��4@}�\��!?U���P��@`�
]��ٿ�HX�b�@,��A�3@ڻ��ߏ!?	x~o�'�@`�
]��ٿ�HX�b�@,��A�3@ڻ��ߏ!?	x~o�'�@�����ٿ����@��� 4@�K<�Ə!?�j}��)�@�����ٿ����@��� 4@�K<�Ə!?�j}��)�@s�d3��ٿ�d����@?Y�X��3@��˟ԏ!?S����@>`�~�ٿ9��1�e�@��~W 4@A֝UЏ!?�R�U$!�@>`�~�ٿ9��1�e�@��~W 4@A֝UЏ!?�R�U$!�@>`�~�ٿ9��1�e�@��~W 4@A֝UЏ!?�R�U$!�@>`�~�ٿ9��1�e�@��~W 4@A֝UЏ!?�R�U$!�@�!�:��ٿ�|Nt��@&�����3@�>(���!?&{i��`�@�!�:��ٿ�|Nt��@&�����3@�>(���!?&{i��`�@����ٿ�$dDD�@���3@W�Fʏ!?%s��8�@P{W&�ٿXd]���@ �c���3@��p��!?t�dݢ�@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@ب�H��ٿطwu��@(�TJ@�3@ʁ�ō�!?��߉���@�Nb
ˮٿ/w�>��@w�	\��3@��|CM�!?h��=60�@�Nb
ˮٿ/w�>��@w�	\��3@��|CM�!?h��=60�@݆}�z�ٿ�,dN4&�@��ި� 4@]{� L�!?�����@݆}�z�ٿ�,dN4&�@��ި� 4@]{� L�!?�����@E �a�ٿ���-�h�@cf����3@��n$�!?��H 6~�@E �a�ٿ���-�h�@cf����3@��n$�!?��H 6~�@E �a�ٿ���-�h�@cf����3@��n$�!?��H 6~�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@��U��ٿ'YTus��@�|��3@s�E���!?N3�}�@F��ՠٿU��ƍu�@g�,y 4@��ȏ!?��4���@F��ՠٿU��ƍu�@g�,y 4@��ȏ!?��4���@F��ՠٿU��ƍu�@g�,y 4@��ȏ!?��4���@F��ՠٿU��ƍu�@g�,y 4@��ȏ!?��4���@�/Рٿ%��ݏ�@ �Y���3@�L� ��!?���r��@�/Рٿ%��ݏ�@ �Y���3@�L� ��!?���r��@��u��ٿ{I� ��@�H�zu4@�PA͏!?K�${�@��u��ٿ{I� ��@�H�zu4@�PA͏!?K�${�@��u��ٿ{I� ��@�H�zu4@�PA͏!?K�${�@��u��ٿ{I� ��@�H�zu4@�PA͏!?K�${�@A����ٿ�C��r��@�7�տ�3@6Թ��!?|h���@A����ٿ�C��r��@�7�տ�3@6Թ��!?|h���@A����ٿ�C��r��@�7�տ�3@6Թ��!?|h���@A����ٿ�C��r��@�7�տ�3@6Թ��!?|h���@���$��ٿ�]IW���@zyc�� 4@��D�!?ۥ�ƚ�@	�k��ٿ�0`!��@���� 4@���c��!?G~\�G��@	�k��ٿ�0`!��@���� 4@���c��!?G~\�G��@	�k��ٿ�0`!��@���� 4@���c��!?G~\�G��@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@jο���ٿU�PIFY�@s���4@!>Ed��!?� | =�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@o<sHïٿ�o����@R��{�4@O��ȓ�!?��X�'�@�n[��ٿ%f`w ��@�S(և4@?�5���!?�X����@�n[��ٿ%f`w ��@�S(և4@?�5���!?�X����@�n[��ٿ%f`w ��@�S(և4@?�5���!?�X����@�n[��ٿ%f`w ��@�S(և4@?�5���!?�X����@�n[��ٿ%f`w ��@�S(և4@?�5���!?�X����@:�5��ٿ�e/���@Eo4@\�(uՏ!?�<�2���@:�5��ٿ�e/���@Eo4@\�(uՏ!?�<�2���@:�5��ٿ�e/���@Eo4@\�(uՏ!?�<�2���@:�5��ٿ�e/���@Eo4@\�(uՏ!?�<�2���@:�5��ٿ�e/���@Eo4@\�(uՏ!?�<�2���@.�0{̬ٿ+uEi�h�@�'��>4@Su
��!?��<Q��@, ���ٿ�Q�0�@i��4@90pr�!?�4}¤�@, ���ٿ�Q�0�@i��4@90pr�!?�4}¤�@�cV�ٿ�-��@�$YP�4@�߾�c�!?{��	�<�@|P39��ٿ������@�|�4@�^*5y�!?܁�S���@|P39��ٿ������@�|�4@�^*5y�!?܁�S���@�h��s�ٿ��<t��@3�D$� 4@F��#��!?Y��\���@`��`�ٿ��f�0G�@X]���4@]^�a��!?��_�O(�@�q,D�ٿ���\��@~�T���3@��MV �!?!ӿM;�@�q,D�ٿ���\��@~�T���3@��MV �!?!ӿM;�@�q,D�ٿ���\��@~�T���3@��MV �!?!ӿM;�@���;��ٿ[� �D��@~��3@�D�:L�!?�RAu�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@m�����ٿ���M�@�=�| 4@���r�!?�����v�@�c�T�ٿ_�n����@J)�c� 4@{U�*n�!?E�kj�;�@�c�T�ٿ_�n����@J)�c� 4@{U�*n�!?E�kj�;�@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@���O�ٿs����Q�@�~Go��3@-�Y�g�!?I��c@��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@R?f�F�ٿ����?��@�ݤ���3@����!?�"�]��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@�~�P��ٿ+�M����@�9�!��3@�A�м�!?��I�_��@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@������ٿv@�PH�@�ۀ�2 4@
D�ڣ�!?t��$�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@�nD�қٿn�$jXG�@��I��3@�>�w�!?�O��מ�@ػ���ٿ�n�\|A�@�Br�!�3@��3m��!?OR�`��@ػ���ٿ�n�\|A�@�Br�!�3@��3m��!?OR�`��@�\"���ٿ�r����@�:�3�3@����e�!?�4�5��@�%@դٿ�Vh���@*)79\�3@��J�!?�0���@�%@դٿ�Vh���@*)79\�3@��J�!?�0���@@�v(�ٿ�!o�m~�@�V���3@h���K�!?�N�H*��@���[��ٿx��N*�@��]R� 4@�p�:��!?2��ɗ�@���[��ٿx��N*�@��]R� 4@�p�:��!?2��ɗ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@��3��ٿ$�ȭf��@�?�Q4@d�Ï!?�D�3ڈ�@�8�yN�ٿ�����@�iy�� 4@�j�ҏ!?#���@�8�yN�ٿ�����@�iy�� 4@�j�ҏ!?#���@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�=P畑ٿbc��!u�@;�=� 4@�;���!?�3	R��@�K�e��ٿ��
W��@m�<�4@e��p��!?�^d�@�K�e��ٿ��
W��@m�<�4@e��p��!?�^d�@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@��+�ٿ�f7`;�@E�o[4@$r�Ï!?\%Q���@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@#��nB�ٿ7�46Z�@�5��� 4@}�`E^�!?���(7�@Y,�㲦ٿCay�@-5�JS4@ќ!-�!?���_��@Y,�㲦ٿCay�@-5�JS4@ќ!-�!?���_��@�$�ٿ\\�W�@� �e'4@�U�#0�!?š}��@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@SP�P�ٿ^��P���@4���4@���n�!?����i�@ֽ�Z�ٿ�&��*�@軒���3@Q �A�!?v��v<�@ֽ�Z�ٿ�&��*�@軒���3@Q �A�!?v��v<�@ֽ�Z�ٿ�&��*�@軒���3@Q �A�!?v��v<�@ֽ�Z�ٿ�&��*�@軒���3@Q �A�!?v��v<�@v.�&�ٿ������@̦�$��3@6g�!?q����d�@^���z�ٿ���j�/�@t�|zB�3@W��x��!?g����@^���z�ٿ���j�/�@t�|zB�3@W��x��!?g����@�
3�ٿ�m>�e��@�+ɤ14@3+�j�!?j������@�
3�ٿ�m>�e��@�+ɤ14@3+�j�!?j������@�
3�ٿ�m>�e��@�+ɤ14@3+�j�!?j������@�
3�ٿ�m>�e��@�+ɤ14@3+�j�!?j������@�
3�ٿ�m>�e��@�+ɤ14@3+�j�!?j������@�\��.�ٿ�4�V<�@��^.�4@T{X��!?���h��@�\��.�ٿ�4�V<�@��^.�4@T{X��!?���h��@�\��.�ٿ�4�V<�@��^.�4@T{X��!?���h��@�\��.�ٿ�4�V<�@��^.�4@T{X��!?���h��@�\��.�ٿ�4�V<�@��^.�4@T{X��!?���h��@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@��糡ٿ�������@Q�
�� 4@+�i�F�!?�+͠8�@�RI��ٿhµ�{�@^�801 4@�M��O�!?D�"����@�RI��ٿhµ�{�@^�801 4@�M��O�!?D�"����@�RI��ٿhµ�{�@^�801 4@�M��O�!?D�"����@�RI��ٿhµ�{�@^�801 4@�M��O�!?D�"����@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@�R�-g�ٿ�����@��T84@G��/�!?��
l&�@P���S�ٿ9��j+Z�@�1k4@����!?Y:C�ƀ�@P���S�ٿ9��j+Z�@�1k4@����!?Y:C�ƀ�@P���S�ٿ9��j+Z�@�1k4@����!?Y:C�ƀ�@P���S�ٿ9��j+Z�@�1k4@����!?Y:C�ƀ�@:�R$U�ٿ{�v�%��@�zU�3@��=@��!?x�!'�6�@bdi#��ٿ��^F�@��ěk�3@�����!?9�j����@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@+G�W��ٿ�_Ǆ�r�@0���S 4@�!rϏ!?�F��%3�@��g��ٿ1����G�@lN! 4@L0
6Ə!? �xI]�@��g��ٿ1����G�@lN! 4@L0
6Ə!? �xI]�@��g��ٿ1����G�@lN! 4@L0
6Ə!? �xI]�@��g��ٿ1����G�@lN! 4@L0
6Ə!? �xI]�@��g��ٿ1����G�@lN! 4@L0
6Ə!? �xI]�@:A���ٿ)i�3��@��Қ� 4@��l��!?�)�����@:A���ٿ)i�3��@��Қ� 4@��l��!?�)�����@:A���ٿ)i�3��@��Қ� 4@��l��!?�)�����@:A���ٿ)i�3��@��Қ� 4@��l��!?�)�����@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@�V��`�ٿV�DD��@Nxvg� 4@A@=�U�!?��e��@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@ܤ�`��ٿ�j,����@���A 4@��ϸX�!?���Ix�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@���d�ٿm�ug�g�@ U��3@�8�"�!?p�K�ϣ�@�Ρ��ٿ��.G\��@���h 4@`��!?(�|���@�Ρ��ٿ��.G\��@���h 4@`��!?(�|���@Qw�'$�ٿ���ji��@�*�� 4@H��̏!?����@Qw�'$�ٿ���ji��@�*�� 4@H��̏!?����@�~ MU�ٿ�J%�@��>���3@� q��!?�T��|��@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@v;�G֚ٿ�=cҤ�@Xu�4@����!?+������@\$9'�ٿb&�[/�@f���� 4@�Cmn��!?䢒��r�@\$9'�ٿb&�[/�@f���� 4@�Cmn��!?䢒��r�@\$9'�ٿb&�[/�@f���� 4@�Cmn��!?䢒��r�@\$9'�ٿb&�[/�@f���� 4@�Cmn��!?䢒��r�@\$9'�ٿb&�[/�@f���� 4@�Cmn��!?䢒��r�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�耲�ٿ���q�@��M��3@)�`
��!?�Ic�U�@�O� �ٿUZ)'���@[Lc��3@�К�k�!?��[�ʦ�@�xVU�ٿ�C�e��@Ƴ��3@�D���!?�T�����@�xVU�ٿ�C�e��@Ƴ��3@�D���!?�T�����@�xVU�ٿ�C�e��@Ƴ��3@�D���!?�T�����@�xVU�ٿ�C�e��@Ƴ��3@�D���!?�T�����@�xVU�ٿ�C�e��@Ƴ��3@�D���!?�T�����@T���ٿz�[�"�@�p����3@���я!?鐲��L�@T���ٿz�[�"�@�p����3@���я!?鐲��L�@T���ٿz�[�"�@�p����3@���я!?鐲��L�@Lt"��ٿ���>H��@c �#4@�˯���!?j�l�v�@Lt"��ٿ���>H��@c �#4@�˯���!?j�l�v�@� X�s�ٿ���k��@��f 4@��w:k�!?Ս����@� X�s�ٿ���k��@��f 4@��w:k�!?Ս����@� X�s�ٿ���k��@��f 4@��w:k�!?Ս����@� X�s�ٿ���k��@��f 4@��w:k�!?Ս����@p���"�ٿ�&��p�@���F4@�xs��!??�2S��@�̇ղ�ٿ4%<9�5�@eL�)O4@y��gҏ!?��] �@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@���D��ٿaԊ�@��@�V�O64@���d�!?y^{���@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@�*
\�ٿ���Y���@渐ѥ 4@�1ʏ��!?_����@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Y�����ٿA��z�@�] �A4@Zх�Ə!?�/yO���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@Uv~{6�ٿ�;��{�@^�F�� 4@�_2�!?��_���@��"v6�ٿ��d�,*�@�����3@@���W�!?��b����@��"v6�ٿ��d�,*�@�����3@@���W�!?��b����@��"v6�ٿ��d�,*�@�����3@@���W�!?��b����@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@��ǡ�ٿ0
+��*�@����W�3@9���я!?	���$�@�|o��ٿcڻ��(�@�����4@�<&�!?��}t&R�@�8˧ٿ�̕�@���bT�3@;��!��!?��6���@�8˧ٿ�̕�@���bT�3@;��!��!?��6���@�8˧ٿ�̕�@���bT�3@;��!��!?��6���@�8˧ٿ�̕�@���bT�3@;��!��!?��6���@�8˧ٿ�̕�@���bT�3@;��!��!?��6���@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@}P����ٿ��K�7?�@��[�a 4@ �䕚�!?V�:-+��@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�ջ#�ٿ�Ak(O|�@�$��3@���͏!?��)�3�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�WΥٿ5Ym�Z�@�C��4@�߯͏!?�G%c�o�@�g�ٿ� ��#�@t�j:4@�;��w�!?x#�g1
�@�g�ٿ� ��#�@t�j:4@�;��w�!?x#�g1
�@N�r2�ٿ���B�_�@%w�- 4@*��O�!?\�����@N�r2�ٿ���B�_�@%w�- 4@*��O�!?\�����@N�r2�ٿ���B�_�@%w�- 4@*��O�!?\�����@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@&qȇ�ٿo�Z���@�=n�p�3@��@ҏ!?�J�|;V�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@��Kq�ٿ���}��@Z�ʧ��3@e&�3L�!?g�֫IU�@;NW���ٿn������@F`A� 4@���ŏ�!?
��a���@;NW���ٿn������@F`A� 4@���ŏ�!?
��a���@x���ٿ��	T��@)��r��3@�����!?3wo��@x���ٿ��	T��@)��r��3@�����!?3wo��@x���ٿ��	T��@)��r��3@�����!?3wo��@x���ٿ��	T��@)��r��3@�����!?3wo��@jŰ�ٿ�
�+�@�+�;4@L�#�!?������@jŰ�ٿ�
�+�@�+�;4@L�#�!?������@jŰ�ٿ�
�+�@�+�;4@L�#�!?������@jŰ�ٿ�
�+�@�+�;4@L�#�!?������@��w��ٿJ�K����@tG 4@�ˏ!?H�J����@��w��ٿJ�K����@tG 4@�ˏ!?H�J����@_�4�ãٿX�"�P�@IڮdX4@����l�!?�|�k��@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�cΚ~�ٿ��_�}r�@�f����3@]^7j�!?��O���@�!3�ٿ��3o	��@��S�4@i���m�!?a������@�!3�ٿ��3o	��@��S�4@i���m�!?a������@�!3�ٿ��3o	��@��S�4@i���m�!?a������@�!3�ٿ��3o	��@��S�4@i���m�!?a������@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�8�菟ٿ�p��+��@���U�4@�Ɇ�l�!?�獢�@�(��ٿ�����@�n�4@׭��@�!?|�Dr��@�(��ٿ�����@�n�4@׭��@�!?|�Dr��@�(��ٿ�����@�n�4@׭��@�!?|�Dr��@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@GEM*s�ٿ\d��D�@9]��4@����e�!?�,����@2�GI�ٿ��.m��@���� 4@�r=^��!?W����@2�GI�ٿ��.m��@���� 4@�r=^��!?W����@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@38︔ٿ�2�����@H�� 4@��3��!?<2�n1d�@��
�ٿT�_R�@�mK'��3@�V�$s�!?����@��
�ٿT�_R�@�mK'��3@�V�$s�!?����@��
�ٿT�_R�@�mK'��3@�V�$s�!?����@��
�ٿT�_R�@�mK'��3@�V�$s�!?����@��
�ٿT�_R�@�mK'��3@�V�$s�!?����@���ͥٿ���w(��@&5#�4@)�Ѵ��!?�����@���ͥٿ���w(��@&5#�4@)�Ѵ��!?�����@���ͥٿ���w(��@&5#�4@)�Ѵ��!?�����@���ͥٿ���w(��@&5#�4@)�Ѵ��!?�����@���ٿ�����@}�PM64@e��ҏ!?���*�@���ٿ�����@}�PM64@e��ҏ!?���*�@���ٿ�����@}�PM64@e��ҏ!?���*�@���ٿ�����@}�PM64@e��ҏ!?���*�@���ٿ�����@}�PM64@e��ҏ!?���*�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@޷��0�ٿ�J[�`�@O���l 4@L�7��!?�4��m�@g��YA�ٿAgxٶ��@��UE��3@�,q�ߏ!?2{�92�@g��YA�ٿAgxٶ��@��UE��3@�,q�ߏ!?2{�92�@g��YA�ٿAgxٶ��@��UE��3@�,q�ߏ!?2{�92�@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@_-�$U�ٿI{+�]�@�A�� 4@�����!?�{}���@�x��ٿ������@�>@*s4@p"��W�!?����n�@),E
��ٿ��}��r�@MCC[� 4@4y���!?�O�w���@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@�r�&ޡٿT� �� �@��{�4@6�r�R�!?e��n��@r�����ٿX�v���@9���s�3@�]�t��!?F4	Md��@r�����ٿX�v���@9���s�3@�]�t��!?F4	Md��@r�����ٿX�v���@9���s�3@�]�t��!?F4	Md��@r�����ٿX�v���@9���s�3@�]�t��!?F4	Md��@r�����ٿX�v���@9���s�3@�]�t��!?F4	Md��@�ɛ�?�ٿF9��}�@'ۜ�4@p�g=�!?�}@�l��@�ɛ�?�ٿF9��}�@'ۜ�4@p�g=�!?�}@�l��@�ɛ�?�ٿF9��}�@'ۜ�4@p�g=�!?�}@�l��@�L�w��ٿ*��6�;�@3=6pg�3@�SE~�!?��[(��@�L�w��ٿ*��6�;�@3=6pg�3@�SE~�!?��[(��@�l����ٿ*��*R�@9�Q�3@��Ǐ!?�����@��
��ٿ_�8A��@1f�4@c���ҏ!?���Ņr�@��
��ٿ_�8A��@1f�4@c���ҏ!?���Ņr�@��
��ٿ_�8A��@1f�4@c���ҏ!?���Ņr�@��
��ٿ_�8A��@1f�4@c���ҏ!?���Ņr�@�Ȱ��ٿ=q`4���@C�;ڭ�3@V��ex�!?��u��@��$��ٿ��kT�2�@Q�q��3@�T��l�!?n�O�@��$��ٿ��kT�2�@Q�q��3@�T��l�!?n�O�@��$��ٿ��kT�2�@Q�q��3@�T��l�!?n�O�@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@�}�ʨٿ�ؾ���@o��[p 4@*��ޭ�!?�N_c$��@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@���Z�ٿ]@�Y���@#Hu!� 4@�� Ǐ!??|����@S����ٿ��#Kj�@��\�4@^���!?��;�@S����ٿ��#Kj�@��\�4@^���!?��;�@S����ٿ��#Kj�@��\�4@^���!?��;�@'���}�ٿ��3�C�@���Õ4@sT�Q֏!?E���w�@'���}�ٿ��3�C�@���Õ4@sT�Q֏!?E���w�@'���}�ٿ��3�C�@���Õ4@sT�Q֏!?E���w�@�h	�G�ٿ=hb	W�@n��8-4@�~�u��!?�z�b�y�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�&Өr�ٿ}3:,���@��y 4@����!?�j�KF�@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@�]�2��ٿ�u�Ǒ��@�ar�6 4@2�	Z��!?	�Mf��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@���äٿ�Og���@��e�� 4@��J���!?w�Fn��@eӼٿ��Wwb�@~6
1��3@gY��!?���C��@eӼٿ��Wwb�@~6
1��3@gY��!?���C��@sj73�ٿ}>&Շe�@~�=iG�3@��n�ӏ!?���-g��@sj73�ٿ}>&Շe�@~�=iG�3@��n�ӏ!?���-g��@sj73�ٿ}>&Շe�@~�=iG�3@��n�ӏ!?���-g��@sj73�ٿ}>&Շe�@~�=iG�3@��n�ӏ!?���-g��@I;$��ٿ�J��M�@!��;��3@U}�R�!?������@%B�T6�ٿ.7�J�S�@\�$7� 4@�o����!?Tk�/���@%B�T6�ٿ.7�J�S�@\�$7� 4@�o����!?Tk�/���@%B�T6�ٿ.7�J�S�@\�$7� 4@�o����!?Tk�/���@%B�T6�ٿ.7�J�S�@\�$7� 4@�o����!?Tk�/���@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@�P���ٿ������@���3@�3G��!?2��y�@!`y�ٿ��|��@
�L]�3@
�����!?�G�R(!�@���ϟٿ��:����@9F=x>�3@��=�֏!?���4�=�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@9$�唙ٿ��i:��@�0���3@$(��Џ!?��Cf�@{���ٿ������@N��f� 4@��Q�!?�&�op��@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@�TpƬ�ٿi�%n,��@vRҚ� 4@��eZ�!?�cU����@0��Ťٿ�v�d���@�ߑ0 4@���%�!?�E%��@�UE�ٿ뺨��@�]�4@!봂��!?��V���@�UE�ٿ뺨��@�]�4@!봂��!?��V���@�UE�ٿ뺨��@�]�4@!봂��!?��V���@�UE�ٿ뺨��@�]�4@!봂��!?��V���@�UE�ٿ뺨��@�]�4@!봂��!?��V���@�UE�ٿ뺨��@�]�4@!봂��!?��V���@������ٿ��`}�@t��K4@���H�!?3��pt�@������ٿ��`}�@t��K4@���H�!?3��pt�@������ٿ��`}�@t��K4@���H�!?3��pt�@������ٿ��`}�@t��K4@���H�!?3��pt�@L�+H�ٿ)�F)B��@䰙��4@�S�`o�!?
⊙��@L�+H�ٿ)�F)B��@䰙��4@�S�`o�!?
⊙��@L�+H�ٿ)�F)B��@䰙��4@�S�`o�!?
⊙��@L�+H�ٿ)�F)B��@䰙��4@�S�`o�!?
⊙��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@�"�z�ٿ�$�9p�@�xry� 4@*epIݏ!?!6:j��@<�Q��ٿ"�s�P��@Ȳ\��4@�����!?�`(�o�@<�Q��ٿ"�s�P��@Ȳ\��4@�����!?�`(�o�@ߨ;p^�ٿ�H 1�7�@�T䜝 4@�T�G�!?Xg�Q�@�a ���ٿ}�޵*�@Pj 4@r!��ɏ!?��&
�@~$g[�ٿA���$��@ة��3@�+���!?��Ѩ�6�@~$g[�ٿA���$��@ة��3@�+���!?��Ѩ�6�@~$g[�ٿA���$��@ة��3@�+���!?��Ѩ�6�@��F���ٿQ������@�J٨�3@6�n��!?"�8���@��F���ٿQ������@�J٨�3@6�n��!?"�8���@��F���ٿQ������@�J٨�3@6�n��!?"�8���@�t�q�ٿ�~.,��@�!��3@�}W��!?E�Ttб�@�t�q�ٿ�~.,��@�!��3@�}W��!?E�Ttб�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@�h!:�ٿ q�e���@Y]�xx 4@���!?�hon�Z�@����n�ٿo�]Tz�@;z#�=�3@�j~U��!?Fk�.�@����n�ٿo�]Tz�@;z#�=�3@�j~U��!?Fk�.�@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@����K�ٿ���%g��@.HJ�I4@s�-��!?��T��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@&�A�ٿV>ȓ�U�@�k
���3@ç1���!?ct�Ŭ��@f�l;��ٿ����5�@ �~��3@�P�Di�!?���V���@f�l;��ٿ����5�@ �~��3@�P�Di�!?���V���@f�l;��ٿ����5�@ �~��3@�P�Di�!?���V���@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@��?^��ٿAaJOL�@�]"� 4@����c�!?��N�2��@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@
����ٿB~��O��@$o�4@<�#��!?��?a�@n��m�ٿYf��2��@��۸4@ͤ�;��!?�
V�;e�@�%f�ٿ?�w���@ѕSQ4@��d�!?��c�@�%f�ٿ?�w���@ѕSQ4@��d�!?��c�@�%f�ٿ?�w���@ѕSQ4@��d�!?��c�@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���{��ٿfݡGg@�@.�]q/ 4@Ut��!?;�L��@���!�ٿ�G#PU�@��� 4@�����!?�8�-�@���!�ٿ�G#PU�@��� 4@�����!?�8�-�@���!�ٿ�G#PU�@��� 4@�����!?�8�-�@��f�H�ٿ8eQe��@�B/�4@v`���!?��M$�2�@��f�H�ٿ8eQe��@�B/�4@v`���!?��M$�2�@��f�H�ٿ8eQe��@�B/�4@v`���!?��M$�2�@��f�H�ٿ8eQe��@�B/�4@v`���!?��M$�2�@̶���ٿ���5�@M��c�4@62�y�!?/0�#7�@�MV��ٿ#��%��@4��|b4@�PŀG�!?DlAi��@>���,�ٿunܸ���@т2JM4@��3��!?z�37�@>���,�ٿunܸ���@т2JM4@��3��!?z�37�@>���,�ٿunܸ���@т2JM4@��3��!?z�37�@>���,�ٿunܸ���@т2JM4@��3��!?z�37�@R!R���ٿ��#����@~�]��4@�x��!?�S.KA�@R!R���ٿ��#����@~�]��4@�x��!?�S.KA�@R!R���ٿ��#����@~�]��4@�x��!?�S.KA�@R!R���ٿ��#����@~�]��4@�x��!?�S.KA�@R!R���ٿ��#����@~�]��4@�x��!?�S.KA�@���N�ٿ�v���#�@}NL��3@�iiB��!?���k�@���N�ٿ�v���#�@}NL��3@�iiB��!?���k�@�	I
!�ٿf9��x=�@U�P���3@�]�}��!?��o��@Q�b8�ٿڇD�k��@5��g� 4@{$C��!?k1R���@��d`�ٿ�$E�ڀ�@�~d��3@������!?I�@���@��d`�ٿ�$E�ڀ�@�~d��3@������!?I�@���@c�'�ʥٿ_7ޫ��@�b�ܹ 4@�C�U�!?@*56��@c�'�ʥٿ_7ޫ��@�b�ܹ 4@�C�U�!?@*56��@c�'�ʥٿ_7ޫ��@�b�ܹ 4@�C�U�!?@*56��@
xzA�ٿn��S&�@���\�4@�ؠ��!?��~���@
xzA�ٿn��S&�@���\�4@�ؠ��!?��~���@��L�ۢٿ7�����@�ыb4@ ?�}Q�!?	�&Y�@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@�����ٿ��_SR-�@a$�h4@�TQ'Ə!?�6�_��@9d�>Δٿ {���@�<1Q 4@��.g��!?�ɾ�x�@9d�>Δٿ {���@�<1Q 4@��.g��!?�ɾ�x�@9d�>Δٿ {���@�<1Q 4@��.g��!?�ɾ�x�@9d�>Δٿ {���@�<1Q 4@��.g��!?�ɾ�x�@Ì��ٿt@�jF�@�'^ 4@̣"{c�!?�����7�@Ì��ٿt@�jF�@�'^ 4@̣"{c�!?�����7�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@����ܛٿ��T��h�@"�ܮv4@2�`��!?�Vc��,�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@uO�F�ٿ4=����@�(�4@8�ھ��!?��j3�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@�Yi�ٿ�]Gco��@*�R4o4@@Ȃ���!?J�;:;�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��b*��ٿQB�5�x�@i�g�4@��yɤ�!?��Q�@��A�ٿ���Zq�@m��� 4@���nя!?%�Vmi��@��A�ٿ���Zq�@m��� 4@���nя!?%�Vmi��@q�-㘫ٿ�8��~�@ ��a� 4@脹�ď!?�s���@q�-㘫ٿ�8��~�@ ��a� 4@脹�ď!?�s���@q�-㘫ٿ�8��~�@ ��a� 4@脹�ď!?�s���@q�-㘫ٿ�8��~�@ ��a� 4@脹�ď!?�s���@����ٿ��ŗ��@%8� ��3@I�ی_�!?5o�π�@�c��éٿ��z;}��@�s�{�3@��DN!�!?��!E�@��V,ƭٿ��k�_�@��G64@7����!?��;����@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@��Yҧٿ[��u���@p�x�Y4@�H�Y�!?��l��@D���ٿ��'�5P�@7_Y�.4@Ʋ!*֏!? ��خ��@D���ٿ��'�5P�@7_Y�.4@Ʋ!*֏!? ��خ��@D���ٿ��'�5P�@7_Y�.4@Ʋ!*֏!? ��خ��@D���ٿ��'�5P�@7_Y�.4@Ʋ!*֏!? ��خ��@�h����ٿ�\�y&��@Mw����3@]�F׷�!?O!\u�P�@LUOȀ�ٿ�D����@�zw�3@u�j�!?#<�3>��@LUOȀ�ٿ�D����@�zw�3@u�j�!?#<�3>��@N}q+�ٿ�&��Y��@��7n|�3@^��ʏ!?�W���@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@�6(`��ٿ6�3�`5�@ĳ�I4@�R-}r�!?va��h�@h�D�ٿ�Lh��@���4@E���l�!?
A|��l�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@t�ٿ��t�ER�@��D5` 4@� �&��!?sm%@�@R��M��ٿ��hɀB�@*[���4@�	���!?0���|m�@R��M��ٿ��hɀB�@*[���4@�	���!?0���|m�@R��M��ٿ��hɀB�@*[���4@�	���!?0���|m�@R��M��ٿ��hɀB�@*[���4@�	���!?0���|m�@R��M��ٿ��hɀB�@*[���4@�	���!?0���|m�@�����ٿ�8���@(+���3@��2��!?L:B���@p) �ٿ}I4����@>�.M��3@�����!?D���n�@�>�U�ٿ�L��=~�@e���64@�?mM}�!?��z&*�@�>�U�ٿ�L��=~�@e���64@�?mM}�!?��z&*�@�&��r�ٿm��b��@���x��3@Nb�^��!?�Z���|�@�&��r�ٿm��b��@���x��3@Nb�^��!?�Z���|�@�&��r�ٿm��b��@���x��3@Nb�^��!?�Z���|�@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@_�'G��ٿc���@�]�> 4@e��z�!?[m���@Q�K�ٿigrI���@�Cc�=4@��A܏!?��_h�@Q�K�ٿigrI���@�Cc�=4@��A܏!?��_h�@Q�K�ٿigrI���@�Cc�=4@��A܏!?��_h�@Q�K�ٿigrI���@�Cc�=4@��A܏!?��_h�@E�E�ٿK�WX��@���F 4@���F��!?��/���@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@=��@�ٿ�}$,.��@�p���3@�M`@��!?��OZ�@	�d�2�ٿ2���
��@�����4@sN\{�!?��4���@q?�>�ٿq.�w�@�n\��4@R��v��!?��M{�@�Ӄ;�ٿ�f�z'�@ }`O4@4:([r�!?$��}� �@�Ӄ;�ٿ�f�z'�@ }`O4@4:([r�!?$��}� �@�Ӄ;�ٿ�f�z'�@ }`O4@4:([r�!?$��}� �@�Ӄ;�ٿ�f�z'�@ }`O4@4:([r�!?$��}� �@�Ӄ;�ٿ�f�z'�@ }`O4@4:([r�!?$��}� �@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@����Ǡٿ	��Q��@գ%�+4@�U���!?��$�0��@x��$�ٿi-m�2^�@4�\��3@^�6���!?��JS ��@4�ѝ^�ٿ�5���@��j�3@"\��K�!?s����@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@_��+�ٿOX<~���@ �?��3@=�}��!?mVB(�t�@C���"�ٿ�
L;��@���3@Q��V~�!?��m��@B�[@/�ٿ������@�n&���3@��g죏!?W�Vp��@B�[@/�ٿ������@�n&���3@��g죏!?W�Vp��@B�[@/�ٿ������@�n&���3@��g죏!?W�Vp��@���ݼ�ٿ�Ң�h�@�*7�4@�]Bd�!?X�(���@65�릞ٿ��c]�H�@Hj7��4@�.��y�!?�G����@65�릞ٿ��c]�H�@Hj7��4@�.��y�!?�G����@��l?�ٿ��$]�@q�Մ� 4@ dj�ʏ!?JH:�#�@��l?�ٿ��$]�@q�Մ� 4@ dj�ʏ!?JH:�#�@��l?�ٿ��$]�@q�Մ� 4@ dj�ʏ!?JH:�#�@~�Dv��ٿʞ� \#�@�]^�� 4@8��!?�ۑ���@����ٿx�*��@ӆⓣ4@��%T�!?��]���@����ٿx�*��@ӆⓣ4@��%T�!?��]���@����ٿx�*��@ӆⓣ4@��%T�!?��]���@����ٿx�*��@ӆⓣ4@��%T�!?��]���@����ٿx�*��@ӆⓣ4@��%T�!?��]���@��|��ٿ���O�@�h�4@~��M�!?X����@��|��ٿ���O�@�h�4@~��M�!?X����@��|��ٿ���O�@�h�4@~��M�!?X����@��|��ٿ���O�@�h�4@~��M�!?X����@��|��ٿ���O�@�h�4@~��M�!?X����@�o�:N�ٿ����|��@�����4@��M��!?��?�J��@�o�:N�ٿ����|��@�����4@��M��!?��?�J��@�a.5�ٿʙ�o���@h),]4@�8@��!?xk7���@�a.5�ٿʙ�o���@h),]4@�8@��!?xk7���@�a.5�ٿʙ�o���@h),]4@�8@��!?xk7���@�a.5�ٿʙ�o���@h),]4@�8@��!?xk7���@�a.5�ٿʙ�o���@h),]4@�8@��!?xk7���@i�UC4�ٿ����r�@M�)F�4@���m�!?D��o�@i�UC4�ٿ����r�@M�)F�4@���m�!?D��o�@i�UC4�ٿ����r�@M�)F�4@���m�!?D��o�@i�UC4�ٿ����r�@M�)F�4@���m�!?D��o�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@�6�0�ٿ�{�!C��@�*�/ 4@����!?#T�[qu�@sM�*Ѣٿ[�f���@>�2�a�3@U$!s�!?4qztR�@sM�*Ѣٿ[�f���@>�2�a�3@U$!s�!?4qztR�@sM�*Ѣٿ[�f���@>�2�a�3@U$!s�!?4qztR�@(�%7_�ٿc���e�@�2�[ 4@�y��f�!?n��Di�@(�%7_�ٿc���e�@�2�[ 4@�y��f�!?n��Di�@(�%7_�ٿc���e�@�2�[ 4@�y��f�!?n��Di�@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@踬ћٿ@@5�i�@H{��L 4@H�H���!?�n�>F��@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@K�cU�ٿ �[�)�@k�E� 4@��Aڏ!?$��E�@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@���B�ٿ���Lf��@"K
��4@��7�ݏ!?�..d���@I��]s�ٿ�
ra��@��, �4@tY��̏!?:Z����@I��]s�ٿ�
ra��@��, �4@tY��̏!?:Z����@I��]s�ٿ�
ra��@��, �4@tY��̏!?:Z����@�$=�ٿz�����@�O�` 4@�W�ُ!?1W��@�$=�ٿz�����@�O�` 4@�W�ُ!?1W��@�$=�ٿz�����@�O�` 4@�W�ُ!?1W��@�$=�ٿz�����@�O�` 4@�W�ُ!?1W��@
�x��ٿ����|�@E}�� 4@k�Ɉ�!?���sǃ�@
�x��ٿ����|�@E}�� 4@k�Ɉ�!?���sǃ�@�/�ٿd|I)���@��4@�0�}k�!?߁
���@�/�ٿd|I)���@��4@�0�}k�!?߁
���@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@k���+�ٿ�=�Q���@]��E�4@�z ��!?uQ�7Y��@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@o���ٿ��Q�[�@vdN� 4@���֋�!?�r�O�p�@�Ɵ	СٿAU��MM�@*O(4@��G�F�!?p&#�v�@�kz�ٿ���g�p�@:���s4@��c�ُ!?�.�2��@�kz�ٿ���g�p�@:���s4@��c�ُ!?�.�2��@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@9Bm���ٿ}��}O��@�0��4@6�T��!?S��bC-�@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@���F�ٿo^�d%��@�c[\4@��)h��!?�H��.��@�V��g�ٿrξ����@���x 4@�����!?������@�V��g�ٿrξ����@���x 4@�����!?������@Ǎ퍙ٿX����@{�ueM4@�3 dŏ!?C9�s��@Ǎ퍙ٿX����@{�ueM4@�3 dŏ!?C9�s��@Ǎ퍙ٿX����@{�ueM4@�3 dŏ!?C9�s��@�,f��ٿ$���p��@� �j�4@ܫ\/��!?@���c�@�,f��ٿ$���p��@� �j�4@ܫ\/��!?@���c�@�,f��ٿ$���p��@� �j�4@ܫ\/��!?@���c�@�,f��ٿ$���p��@� �j�4@ܫ\/��!?@���c�@f�ᦘ�ٿZ0r6���@�c��F4@9p����!?3G���\�@f�ᦘ�ٿZ0r6���@�c��F4@9p����!?3G���\�@R�9P�ٿ34����@D�q}g4@��C���!?����@R�9P�ٿ34����@D�q}g4@��C���!?����@R�9P�ٿ34����@D�q}g4@��C���!?����@R�9P�ٿ34����@D�q}g4@��C���!?����@R�9P�ٿ34����@D�q}g4@��C���!?����@R�9P�ٿ34����@D�q}g4@��C���!?����@�_jF��ٿ-U�)�@��lZ��3@�ƅl��!?���k���@�_jF��ٿ-U�)�@��lZ��3@�ƅl��!?���k���@�_jF��ٿ-U�)�@��lZ��3@�ƅl��!?���k���@�_jF��ٿ-U�)�@��lZ��3@�ƅl��!?���k���@�_jF��ٿ-U�)�@��lZ��3@�ƅl��!?���k���@;W��ٿ��T�@�Dj���3@vcꠓ�!? �w����@;W��ٿ��T�@�Dj���3@vcꠓ�!? �w����@�8����ٿ�`�L�@�[-�4@�2c��!?8�|����@�8����ٿ�`�L�@�[-�4@�2c��!?8�|����@G`/?�ٿ}��`�;�@X�K�g 4@�~���!?�$��S�@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@r� ښٿd�Gt���@4`���4@~��ؕ�!?�W^aW��@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@���2�ٿ|�o�6�@��.�O�3@�x%Aӏ!?ȴ�u,�@@V��!�ٿ��Q��@�HW�4@[�ۏ!?��M�vz�@@V��!�ٿ��Q��@�HW�4@[�ۏ!?��M�vz�@U;����ٿ�Μ���@�,��I4@�$튠�!??}H�# �@���Ap�ٿyvVlw��@��Hg� 4@vX"��!?8}d�@���Ap�ٿyvVlw��@��Hg� 4@vX"��!?8}d�@�B���ٿk򇭑��@��`��3@�/@���!?~���@�B���ٿk򇭑��@��`��3@�/@���!?~���@�B���ٿk򇭑��@��`��3@�/@���!?~���@�&a�v�ٿ�DH���@r����3@���4��!?������@����ٿEc9����@�����3@\I���!?�N���@����ٿEc9����@�����3@\I���!?�N���@����ٿEc9����@�����3@\I���!?�N���@�ihK�ٿ"�r���@�&	=�3@y�|~�!?v�2�,A�@�ihK�ٿ"�r���@�&	=�3@y�|~�!?v�2�,A�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@��tlߥٿ,�0�6��@���T)�3@������!?$��p�H�@f8�\�ٿ5���@�i �h�3@Z=�F�!?H[r ��@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@� q��ٿJ�"j�@t!�i^�3@�V:���!?ٚ\����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�E�p�ٿ?r�Cd��@��l�r 4@g�%�ҏ!?�4.����@�w��ٿ{u�����@�嗎)�3@�c�ԏ!?_�ҢO��@�w��ٿ{u�����@�嗎)�3@�c�ԏ!?_�ҢO��@�w��ٿ{u�����@�嗎)�3@�c�ԏ!?_�ҢO��@���ٿ	�x��N�@�X�)��3@1QV&��!?%�1 :�@���ٿ	�x��N�@�X�)��3@1QV&��!?%�1 :�@0JY�_�ٿ�$$�t�@�gЦ4@�<a��!?7AH��@0JY�_�ٿ�$$�t�@�gЦ4@�<a��!?7AH��@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@��\��ٿ�"�Em�@� �� 4@��I4��!?�����@���ܭٿ�?|���@��:{��3@��Sm�!?��熱��@���ܭٿ�?|���@��:{��3@��Sm�!?��熱��@�?�k��ٿU�<���@�zIv� 4@;!s��!?�9���@$I̷6�ٿ��r���@%�k?;4@D��r�!?T�坷�@$I̷6�ٿ��r���@%�k?;4@D��r�!?T�坷�@$I̷6�ٿ��r���@%�k?;4@D��r�!?T�坷�@,V��ٿ�]wc��@�<�}4@$}4��!?�"����@,V��ٿ�]wc��@�<�}4@$}4��!?�"����@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�0��ٿ��(E���@�
{Hs4@���m��!?�8犀!�@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@�E�ٿǼLT!��@ֲȸ4@#5"ɣ�!?>��� ��@���5(�ٿn�����@JLsZ4@$ujbO�!?D���ze�@���5(�ٿn�����@JLsZ4@$ujbO�!?D���ze�@v���ߦٿ�-�X�@r�7BF4@H�8V��!?��nq��@v���ߦٿ�-�X�@r�7BF4@H�8V��!?��nq��@ܻ@�4�ٿ�U�(�@k �4m�3@��Om�!?�<�a�u�@ܻ@�4�ٿ�U�(�@k �4m�3@��Om�!?�<�a�u�@ܻ@�4�ٿ�U�(�@k �4m�3@��Om�!?�<�a�u�@s�g�ٿN:�3��@�I����3@J���!?�Dq��@s�g�ٿN:�3��@�I����3@J���!?�Dq��@s�g�ٿN:�3��@�I����3@J���!?�Dq��@�阼8�ٿ�֙ʥ��@������3@���c��!?��r��@�阼8�ٿ�֙ʥ��@������3@���c��!?��r��@ǣ�]��ٿM�M���@�"����3@^ɐ���!?iL�ܣ�@o���ٿ������@.ȇZ 4@�����!?ϵ���@o���ٿ������@.ȇZ 4@�����!?ϵ���@�|���ٿ[�~��@�E��[ 4@��oz�!?���h��@��ԑ�ٿ�u^�(w�@HE���3@cjn?�!?�5�����@��ԑ�ٿ�u^�(w�@HE���3@cjn?�!?�5�����@�����ٿJtpv�@ KF2� 4@L��8�!?��J&�@�����ٿJtpv�@ KF2� 4@L��8�!?��J&�@�i���ٿ�CD��@���4@���I�!?����@�i���ٿ�CD��@���4@���I�!?����@+v���ٿ`D&�V��@7LR 4@�!?�!r��@+v���ٿ`D&�V��@7LR 4@�!?�!r��@+v���ٿ`D&�V��@7LR 4@�!?�!r��@+v���ٿ`D&�V��@7LR 4@�!?�!r��@+v���ٿ`D&�V��@7LR 4@�!?�!r��@���'M�ٿJ����@=�ww 4@u���p�!?L��F���@���'M�ٿJ����@=�ww 4@u���p�!?L��F���@���'M�ٿJ����@=�ww 4@u���p�!?L��F���@���'M�ٿJ����@=�ww 4@u���p�!?L��F���@���'M�ٿJ����@=�ww 4@u���p�!?L��F���@���z�ٿ���#E��@��=)4@�}���!?���+Nf�@���z�ٿ���#E��@��=)4@�}���!?���+Nf�@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@Ԝ�.w�ٿ�9�ժ��@�<Xi��3@>W�』!?�~v���@������ٿ�9|Y���@�?,  4@&�&3��!?7�����@������ٿ�9|Y���@�?,  4@&�&3��!?7�����@������ٿ�9|Y���@�?,  4@&�&3��!?7�����@������ٿ�9|Y���@�?,  4@&�&3��!?7�����@&��o�ٿ:��3e��@��'�� 4@%�g��!?�":.*�@&��o�ٿ:��3e��@��'�� 4@%�g��!?�":.*�@&��o�ٿ:��3e��@��'�� 4@%�g��!?�":.*�@�0�	{�ٿ7������@*d�Pv4@U�)��!?�>4��#�@�0�	{�ٿ7������@*d�Pv4@U�)��!?�>4��#�@�0�	{�ٿ7������@*d�Pv4@U�)��!?�>4��#�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@��P�ݧٿ�>�zc��@^g{a� 4@N���p�!?��\53G�@j�����ٿp��ڽ|�@�S�K4@�Z�)͏!?�D�F%��@j�����ٿp��ڽ|�@�S�K4@�Z�)͏!?�D�F%��@j�����ٿp��ڽ|�@�S�K4@�Z�)͏!?�D�F%��@ǆ�#��ٿ&?���K�@ktqh�3@�H�)ҏ!?��@�{�@y�r�ٿ܋K9p��@��!m 4@�r߾�!?�u����@y�r�ٿ܋K9p��@��!m 4@�r߾�!?�u����@y�r�ٿ܋K9p��@��!m 4@�r߾�!?�u����@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@�o`�ٿ�P/��@�mj��3@%�H��!?��G�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@��t(_�ٿ"g��s�@~����4@���!?G��$�@�K�/&�ٿ3GV�V�@�$f 4@�����!?b�L�Mr�@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�!,3��ٿE�;�Y��@-B��3@����!?�� ��@�\��^�ٿ�=�i�u�@/���u 4@��?q��!?�#ך��@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@�{�ٿ$��`k��@r��rj4@��CՇ�!?�Ń����@��`�Ȧٿ��hhP��@�� S! 4@3��s��!?ݰ�y9��@��`�Ȧٿ��hhP��@�� S! 4@3��s��!?ݰ�y9��@��`�Ȧٿ��hhP��@�� S! 4@3��s��!?ݰ�y9��@��`�Ȧٿ��hhP��@�� S! 4@3��s��!?ݰ�y9��@�p]�\�ٿfnV�K^�@�	'�3@��|h��!?�5��P��@�p]�\�ٿfnV�K^�@�	'�3@��|h��!?�5��P��@�p]�\�ٿfnV�K^�@�	'�3@��|h��!?�5��P��@�p]�\�ٿfnV�K^�@�	'�3@��|h��!?�5��P��@�p]�\�ٿfnV�K^�@�	'�3@��|h��!?�5��P��@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@9j�!4�ٿ�}�$M��@��8Ze�3@:��ٮ�!?��+c���@#�� �ٿs�?a��@�[�4�3@2[�k��!?u��i�!�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@C�(���ٿlb�X�@W��\3�3@�$���!?f�45�@��Zo�ٿ
MM7|��@�C�O��3@�Ãݧ�!?|`�C�c�@/M�ٿs���'��@H�>�3@�`��!?�!�j��@/M�ٿs���'��@H�>�3@�`��!?�!�j��@/M�ٿs���'��@H�>�3@�`��!?�!�j��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@1��N�ٿg��c��@��9��3@��Y�!?�ePa>��@ߣ~�4�ٿa� A߯�@����3@;�'�T�!?�=o��@ߣ~�4�ٿa� A߯�@����3@;�'�T�!?�=o��@ߣ~�4�ٿa� A߯�@����3@;�'�T�!?�=o��@ߣ~�4�ٿa� A߯�@����3@;�'�T�!?�=o��@��2�ٿ+ӊ���@xEa���3@@i ϥ�!?z��[�D�@���ٿ&*�#�?�@�>�v��3@�22j��!?и��9��@G6\�ٿ��Z��t�@��k��3@���8�!?�#$E���@G6\�ٿ��Z��t�@��k��3@���8�!?�#$E���@G6\�ٿ��Z��t�@��k��3@���8�!?�#$E���@Q��Ġٿ�=�β��@2,U� 4@�-@�U�!?�u�"���@T5O�ٿ�d�����@��/^k�3@9��ժ�!?�����@T5O�ٿ�d�����@��/^k�3@9��ժ�!?�����@T5O�ٿ�d�����@��/^k�3@9��ժ�!?�����@T5O�ٿ�d�����@��/^k�3@9��ժ�!?�����@T5O�ٿ�d�����@��/^k�3@9��ժ�!?�����@����՜ٿO������@��b  4@;����!?�TT���@����՜ٿO������@��b  4@;����!?�TT���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@?��_�ٿ)Vk�s��@}�4@����!?���l���@�{�hT�ٿat���@��^
4@�q��ԏ!?a�57��@�{�hT�ٿat���@��^
4@�q��ԏ!?a�57��@�{�hT�ٿat���@��^
4@�q��ԏ!?a�57��@?7�ױٿl�{�5��@!~	F�4@RcM�ޏ!?�S=�@i��L�ٿ�K橼��@�m1O4@�p(�o�!?IR )���@i��L�ٿ�K橼��@�m1O4@�p(�o�!?IR )���@��y.�ٿ��A�2�@~l��R 4@o#+��!?��M��@��y.�ٿ��A�2�@~l��R 4@o#+��!?��M��@��y.�ٿ��A�2�@~l��R 4@o#+��!?��M��@��y.�ٿ��A�2�@~l��R 4@o#+��!?��M��@��y.�ٿ��A�2�@~l��R 4@o#+��!?��M��@�h��[�ٿ�j{��@�[�T�4@,f�p�!?d�2(jg�@�Ɋw�ٿ|�	�/�@>'Ud4@�)�!?2^ӹL��@�,�ȟٿ,\�L��@Ơ�4@���Z-�!?߰�J�@*6��ٿ�5z�@;ɐ�34@�ۯe�!?����)�@*6��ٿ�5z�@;ɐ�34@�ۯe�!?����)�@*6��ٿ�5z�@;ɐ�34@�ۯe�!?����)�@*6��ٿ�5z�@;ɐ�34@�ۯe�!?����)�@�m�\ɪٿ{��T��@��c� 4@8V��!?�f?�A�@�ʙVN�ٿ�e/�r.�@ SOs�4@�6�[�!?p��Qy�@�ʙVN�ٿ�e/�r.�@ SOs�4@�6�[�!?p��Qy�@�ʙVN�ٿ�e/�r.�@ SOs�4@�6�[�!?p��Qy�@�ʙVN�ٿ�e/�r.�@ SOs�4@�6�[�!?p��Qy�@�ʙVN�ٿ�e/�r.�@ SOs�4@�6�[�!?p��Qy�@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�Ӝ�ٿH߹�)T�@���I��3@�uG�i�!?l��z��@�1+מٿ��'����@���3@����Z�!?��ql��@�1+מٿ��'����@���3@����Z�!?��ql��@�1+מٿ��'����@���3@����Z�!?��ql��@�1+מٿ��'����@���3@����Z�!?��ql��@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@_ǠƘ�ٿ!(�-�e�@��^�w4@J32ں�!?�! �.�@�lB>�ٿ��>��J�@����5 4@o�䝏!?��[��@�lB>�ٿ��>��J�@����5 4@o�䝏!?��[��@�lB>�ٿ��>��J�@����5 4@o�䝏!?��[��@�lB>�ٿ��>��J�@����5 4@o�䝏!?��[��@���/�ٿ��M�2J�@�va4@r����!?eg��H�@���/�ٿ��M�2J�@�va4@r����!?eg��H�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@��A�ٿc3��\��@���ѯ 4@< J��!?MBKFd~�@�	:
��ٿ������@�4��4@4��%͏!?��ƨ�%�@�	:
��ٿ������@�4��4@4��%͏!?��ƨ�%�@�	:
��ٿ������@�4��4@4��%͏!?��ƨ�%�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@E@B��ٿ�����y�@�G�BQ 4@x�=�Տ!?���R?�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@KAtZ�ٿNK��A��@��f�� 4@��O�!?��Q�@
ڂQ�ٿe-��.n�@}[L�4@p܎��!?����k��@
ڂQ�ٿe-��.n�@}[L�4@p܎��!?����k��@Y���^�ٿ���˨�@wԦ! 4@F����!?����@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@w�h�Ūٿ����u�@0e/E�4@�s�]��!?d�{io�@X61�ٿ4��1�:�@��r�� 4@t�J&N�!?b�y��@X61�ٿ4��1�:�@��r�� 4@t�J&N�!?b�y��@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@ωGҨٿ�d{8m�@} 4@��lF�!?���/�@���|�ٿ�Em����@���K7 4@!��Z��!?���
�x�@���|�ٿ�Em����@���K7 4@!��Z��!?���
�x�@���|�ٿ�Em����@���K7 4@!��Z��!?���
�x�@���|�ٿ�Em����@���K7 4@!��Z��!?���
�x�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@��)��ٿ�t�l��@ߔN|�4@hΚ�o�!?t2jj�D�@aM��S�ٿxh�us'�@*�,4@ڟ4O�!?�����@aM��S�ٿxh�us'�@*�,4@ڟ4O�!?�����@�9�y�ٿ��-i;�@���a4@E��~�!?h5-��k�@�9�y�ٿ��-i;�@���a4@E��~�!?h5-��k�@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�1�3�ٿu�1W��@=�a���3@�P8�v�!?�ڡC���@�7Lg��ٿF�Rڱc�@(��3�3@��)/��!?��ny��@�7Lg��ٿF�Rڱc�@(��3�3@��)/��!?��ny��@�7Lg��ٿF�Rڱc�@(��3�3@��)/��!?��ny��@�7Lg��ٿF�Rڱc�@(��3�3@��)/��!?��ny��@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@L�hM�ٿ#�\*��@t	�Zz 4@trQOi�!?8��'x�@�Em��ٿ�a�޴��@!T��4@�Or�!?D��#���@MA���ٿ2���<��@�s�}+4@S��X�!?\+Z��A�@MA���ٿ2���<��@�s�}+4@S��X�!?\+Z��A�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@.mb��ٿ)U	�ġ�@��.+4@��\�!?>ݥ�[�@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@�d�!�ٿ�.����@�uZ:� 4@p@ S~�!?��H5���@���u�ٿ��r��@K��dy 4@:��ď!?��\��Z�@�>����ٿ�'���@�{���3@_{�+��!?l�V���@OopPs�ٿ/��":�@B\O�4@������!?W�<X,�@7L���ٿ���X�@�� 4@6ZhG�!?bMg*4<�@7L���ٿ���X�@�� 4@6ZhG�!?bMg*4<�@7L���ٿ���X�@�� 4@6ZhG�!?bMg*4<�@7L���ٿ���X�@�� 4@6ZhG�!?bMg*4<�@7L���ٿ���X�@�� 4@6ZhG�!?bMg*4<�@�$:.��ٿ�� ���@���� 4@��}5��!?t�����@�$:.��ٿ�� ���@���� 4@��}5��!?t�����@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@��C �ٿ\�b5k�@IG7с�3@&8|�!?$3�L<�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@�
�ٿ�<��Z�@�؎���3@{�d���!?�+�@!j���ٿ`�D)R�@�!kcp�3@~���!?�]�=���@!j���ٿ`�D)R�@�!kcp�3@~���!?�]�=���@!j���ٿ`�D)R�@�!kcp�3@~���!?�]�=���@!j���ٿ`�D)R�@�!kcp�3@~���!?�]�=���@!j���ٿ`�D)R�@�!kcp�3@~���!?�]�=���@eH�26�ٿ�n9$��@�I�6C�3@.�L�~�!?�j�%��@eH�26�ٿ�n9$��@�I�6C�3@.�L�~�!?�j�%��@eH�26�ٿ�n9$��@�I�6C�3@.�L�~�!?�j�%��@�?��ٿ�ߟ@���@l�w34@c�N�!?S�n���@���n�ٿS��ND��@��~5(4@ A
�V�!?,9Z����@���n�ٿS��ND��@��~5(4@ A
�V�!?,9Z����@���n�ٿS��ND��@��~5(4@ A
�V�!?,9Z����@���n�ٿS��ND��@��~5(4@ A
�V�!?,9Z����@���n�ٿS��ND��@��~5(4@ A
�V�!?,9Z����@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@&*�ݳ�ٿ��K	c�@bC>v�4@\�x!?D�}V�*�@A�ۗٿ�xw:h�@r����4@�uo��!?2~���@~���ٿ��M�@��E�4@ۿ��؏!?��m�'��@�.���ٿm>���@>�}��4@{��!?=8�VZ�@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@A�5��ٿY��ZH�@�k���4@NDW��!?�
szX��@��" �ٿ��\B�@v���3@¯��!?�Fg��@��" �ٿ��\B�@v���3@¯��!?�Fg��@��" �ٿ��\B�@v���3@¯��!?�Fg��@��" �ٿ��\B�@v���3@¯��!?�Fg��@��" �ٿ��\B�@v���3@¯��!?�Fg��@��" �ٿ��\B�@v���3@¯��!?�Fg��@<<��ٿ�"�h�'�@��y: 4@IMI��!?m�4b�n�@<<��ٿ�"�h�'�@��y: 4@IMI��!?m�4b�n�@תMA�ٿ��|�@J`�c�3@l�(ʏ!?mҠ1��@תMA�ٿ��|�@J`�c�3@l�(ʏ!?mҠ1��@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@�|@+%�ٿL��d�6�@T�)K� 4@i����!?���I�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@`6x@�ٿ���4���@R�Hx4@�P��!?�Wh�x�@�Ln0�ٿ]ÂN0��@�S�F<4@wѢk��!?bXz��D�@�Ln0�ٿ]ÂN0��@�S�F<4@wѢk��!?bXz��D�@6�z�r�ٿ��	����@>p�K� 4@�Qy봏!?.�n[S�@6�z�r�ٿ��	����@>p�K� 4@�Qy봏!?.�n[S�@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@�͵:�ٿb��n�@�ǯW 4@��jr��!?XM���@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@a!�˘ٿ�yU�|�@҄�� 4@�YȺ��!?n�� �@�tz~ٕٿ�% )v��@�ƕ 4@)M���!?��yY���@�tz~ٕٿ�% )v��@�ƕ 4@)M���!?��yY���@�tz~ٕٿ�% )v��@�ƕ 4@)M���!?��yY���@>ˣ�ٿ���S�@$ h�4@a���!?Kۿ�}�@>ˣ�ٿ���S�@$ h�4@a���!?Kۿ�}�@>ˣ�ٿ���S�@$ h�4@a���!?Kۿ�}�@>ˣ�ٿ���S�@$ h�4@a���!?Kۿ�}�@�ԋ�Șٿ��I��@@��&4@���ȏ!?~�!9R�@�ԋ�Șٿ��I��@@��&4@���ȏ!?~�!9R�@�ԋ�Șٿ��I��@@��&4@���ȏ!?~�!9R�@�ԋ�Șٿ��I��@@��&4@���ȏ!?~�!9R�@T=Pݖٿ�Y�J�#�@�(ڣ0�3@���!��!?Yq�����@��ZW��ٿaE�9"��@�n۵Y�3@4=�nُ!?�����@��ZW��ٿaE�9"��@�n۵Y�3@4=�nُ!?�����@��ZW��ٿaE�9"��@�n۵Y�3@4=�nُ!?�����@��ZW��ٿaE�9"��@�n۵Y�3@4=�nُ!?�����@'�"�ˑٿn!��U��@�����3@��6��!?�����@��}��ٿvŘ��@�C>�{�3@�_���!?��@C�u�@��}��ٿvŘ��@�C>�{�3@�_���!?��@C�u�@��}��ٿvŘ��@�C>�{�3@�_���!?��@C�u�@���B�ٿ�w����@�yv��3@�5�!?�[YgX��@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@�v���ٿ"�i����@�j̻�3@-z��}�!?���.(�@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@b�Oߜٿ���N>��@^����3@*̌y�!?�	;���@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@H�:;�ٿ���7��@9ܡ�W 4@c2&�s�!?��|����@o{xb�ٿ�����@�h"u 4@\�F�k�!?`I5�
��@o{xb�ٿ�����@�h"u 4@\�F�k�!?`I5�
��@o{xb�ٿ�����@�h"u 4@\�F�k�!?`I5�
��@�Ʉ��ٿ��w<��@�;���3@u9�C�!?���&'�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@s}� $�ٿ�6����@$�8�� 4@=����!?G��<�@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@P�ofY�ٿ��l����@'�	E1 4@��U���!?��X���@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�Z���ٿb0XL��@�D �4@�*$v͏!?.mH7u��@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�.剢ٿ9�2�`�@���S4@����ŏ!?���
�@�T��ٿ��*ez�@tDK| 4@�=�	��!?*bs�-��@�T��ٿ��*ez�@tDK| 4@�=�	��!?*bs�-��@�T��ٿ��*ez�@tDK| 4@�=�	��!?*bs�-��@�>ڡ��ٿ�X4b�@l7D& 4@��fm�!?�,�!�@�>ڡ��ٿ�X4b�@l7D& 4@��fm�!?�,�!�@�ȴJ��ٿ�A�#e�@_̌h�3@�3v�!?�o�˟!�@�ȴJ��ٿ�A�#e�@_̌h�3@�3v�!?�o�˟!�@�ȴJ��ٿ�A�#e�@_̌h�3@�3v�!?�o�˟!�@�M����ٿ)k����@f�6��3@��pzW�!?8��uTy�@�M����ٿ)k����@f�6��3@��pzW�!?8��uTy�@~=wj�ٿ@��4��@����) 4@�����!?ݿa��*�@87s̲�ٿ^��|���@��"T��3@_�bnX�!?q��vI�@(���6�ٿ�]�5��@�ߖ�4@�%��!?��˞�@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@	�q�ٿď�1���@4�}/|4@����!?V0�����@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@\x|�	�ٿ>*󣻳�@��^]S4@�����!?�V��O�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�yA�s�ٿ��� i��@��t�	4@�umt��!?CV��K�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@�`o���ٿ*�|���@6�a� 4@#@,���!?�E��}�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@k��K��ٿ�O2�+��@:��?4@�C��!?�Ѥ�s?�@ Ek_.�ٿ������@�Ye�� 4@32��q�!?��?�<�@ Ek_.�ٿ������@�Ye�� 4@32��q�!?��?�<�@ Ek_.�ٿ������@�Ye�� 4@32��q�!?��?�<�@ Ek_.�ٿ������@�Ye�� 4@32��q�!?��?�<�@ Ek_.�ٿ������@�Ye�� 4@32��q�!?��?�<�@3	)Śٿ�!B���@T��e4@jr��!?��H;���@3	)Śٿ�!B���@T��e4@jr��!?��H;���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@�9�y��ٿ|�B�b��@d����3@�Y~�!?L�9���@��*a�ٿ._c��@�ǧ�3@��2���!?W��[��@��.���ٿ�SC���@;|<N� 4@��ď!?�<�̽V�@�K����ٿ�跘��@�����3@&��ބ�!?�Z?��.�@�K����ٿ�跘��@�����3@&��ބ�!?�Z?��.�@�d��ٿk�"�N��@�K�Kt 4@G0Z ��!?��Enz��@�d��ٿk�"�N��@�K�Kt 4@G0Z ��!?��Enz��@�d��ٿk�"�N��@�K�Kt 4@G0Z ��!?��Enz��@�Ecw؟ٿ�u���@y7_��3@�Ji���!?���N��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@3�66�ٿ���YP��@�(��9 4@�l�ׄ�!?x^��@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@�x���ٿ��IA��@iD��Q�3@�u����!?�z��I:�@q쥳y�ٿ��6���@����9 4@wb4֒�!?WaDI<�@q쥳y�ٿ��6���@����9 4@wb4֒�!?WaDI<�@���o��ٿ~_���@V⫭ 4@�K߶�!?/NM�A�@���o��ٿ~_���@V⫭ 4@�K߶�!?/NM�A�@���o��ٿ~_���@V⫭ 4@�K߶�!?/NM�A�@���o��ٿ~_���@V⫭ 4@�K߶�!?/NM�A�@�@d�ٿ����@���� 4@}!�[��!?T���@�@d�ٿ����@���� 4@}!�[��!?T���@�U�e�ٿ��d�ĕ�@&떼S 4@u����!?��抽�@�U�e�ٿ��d�ĕ�@&떼S 4@u����!?��抽�@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@��1�ٿ�a-�e��@��F� 4@�혁�!?�Xt����@s�x3��ٿ|�k�r�@�K� 4@e׫�I�!?��z���@s�x3��ٿ|�k�r�@�K� 4@e׫�I�!?��z���@s�x3��ٿ|�k�r�@�K� 4@e׫�I�!?��z���@s�x3��ٿ|�k�r�@�K� 4@e׫�I�!?��z���@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@��i�
�ٿX�5�g�@,~˴�3@�[e��!?��-؎�@���ɰٿ����C�@��㠛�3@@S[Xh�!?�R�����@�]�֩ٿ�d� ��@�Y@0 4@�QG�!?�wSL&�@�]�֩ٿ�d� ��@�Y@0 4@�QG�!?�wSL&�@�]�֩ٿ�d� ��@�Y@0 4@�QG�!?�wSL&�@�]�֩ٿ�d� ��@�Y@0 4@�QG�!?�wSL&�@��Z��ٿm���`��@|Rۆ+ 4@��VM�!?�%��-R�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@���D�ٿ8[x���@���3m4@qF؊.�!?�w��"�@��$�ٿ�Y�U�c�@u�ߍO4@z���K�!?L'�nr�@Q8���ٿ��lU���@�1xZ 4@��u]�!?8��K��@ze=�=�ٿ�5��2��@����4@�`�W�!?�������@ze=�=�ٿ�5��2��@����4@�`�W�!?�������@ze=�=�ٿ�5��2��@����4@�`�W�!?�������@	�����ٿ��ˎϜ�@��Q4@8���!?9g[Z*��@	�����ٿ��ˎϜ�@��Q4@8���!?9g[Z*��@	�����ٿ��ˎϜ�@��Q4@8���!?9g[Z*��@	�����ٿ��ˎϜ�@��Q4@8���!?9g[Z*��@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@��c��ٿ{=dML�@߫�4@�����!?S�H{AD�@�$�(�ٿ�Zd���@��!�4@p�]岏!?����y��@�$�(�ٿ�Zd���@��!�4@p�]岏!?����y��@I�h�ٿ�H�n�@��*`�4@�g�Ǐ!?�2HD���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@3�wU�ٿY�R�5��@{��U4@?!�+^�!?��;���@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@q���ҧٿ:�pZ��@a�+i4@�)�莏!?����d��@�ٺx�ٿ�|j�S�@, 	7v 4@ ՞���!?�]�-��@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@�;���ٿ>t>����@8y��4@�*Uh��!?��ڭ6�@��c�4�ٿ�HB��@j���4@��e��!?���\��@��c�4�ٿ�HB��@j���4@��e��!?���\��@��c�4�ٿ�HB��@j���4@��e��!?���\��@�[��ٿGVB�|�@{�'bY 4@����!?8n��~�@�[��ٿGVB�|�@{�'bY 4@����!?8n��~�@�[��ٿGVB�|�@{�'bY 4@����!?8n��~�@��O�ٿ�`�j�T�@h�= 4@�y��Ϗ!?�M�T_��@ˏ��ٿ�R=���@$}N�]�3@���}�!?��2s��@ˏ��ٿ�R=���@$}N�]�3@���}�!?��2s��@Y��ٿI���z�@�瀅�3@/�˲ڏ!?��-}v|�@Y��ٿI���z�@�瀅�3@/�˲ڏ!?��-}v|�@Y��ٿI���z�@�瀅�3@/�˲ڏ!?��-}v|�@Y��ٿI���z�@�瀅�3@/�˲ڏ!?��-}v|�@Y��ٿI���z�@�瀅�3@/�˲ڏ!?��-}v|�@��/�ٿ&x|��@��V ��3@W�L��!?p���~�@��/�ٿ&x|��@��V ��3@W�L��!?p���~�@�+/s��ٿ|�:�i�@W�i	� 4@�eC|��!?y�Մ`��@�f��ٿ]�։E�@�(�z��3@ ��R��!?g�U�[��@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@(/��ٿF��d��@'@T�3@F�z3��!?H[X>�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��a7i�ٿ(����7�@"t�3j4@4�c7P�!?�S<Zh�@��Wb��ٿJu�j�@�N�x)4@̀.j�!?Ԡ^���@��Wb��ٿJu�j�@�N�x)4@̀.j�!?Ԡ^���@sݪI��ٿ���Ȼ�@�z��*4@)��\�!?��<���@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@?эCΦٿ�R�km:�@hC.4@��{�!?{��(9�@�c-���ٿ'۠�A�@)�%�8 4@� H3r�!?�X���@g.�ٿ����k�@�����3@��x]�!?��+<�@g.�ٿ����k�@�����3@��x]�!?��+<�@g.�ٿ����k�@�����3@��x]�!?��+<�@g.�ٿ����k�@�����3@��x]�!?��+<�@�AVl��ٿ8p���@�o��3@����v�!?kN%ܖ�@�AVl��ٿ8p���@�o��3@����v�!?kN%ܖ�@�AVl��ٿ8p���@�o��3@����v�!?kN%ܖ�@�AVl��ٿ8p���@�o��3@����v�!?kN%ܖ�@�AVl��ٿ8p���@�o��3@����v�!?kN%ܖ�@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@T0�Q.�ٿ����,F�@s�t	� 4@�pzF��!?Q6���@�_;�£ٿX9��.��@E��f\ 4@>l�9�!?D.���N�@�_;�£ٿX9��.��@E��f\ 4@>l�9�!?D.���N�@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@�0kH�ٿX�u}��@�<��4@2Ђܷ�!?����@Z䅍��ٿ#Yǋ�p�@N��m 4@aIۘ�!?�6����@Z䅍��ٿ#Yǋ�p�@N��m 4@aIۘ�!?�6����@��_�H�ٿK�6h��@��'t�3@�|;ny�!?�LW|��@V˭��ٿ)�����@t #ol4@����c�!?�dt��@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@^�J�ٿ��M�@���g� 4@���WΏ!?ڬ�b�_�@�𿬎�ٿǆ���O�@S�@ 4@�7vؒ�!?�%����@�𿬎�ٿǆ���O�@S�@ 4@�7vؒ�!?�%����@�𿬎�ٿǆ���O�@S�@ 4@�7vؒ�!?�%����@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@$�HT�ٿ�(�{���@A�B� 4@����P�!?Դq�;��@nj�\�ٿO%vy��@��u�4@�ҏ!?&}�p@�@nj�\�ٿO%vy��@��u�4@�ҏ!?&}�p@�@nj�\�ٿO%vy��@��u�4@�ҏ!?&}�p@�@1�L�ٿ�蒖�@*����4@=ѭ��!?-��c��@����ٿ��� m��@YD��w4@l����!?��dwJ��@{�̗ٿ���y�@��<�;4@?L��!?�#p�{{�@L����ٿ�Pv�]�@`�>z�4@;�t��!?l �9�'�@L����ٿ�Pv�]�@`�>z�4@;�t��!?l �9�'�@�-Oۜٿb�)U�@�U1΁4@j�U!�!?ЉT�$�@�-Oۜٿb�)U�@�U1΁4@j�U!�!?ЉT�$�@�-Oۜٿb�)U�@�U1΁4@j�U!�!?ЉT�$�@t1���ٿVZ<F���@Ĵt��4@�*'��!?�)腞��@t1���ٿVZ<F���@Ĵt��4@�*'��!?�)腞��@t1���ٿVZ<F���@Ĵt��4@�*'��!?�)腞��@t1���ٿVZ<F���@Ĵt��4@�*'��!?�)腞��@t1���ٿVZ<F���@Ĵt��4@�*'��!?�)腞��@�}�' �ٿ�������@ꁘXA4@�@����!?V����@-���/�ٿ�l��h�@E��� 4@[�����!?kJ$����@-���/�ٿ�l��h�@E��� 4@[�����!?kJ$����@-���/�ٿ�l��h�@E��� 4@[�����!?kJ$����@Tkٖ)�ٿ�Z~׆��@	��, 4@� f��!?23���@��5j��ٿ�nC&��@�ja��3@�_�!?�����@��5j��ٿ�nC&��@�ja��3@�_�!?�����@��5j��ٿ�nC&��@�ja��3@�_�!?�����@}����ٿ��w�I�@u��� 4@)�0u�!?�*�AP��@}����ٿ��w�I�@u��� 4@)�0u�!?�*�AP��@}����ٿ��w�I�@u��� 4@)�0u�!?�*�AP��@dw�ʧٿ��{0�d�@\1qa 4@C��1�!? $�i���@���yx�ٿN��aD�@΁��3@��e:4�!?���2��@hexp�ٿ������@�5�}4@�C/i�!?'H��8H�@׬9 1�ٿ�9�<ł�@	�q�*4@��?�X�!?c��]o��@׬9 1�ٿ�9�<ł�@	�q�*4@��?�X�!?c��]o��@qjUp��ٿ�b�s'�@�:o94@4�o=�!?�	����@qjUp��ٿ�b�s'�@�:o94@4�o=�!?�	����@qjUp��ٿ�b�s'�@�:o94@4�o=�!?�	����@qjUp��ٿ�b�s'�@�:o94@4�o=�!?�	����@qjUp��ٿ�b�s'�@�:o94@4�o=�!?�	����@�Ȧ�ٿ��	M�W�@	�2A4@��Ӌh�!?�,I)\��@�Ȧ�ٿ��	M�W�@	�2A4@��Ӌh�!?�,I)\��@2%�n��ٿ�=�]O��@��K�4@�x�$ҏ!?�5 {���@2%�n��ٿ�=�]O��@��K�4@�x�$ҏ!?�5 {���@�x�<��ٿ2\:v(�@�n�4@��tŏ!?�}���w�@�x�<��ٿ2\:v(�@�n�4@��tŏ!?�}���w�@�x�<��ٿ2\:v(�@�n�4@��tŏ!?�}���w�@�x�<��ٿ2\:v(�@�n�4@��tŏ!?�}���w�@�x�<��ٿ2\:v(�@�n�4@��tŏ!?�}���w�@�ǋ(�ٿ=s�K�@��:4@ /&��!?�*f�iU�@�7N�ٿQ8T�g��@2_�5�4@MJ�j��!?�9s�Z �@�G쒯ٿ�����@ˠ��X 4@'~w�l�!?�������@�G쒯ٿ�����@ˠ��X 4@'~w�l�!?�������@�G쒯ٿ�����@ˠ��X 4@'~w�l�!?�������@f3��ٿ���,��@.��- 4@y�(��!?�ǎ��y�@f3��ٿ���,��@.��- 4@y�(��!?�ǎ��y�@���w�ٿ���jhu�@d�����3@���dC�!?� �q�@���w�ٿ���jhu�@d�����3@���dC�!?� �q�@���w�ٿ���jhu�@d�����3@���dC�!?� �q�@���w�ٿ���jhu�@d�����3@���dC�!?� �q�@X{����ٿ} ��w�@�$f�b4@���LJ�!?s�a�\��@X{����ٿ} ��w�@�$f�b4@���LJ�!?s�a�\��@X{����ٿ} ��w�@�$f�b4@���LJ�!?s�a�\��@X{����ٿ} ��w�@�$f�b4@���LJ�!?s�a�\��@X{����ٿ} ��w�@�$f�b4@���LJ�!?s�a�\��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@���FA�ٿ�em;L�@���3@ed�U�!? �ԏ)��@<4�7�ٿ��[w���@|����3@�¹"��!?�#�;���@<4�7�ٿ��[w���@|����3@�¹"��!?�#�;���@<4�7�ٿ��[w���@|����3@�¹"��!?�#�;���@<4�7�ٿ��[w���@|����3@�¹"��!?�#�;���@<4�7�ٿ��[w���@|����3@�¹"��!?�#�;���@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@b���ϢٿÞ����@�T+���3@r�u~}�!?	�H��@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@��R�2�ٿ�V0����@�7*�z�3@j/��!?P�d�Y�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@� �ٿ��~�q�@M�A�� 4@�m7��!?�}g�t�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@��®i�ٿ�5�5D�@T8^�	4@)��ȏ!?�녿�	�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@���0�ٿ�0L���@z��j� 4@h����!?���@P�@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@p�X ��ٿ�����@��4U��3@X�v��!?��:B���@9� t��ٿ��Y%��@��)A4@��w9d�!?yb�6-��@9� t��ٿ��Y%��@��)A4@��w9d�!?yb�6-��@9� t��ٿ��Y%��@��)A4@��w9d�!?yb�6-��@9� t��ٿ��Y%��@��)A4@��w9d�!?yb�6-��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@��i���ٿa٘I
�@�)Pj4@S�u��!?���3o��@gG�N��ٿz��U�@���9V4@�VD	��!?!���^R�@gG�N��ٿz��U�@���9V4@�VD	��!?!���^R�@gG�N��ٿz��U�@���9V4@�VD	��!?!���^R�@gG�N��ٿz��U�@���9V4@�VD	��!?!���^R�@gG�N��ٿz��U�@���9V4@�VD	��!?!���^R�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@�U]� �ٿ�r�4U�@Kr�˔�3@Y���!?�B�X�3�@db�}�ٿ�����@v8Qi 4@U���ޏ!?9�H
���@db�}�ٿ�����@v8Qi 4@U���ޏ!?9�H
���@db�}�ٿ�����@v8Qi 4@U���ޏ!?9�H
���@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@N���	�ٿ4��o��@V(��4@������!?a�/QƯ�@���dF�ٿ(��u��@�Ͳ��3@l����!?N.�N��@�؃2p�ٿ�P"��@����i 4@/k+g��!?��)O�y�@xq�ԟٿL��@�S�C� 4@U�rю�!?�SV��@��'��ٿ���>($�@xjD�N4@��R���!?��B�θ�@��'��ٿ���>($�@xjD�N4@��R���!?��B�θ�@��'��ٿ���>($�@xjD�N4@��R���!?��B�θ�@��'��ٿ���>($�@xjD�N4@��R���!?��B�θ�@%�P��ٿ&kS0O��@�����3@� !﯏!?@%�m��@%�P��ٿ&kS0O��@�����3@� !﯏!?@%�m��@%�P��ٿ&kS0O��@�����3@� !﯏!?@%�m��@%�P��ٿ&kS0O��@�����3@� !﯏!?@%�m��@�H����ٿf�{���@�hT��4@鶮j�!?����&��@�H����ٿf�{���@�hT��4@鶮j�!?����&��@�H����ٿf�{���@�hT��4@鶮j�!?����&��@��GO�ٿSX��@}��u�4@�ϓSO�!?"�]X���@��GO�ٿSX��@}��u�4@�ϓSO�!?"�]X���@��c��ٿ��h��@�rM�4@Uʻp�!?�i���@>�*�ٿ�YV�2�@�I�<�4@�[Џ!?�:�n�	�@>�*�ٿ�YV�2�@�I�<�4@�[Џ!?�:�n�	�@>�*�ٿ�YV�2�@�I�<�4@�[Џ!?�:�n�	�@>�*�ٿ�YV�2�@�I�<�4@�[Џ!?�:�n�	�@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@���Lx�ٿ����n��@yc4@�+�ڐ�!?�k�T��@T��+Ηٿ����t��@"{7|�4@�2�n�!?3ؿc��@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@�Tj0l�ٿ*X̀���@d԰4@�o�i�!?������@a��۰�ٿ){�$�@��L��3@�g����!?۵dX��@a��۰�ٿ){�$�@��L��3@�g����!?۵dX��@a��۰�ٿ){�$�@��L��3@�g����!?۵dX��@a��۰�ٿ){�$�@��L��3@�g����!?۵dX��@a��۰�ٿ){�$�@��L��3@�g����!?۵dX��@�Ҷp�ٿ�ѣ���@�A�8� 4@K�Š�!?�װMoG�@�����ٿ��ҏ�t�@���4@�����!?�h�g�t�@�����ٿ��ҏ�t�@���4@�����!?�h�g�t�@���Ƕٿc�b���@,��ު4@�y��!?�-����@���Ƕٿc�b���@,��ު4@�y��!?�-����@���Ƕٿc�b���@,��ު4@�y��!?�-����@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@��:�`�ٿ&�+�۪�@�Tk� 4@��.iƏ!?9�S�<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@F��̷ٿ��/�0��@}�eJ�3@,��@�!?�_��t<�@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@��pذٿ���^t�@�����3@p�IՏ!?�ѻ��@�Sn��ٿ%����@M�� 4@���'֏!?B���A�@�Sn��ٿ%����@M�� 4@���'֏!?B���A�@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@o��h�ٿ�T�p�@eʺ�U 4@3���Q�!?½���@�h&�ٿV@�	���@Rz%� 4@�7K�!?�n��&�@�h&�ٿV@�	���@Rz%� 4@�7K�!?�n��&�@�h&�ٿV@�	���@Rz%� 4@�7K�!?�n��&�@�h&�ٿV@�	���@Rz%� 4@�7K�!?�n��&�@�h&�ٿV@�	���@Rz%� 4@�7K�!?�n��&�@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@+�ɓ��ٿ�`��%��@��s 4@�oc�̏!?ϴ��Z��@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@�(8���ٿ ������@1��c4@ �� ߏ!?\¨���@}�2׭�ٿ��^�@2��}N4@� �|�!?���b�>�@}�2׭�ٿ��^�@2��}N4@� �|�!?���b�>�@}�2׭�ٿ��^�@2��}N4@� �|�!?���b�>�@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@��3�ٿ���Z�@�t�
�4@� �>n�!?�|ù��@�~�/��ٿ�\JCFl�@������3@sK�^�!?�·�'��@�~�/��ٿ�\JCFl�@������3@sK�^�!?�·�'��@x��{,�ٿ�F��D�@(7�FD4@C�rJ5�!?�+���@x��{,�ٿ�F��D�@(7�FD4@C�rJ5�!?�+���@x��{,�ٿ�F��D�@(7�FD4@C�rJ5�!?�+���@x��{,�ٿ�F��D�@(7�FD4@C�rJ5�!?�+���@L�3m��ٿ���?W�@wr���4@gt ǲ�!?E��ۮ�@L�3m��ٿ���?W�@wr���4@gt ǲ�!?E��ۮ�@�r0��ٿ[Y���v�@�?�!D4@�b��ˏ!?&�ӛ��@�r0��ٿ[Y���v�@�?�!D4@�b��ˏ!?&�ӛ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�:ϲ��ٿ������@��T�- 4@�P�я!?/�� ��@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�D4-�ٿ�֜K�@���,n 4@��{��!?5����@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@�����ٿ�t;!$��@��P��3@�\8���!?�
���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@Ʒ�Οٿe<�Zh�@=�!pl 4@�^�+��!?�*iS���@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@��b.�ٿ.����@ڬ� 4@e ~T��!?�Z/P�@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@#��vȧٿ�]�z��@��i[��3@���8�!?	�D��@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@i	둤ٿiRn�4��@,��3@���y�!?Q��p���@��rU�ٿ�$ڼ�X�@0W�F�3@�g2B��!?��;�Z�@	m,V �ٿ��4z;�@���-��3@�DHҏ!?L����%�@	m,V �ٿ��4z;�@���-��3@�DHҏ!?L����%�@	m,V �ٿ��4z;�@���-��3@�DHҏ!?L����%�@	m,V �ٿ��4z;�@���-��3@�DHҏ!?L����%�@	m,V �ٿ��4z;�@���-��3@�DHҏ!?L����%�@C|�d��ٿ��q�!�@JA�4@�c�'܏!?���e�@C|�d��ٿ��q�!�@JA�4@�c�'܏!?���e�@-��R@�ٿV]&iQ�@�z¥��3@�o�d^�!?6��G��@�1��ٿg�"�[4�@p��/�3@�@����!?�>U�q�@U�Ȣٿ~i��=�@�)*(Q4@ς9͟�!?�g~_\Z�@U�Ȣٿ~i��=�@�)*(Q4@ς9͟�!?�g~_\Z�@U�Ȣٿ~i��=�@�)*(Q4@ς9͟�!?�g~_\Z�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@	��;ިٿ�wEP��@�$*�7 4@�dl���!?��D�Ġ�@1ŀ�o�ٿ�Z�2���@������3@�w|܏!?�\R�X�@1ŀ�o�ٿ�Z�2���@������3@�w|܏!?�\R�X�@1ŀ�o�ٿ�Z�2���@������3@�w|܏!?�\R�X�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@0���M�ٿ�.�	d�@�� .O 4@cZJ�!?����[�@F_��!�ٿ���d�@�y>>� 4@7�&7�!?x��}��@F_��!�ٿ���d�@�y>>� 4@7�&7�!?x��}��@F_��!�ٿ���d�@�y>>� 4@7�&7�!?x��}��@F_��!�ٿ���d�@�y>>� 4@7�&7�!?x��}��@F_��!�ٿ���d�@�y>>� 4@7�&7�!?x��}��@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@zS �ٿ8G�7ӧ�@D~Õ 4@Jʻv��!?����ɸ�@��@��ٿ\W�;_�@g��̒ 4@��
���!?!������@���Yܡٿ`sR���@����4@:4�<c�!?p& k�_�@���Yܡٿ`sR���@����4@:4�<c�!?p& k�_�@Pztt��ٿ�o���A�@��<X4@�zI���!?�W��"��@Pztt��ٿ�o���A�@��<X4@�zI���!?�W��"��@e��M�ٿ>�L����@I����4@V�*a�!?)��j�@�M�ٿK��]2��@MB� 4@ꒅ���!?��Q��@�M�ٿK��]2��@MB� 4@ꒅ���!?��Q��@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@Ƞ\��ٿxi��_��@F�K
 4@ҕɟ��!?:�׆O+�@��J��ٿoD=_L��@ z��� 4@��>�p�!?t�Da$��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@�7Y��ٿ\��?j�@X
!�3@BV �Տ!?��2D��@R�V���ٿ�m\�@��C���3@5 �U��!?[��<�@R�V���ٿ�m\�@��C���3@5 �U��!?[��<�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@ju�#�ٿ~��!;|�@��1߮ 4@��e{f�!?df׏I&�@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@����q�ٿ���I"��@S,�(� 4@�-�r�!?��aߌ��@i�ٵT�ٿ�[�3��@dmP���3@�X���!?������@i�ٵT�ٿ�[�3��@dmP���3@�X���!?������@��E=�ٿ�ǚ��@�jF�?�3@�Vaj�!?-����@��E=�ٿ�ǚ��@�jF�?�3@�Vaj�!?-����@�����ٿHǘ�@�3={e 4@�w/?��!?����o��@�����ٿHǘ�@�3={e 4@�w/?��!?����o��@��O�ٿ^�oH��@W��� 4@ʒ�(_�!?�4�Ytc�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@�n��ٿ
ě>���@(w�� 4@��W��!?>���@�@>�˘ٿ��7���@�t�U�4@NA���!?F1Z�n�@>�˘ٿ��7���@�t�U�4@NA���!?F1Z�n�@>�˘ٿ��7���@�t�U�4@NA���!?F1Z�n�@>�˘ٿ��7���@�t�U�4@NA���!?F1Z�n�@�2�⛟ٿ������@y�#�M4@i�/�!?վqM��@�2�⛟ٿ������@y�#�M4@i�/�!?վqM��@�2�⛟ٿ������@y�#�M4@i�/�!?վqM��@�2�⛟ٿ������@y�#�M4@i�/�!?վqM��@:��Ƹ�ٿ�� ���@>�"�4@1��z��!?��/���@Z��u�ٿ�����@|�W+4@ ����!?���o9C�@Z��u�ٿ�����@|�W+4@ ����!?���o9C�@Z��u�ٿ�����@|�W+4@ ����!?���o9C�@�eԫo�ٿ��w���@Ә`� 4@���U��!?�M�	 (�@�eԫo�ٿ��w���@Ә`� 4@���U��!?�M�	 (�@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@d��#�ٿ��-�G�@	f��4@����!?7����@3��b��ٿN&��%�@\�Q4@?�NRя!?{�艧�@_�M8i�ٿ5Dl�FN�@D��s�4@%�&f��!?&��T`�@_�M8i�ٿ5Dl�FN�@D��s�4@%�&f��!?&��T`�@_�M8i�ٿ5Dl�FN�@D��s�4@%�&f��!?&��T`�@�+�Y�ٿ��F���@��$R�4@Y�\鑏!?�$Ӕ4��@�+�Y�ٿ��F���@��$R�4@Y�\鑏!?�$Ӕ4��@�fB �ٿ�L�����@�{��u�3@K��ּ�!?O�G{Cm�@�fB �ٿ�L�����@�{��u�3@K��ּ�!?O�G{Cm�@�fB �ٿ�L�����@�{��u�3@K��ּ�!?O�G{Cm�@<����ٿ�S~ߝ�@�~Q��3@UU~'��!?ӱ!�Og�@<����ٿ�S~ߝ�@�~Q��3@UU~'��!?ӱ!�Og�@<����ٿ�S~ߝ�@�~Q��3@UU~'��!?ӱ!�Og�@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@������ٿp�>���@G�f8 4@F.S��!?,=Q���@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@���@�ٿ�WgC���@E��$�4@Z�0���!?���w��@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@�0ďt�ٿ����Nx�@3z�##4@O��ˏ!?"�/>l�@��"w�ٿj�.4��@��O�4@>濏!?=µ�E(�@��"w�ٿj�.4��@��O�4@>濏!?=µ�E(�@��"w�ٿj�.4��@��O�4@>濏!?=µ�E(�@��"w�ٿj�.4��@��O�4@>濏!?=µ�E(�@$�ʱϪٿ���O���@����4@� i�!?�,�t@��@$�ʱϪٿ���O���@����4@� i�!?�,�t@��@���ٿ��8?�X�@Q/��74@�X�`�!?�t~9��@���ٿ��8?�X�@Q/��74@�X�`�!?�t~9��@���ٿ��8?�X�@Q/��74@�X�`�!?�t~9��@���ٿ��8?�X�@Q/��74@�X�`�!?�t~9��@-a"�ȳٿDCZ!��@ۨϖ��3@�`0��!?d
��3��@-a"�ȳٿDCZ!��@ۨϖ��3@�`0��!?d
��3��@-a"�ȳٿDCZ!��@ۨϖ��3@�`0��!?d
��3��@-a"�ȳٿDCZ!��@ۨϖ��3@�`0��!?d
��3��@-a"�ȳٿDCZ!��@ۨϖ��3@�`0��!?d
��3��@��8u�ٿO�����@'0�I 4@���S�!?�4��M�@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@(ۥFe�ٿ%/�9s�@sz�/4@qb���!?���Ƴ��@���B��ٿ��9Y2��@���k4@^� cx�!?�#�R��@���B��ٿ��9Y2��@���k4@^� cx�!?�#�R��@���B��ٿ��9Y2��@���k4@^� cx�!?�#�R��@f����ٿ;�X�q�@&56;� 4@�JE'��!?���=��@f����ٿ;�X�q�@&56;� 4@�JE'��!?���=��@f����ٿ;�X�q�@&56;� 4@�JE'��!?���=��@f����ٿ;�X�q�@&56;� 4@�JE'��!?���=��@�eh8��ٿo���@��Lo�4@��=���!?�	�)��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@ӄ�/"�ٿg;��τ�@�K�$|4@��#p��!?ei�8��@w��O��ٿ=
�y�@�3�1H 4@��w] �!?06��@w��O��ٿ=
�y�@�3�1H 4@��w] �!?06��@w��O��ٿ=
�y�@�3�1H 4@��w] �!?06��@w��O��ٿ=
�y�@�3�1H 4@��w] �!?06��@w��O��ٿ=
�y�@�3�1H 4@��w] �!?06��@dx�[ҩٿj��z=F�@�c<^� 4@8��9֏!?b�s'.�@dx�[ҩٿj��z=F�@�c<^� 4@8��9֏!?b�s'.�@dx�[ҩٿj��z=F�@�c<^� 4@8��9֏!?b�s'.�@dx�[ҩٿj��z=F�@�c<^� 4@8��9֏!?b�s'.�@A3��ٿ(�����@&@$�V�3@w���Տ!?�)}8��@vm�E"�ٿ����/ �@�q�0��3@����!?D�m\�@T�"ɤ�ٿ?h�u%h�@��{�3@�����!?ʓFs�@T�"ɤ�ٿ?h�u%h�@��{�3@�����!?ʓFs�@T�"ɤ�ٿ?h�u%h�@��{�3@�����!?ʓFs�@T�"ɤ�ٿ?h�u%h�@��{�3@�����!?ʓFs�@T�"ɤ�ٿ?h�u%h�@��{�3@�����!?ʓFs�@Nd��ޝٿ���n�@k���3@;� ~�!?�1�*m��@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@ȞAe��ٿK��v`�@ĵm�� 4@'[�̡�!?����7[�@�����ٿm��'$��@b4��"�3@[�򒉏!?!�)�c�@�����ٿm��'$��@b4��"�3@[�򒉏!?!�)�c�@�����ٿm��'$��@b4��"�3@[�򒉏!?!�)�c�@�6\�ٿB��)�P�@���G�3@�Y漡�!?e�
S�@�6\�ٿB��)�P�@���G�3@�Y漡�!?e�
S�@�6\�ٿB��)�P�@���G�3@�Y漡�!?e�
S�@�u��ٿH�
��r�@<��f� 4@�V@�Ώ!?�������@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@!��h�ٿ
�"��3�@���q�3@��϶��!?*�7���@@�;Ğ�ٿ�0�z��@_�웻�3@�3�r`�!?�.2u���@@�;Ğ�ٿ�0�z��@_�웻�3@�3�r`�!?�.2u���@@�;Ğ�ٿ�0�z��@_�웻�3@�3�r`�!?�.2u���@@�;Ğ�ٿ�0�z��@_�웻�3@�3�r`�!?�.2u���@@�;Ğ�ٿ�0�z��@_�웻�3@�3�r`�!?�.2u���@VD�`ݧٿ胄Dg��@��� 4@/�D�d�!?��pE���@VD�`ݧٿ胄Dg��@��� 4@/�D�d�!?��pE���@VD�`ݧٿ胄Dg��@��� 4@/�D�d�!?��pE���@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�|5�4�ٿ����@�Q��4@�zu�p�!?䧊!'��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@�&�D�ٿŹV��@h{m�:4@�=&y�!?I2Uσ��@8�/�O�ٿ�ZŞ\*�@�y��3@$D�쾏!?|���ݾ�@8�/�O�ٿ�ZŞ\*�@�y��3@$D�쾏!?|���ݾ�@8�/�O�ٿ�ZŞ\*�@�y��3@$D�쾏!?|���ݾ�@8�/�O�ٿ�ZŞ\*�@�y��3@$D�쾏!?|���ݾ�@�Ǖ�ٿhp��fg�@��!d4�3@� ��!?�(����@��l^�ٿ��^��@S�LE�4@|@�h�!?IT�5��@�R��J�ٿ���2��@g��t`4@@����!?�
�.	�@�R��J�ٿ���2��@g��t`4@@����!?�
�.	�@�R��J�ٿ���2��@g��t`4@@����!?�
�.	�@��Lڤٿ��~�S��@~t�q4@�W����!?�{����@�Y8�ٿ�x3�@�9�(0 4@0�ѣ�!?�:�r1��@�Y8�ٿ�x3�@�9�(0 4@0�ѣ�!?�:�r1��@�ѿ�ٿ��$��@ �� 4@p�E�ď!?��rXoC�@�ѿ�ٿ��$��@ �� 4@p�E�ď!?��rXoC�@� �ʪٿ��:�n�@8�2�"4@P�|"�!?Y�/A�@$�\���ٿ�l�k^��@�p <a4@��Z��!?��E#:J�@$�\���ٿ�l�k^��@�p <a4@��Z��!?��E#:J�@$�\���ٿ�l�k^��@�p <a4@��Z��!?��E#:J�@$�\���ٿ�l�k^��@�p <a4@��Z��!?��E#:J�@�3���ٿ���ǩ�@�
�4@�`����!?����	w�@�i6�Z�ٿ'�MSj��@��M�4@7���L�!?A0M��@�i6�Z�ٿ'�MSj��@��M�4@7���L�!?A0M��@�i6�Z�ٿ'�MSj��@��M�4@7���L�!?A0M��@:S�ٿR��M�@ɶ��} 4@�(����!?k���)�@:S�ٿR��M�@ɶ��} 4@�(����!?k���)�@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@���B�ٿ�En��@���9 4@T_\F��!?�ֶr���@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@?��߭ٿ)b�^�i�@�#	�)�3@�%=!?js ����@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@iҟY�ٿN+��@��@���@��3@���=��!?�I�>�@r����ٿcyӌ�}�@q�8�> 4@ؒ����!?�ށ���@r����ٿcyӌ�}�@q�8�> 4@ؒ����!?�ށ���@r����ٿcyӌ�}�@q�8�> 4@ؒ����!?�ށ���@��թٿ�bJ����@�B R�3@���:�!?����,�@��թٿ�bJ����@�B R�3@���:�!?����,�@��թٿ�bJ����@�B R�3@���:�!?����,�@��թٿ�bJ����@�B R�3@���:�!?����,�@��թٿ�bJ����@�B R�3@���:�!?����,�@.�	�6�ٿ�ѣqH�@f����3@G�D#�!?��1ӈ�@.�	�6�ٿ�ѣqH�@f����3@G�D#�!?��1ӈ�@.�	�6�ٿ�ѣqH�@f����3@G�D#�!?��1ӈ�@.�	�6�ٿ�ѣqH�@f����3@G�D#�!?��1ӈ�@x�g�ӗٿ9��i��@!'��14@P�}ń�!?��-�M��@x�g�ӗٿ9��i��@!'��14@P�}ń�!?��-�M��@g����ٿ���ӕ�@/�4@�K�O��!?��I	���@g����ٿ���ӕ�@/�4@�K�O��!?��I	���@g����ٿ���ӕ�@/�4@�K�O��!?��I	���@g����ٿ���ӕ�@/�4@�K�O��!?��I	���@g����ٿ���ӕ�@/�4@�K�O��!?��I	���@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@�U�sN�ٿnv�s��@R�!9{4@E� �8�!?6K� >�@���@�ٿG^P���@���X.4@�ً�S�!?!����@���@�ٿG^P���@���X.4@�ً�S�!?!����@���@�ٿG^P���@���X.4@�ً�S�!?!����@�(�'��ٿ�� �E��@q��4@�?r�!?wZ���@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@� �ο�ٿ�0%��@"ߚE4@'��̘�!?�ctx%�@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@��͖?�ٿP�:c>��@��U��4@�jҏ!?A��a��@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@
 ��ٿ�S����@O�ث~ 4@�Iu���!?�^���6�@X����ٿ�R6�|�@<��2 4@f���E�!?w�/@��@X����ٿ�R6�|�@<��2 4@f���E�!?w�/@��@���I��ٿ��k�@؎�q� 4@��@R_�!?�E��a��@���I��ٿ��k�@؎�q� 4@��@R_�!?�E��a��@��o.`�ٿ�8QAę�@�9�Q��3@��D�׏!?�U����@TP���ٿ]pU>�@S���W4@�� C��!?�N](D�@TP���ٿ]pU>�@S���W4@�� C��!?�N](D�@Z=���ٿ��K�_�@�bb�$4@�@7��!?�>7F���@Z=���ٿ��K�_�@�bb�$4@�@7��!?�>7F���@Z=���ٿ��K�_�@�bb�$4@�@7��!?�>7F���@Z=���ٿ��K�_�@�bb�$4@�@7��!?�>7F���@iw�t��ٿڦ�����@'(i) 4@w����!?u�W���@iw�t��ٿڦ�����@'(i) 4@w����!?u�W���@�9f�ٿ��ja�i�@꧱"t�3@r���!?��j���@�9f�ٿ��ja�i�@꧱"t�3@r���!?��j���@�9f�ٿ��ja�i�@꧱"t�3@r���!?��j���@�9f�ٿ��ja�i�@꧱"t�3@r���!?��j���@�rmc>�ٿ��?-�9�@I��3@x� 	؏!?�����C�@�rmc>�ٿ��?-�9�@I��3@x� 	؏!?�����C�@�rmc>�ٿ��?-�9�@I��3@x� 	؏!?�����C�@�rmc>�ٿ��?-�9�@I��3@x� 	؏!?�����C�@� �@{�ٿ!G�!׷�@��ǃ?4@�:˜�!?[�̰���@� �@{�ٿ!G�!׷�@��ǃ?4@�:˜�!?[�̰���@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@-.��̩ٿ�5�y�@�I�{�4@�m�ӏ!?�k�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@I(ܞe�ٿ{��,��@�.	�z 4@ezy!?�v�ф8�@B|-���ٿ�h ]���@0Tdb 4@�Ŕ'[�!?1�ؕ��@B|-���ٿ�h ]���@0Tdb 4@�Ŕ'[�!?1�ؕ��@B|-���ٿ�h ]���@0Tdb 4@�Ŕ'[�!?1�ؕ��@��&>��ٿ_����@ � �4@� P�!?�ߥWc��@ъն�ٿ]��I���@S�-S��3@���i�!?�2��W��@HT��:�ٿ �^�@�y��( 4@ �Vb�!?@��
3�@HT��:�ٿ �^�@�y��( 4@ �Vb�!?@��
3�@HT��:�ٿ �^�@�y��( 4@ �Vb�!?@��
3�@HT��:�ٿ �^�@�y��( 4@ �Vb�!?@��
3�@HT��:�ٿ �^�@�y��( 4@ �Vb�!?@��
3�@�Wbh�ٿ�[�qK�@�2��� 4@�� 颏!?�gf����@�Wbh�ٿ�[�qK�@�2��� 4@�� 颏!?�gf����@�Wbh�ٿ�[�qK�@�2��� 4@�� 颏!?�gf����@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@_A��7�ٿĀ.��2�@֒Z@4@sm�ӏ!?�8�@��w.�ٿ����@���4@,�r�!?����+	�@��w.�ٿ����@���4@,�r�!?����+	�@r�٭��ٿ�ٝw��@8�t�4@�iVg�!?�8>3Q��@�q �B�ٿ���)b@�@��qE� 4@�b2��!?�5ag(�@��.I��ٿt�&É1�@��m�4@�{D[�!?���W�@��.I��ٿt�&É1�@��m�4@�{D[�!?���W�@���d��ٿ��}��@�
( 4@.Z+P1�!?c�����@���d��ٿ��}��@�
( 4@.Z+P1�!?c�����@���d��ٿ��}��@�
( 4@.Z+P1�!?c�����@^L���ٿ�1���	�@�k"��3@g��V�!?X�����@�
��ٿ'1v[w��@_۫���3@D}B�!?���O�@�
��ٿ'1v[w��@_۫���3@D}B�!?���O�@~��ٿEË]�c�@T߼��3@��e��!?[]!Ḉ�@~��ٿEË]�c�@T߼��3@��e��!?[]!Ḉ�@~��ٿEË]�c�@T߼��3@��e��!?[]!Ḉ�@~��ٿEË]�c�@T߼��3@��e��!?[]!Ḉ�@^.VQ�ٿ����׾�@'�ѡF�3@��~Ţ�!?�ʗ��5�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@Xo"L�ٿ�uL���@
8Y?W�3@M�2���!?���׀�@���k�ٿ�P���U�@�P/�4@�D����!?�-���@�rFx�ٿ�} ���@��ɮ�4@��n�!?j�@�@�rFx�ٿ�} ���@��ɮ�4@��n�!?j�@�@Ѣ�W�ٿ��:3*s�@���F,4@�ż�u�!?@ڋ�s�@j��ҏ�ٿ.4��@�V�Ǝ4@�*�	��!?k43�GJ�@j��ҏ�ٿ.4��@�V�Ǝ4@�*�	��!?k43�GJ�@j��ҏ�ٿ.4��@�V�Ǝ4@�*�	��!?k43�GJ�@��?^�ٿEʵ��Z�@�ы* 4@M��f��!?|���@��?^�ٿEʵ��Z�@�ы* 4@M��f��!?|���@��?^�ٿEʵ��Z�@�ы* 4@M��f��!?|���@��?^�ٿEʵ��Z�@�ы* 4@M��f��!?|���@���G�ٿ��g���@�%����3@=%"�c�!?2h����@���G�ٿ��g���@�%����3@=%"�c�!?2h����@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@+���ٿ�Z�O���@����*�3@�(��V�!?�WH�P��@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@)���ٿ|�캖��@��M��3@�*U��!?����@�8<�ĦٿF�3���@�v-t4@��:Y�!?5~�:+�@���}�ٿ�ԡ{��@�oy�/4@yr5I��!?	G��9�@���}�ٿ�ԡ{��@�oy�/4@yr5I��!?	G��9�@���}�ٿ�ԡ{��@�oy�/4@yr5I��!?	G��9�@���}�ٿ�ԡ{��@�oy�/4@yr5I��!?	G��9�@L���ٿz`]@��@h�� 4@�˝e�!?����@L���ٿz`]@��@h�� 4@�˝e�!?����@hs�9^�ٿ�)��@�2n���3@�4H�!?��e�}o�@f�I�Y�ٿ�{����@��l7�3@Y]��(�!?Y���#�@f�I�Y�ٿ�{����@��l7�3@Y]��(�!?Y���#�@|�h1+�ٿO��W`�@H9h�y 4@��롪�!?c�����@|�h1+�ٿO��W`�@H9h�y 4@��롪�!?c�����@|�h1+�ٿO��W`�@H9h�y 4@��롪�!?c�����@����ͧٿ�u���(�@�*Ԩ� 4@�8+ߏ!?�\C���@����ͧٿ�u���(�@�*Ԩ� 4@�8+ߏ!?�\C���@����ͧٿ�u���(�@�*Ԩ� 4@�8+ߏ!?�\C���@��0�ٿ�XV��'�@��I4@)J3��!?��<�@��0�ٿ�XV��'�@��I4@)J3��!?��<�@x�U�ٿ�H(���@�w���3@�i�ҏ!?ӌ&�8u�@x�U�ٿ�H(���@�w���3@�i�ҏ!?ӌ&�8u�@D��~"�ٿbv�`�@����, 4@���؏!?H�&��@D��~"�ٿbv�`�@����, 4@���؏!?H�&��@D��~"�ٿbv�`�@����, 4@���؏!?H�&��@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@��__'�ٿ9���R��@�jE� 4@i��ȏ!?�t��"�@R �E��ٿ������@��h�S�3@���؏!?*4WƷ�@R �E��ٿ������@��h�S�3@���؏!?*4WƷ�@,d9()�ٿi=-<Y�@�R�WD4@��fR��!?BE�S��@,d9()�ٿi=-<Y�@�R�WD4@��fR��!?BE�S��@,d9()�ٿi=-<Y�@�R�WD4@��fR��!?BE�S��@�Je�ٿ��D�5�@����4@�3�7��!?m��K�@�Je�ٿ��D�5�@����4@�3�7��!?m��K�@�Je�ٿ��D�5�@����4@�3�7��!?m��K�@�Je�ٿ��D�5�@����4@�3�7��!?m��K�@�G��m�ٿ�dC��@�}.��3@U	<k�!?:*�;��@�G��m�ٿ�dC��@�}.��3@U	<k�!?:*�;��@�G��m�ٿ�dC��@�}.��3@U	<k�!?:*�;��@�G��m�ٿ�dC��@�}.��3@U	<k�!?:*�;��@�G��m�ٿ�dC��@�}.��3@U	<k�!?:*�;��@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@����}�ٿ��w=���@������3@u�9�Ï!?4�3' �@��E��ٿ��pݕ�@C�w� 4@N�r�!?��jJx0�@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@��a���ٿ+�0�C��@��~�3@�4.[ɏ!?�1 ��@�y�Φ�ٿD��q��@��:�P 4@�����!?dW�HV�@�y�Φ�ٿD��q��@��:�P 4@�����!?dW�HV�@�y�Φ�ٿD��q��@��:�P 4@�����!?dW�HV�@�y�Φ�ٿD��q��@��:�P 4@�����!?dW�HV�@'�Uӯ�ٿ�A�g��@Z����3@�m
в�!?$��@'�Uӯ�ٿ�A�g��@Z����3@�m
в�!?$��@�D�0=�ٿ�<J���@�U[��3@�̘`�!?�Ѷcf�@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@n�Mm>�ٿ�nĝN�@�~V!B�3@A�﯏!?wQ�fM��@(3����ٿL���@зAT�3@@<8P��!?z�t�5��@(3����ٿL���@зAT�3@@<8P��!?z�t�5��@(3����ٿL���@зAT�3@@<8P��!?z�t�5��@�0�s�ٿ�ࢢ�-�@����3@�����!?�W�j�L�@�0�s�ٿ�ࢢ�-�@����3@�����!?�W�j�L�@����ٿ�H$�ǒ�@�	BKr�3@�+5��!?k����@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@��:�ٿ?�,�[��@"�;���3@#��$�!?B~(H5��@`�{�t�ٿ����C��@FӲ���3@��!?Ц˰*�@`�{�t�ٿ����C��@FӲ���3@��!?Ц˰*�@?F�i�ٿ�M3����@�ɔU��3@�����!?g�s��S�@?F�i�ٿ�M3����@�ɔU��3@�����!?g�s��S�@[�Q�ٿ������@������3@�Dm�Ǐ!?�O�;��@[�Q�ٿ������@������3@�Dm�Ǐ!?�O�;��@[�Q�ٿ������@������3@�Dm�Ǐ!?�O�;��@[�Q�ٿ������@������3@�Dm�Ǐ!?�O�;��@ڸ�#;�ٿ-�<ĝx�@ΛDG� 4@�Z�я!?Ӑ�q��@ڸ�#;�ٿ-�<ĝx�@ΛDG� 4@�Z�я!?Ӑ�q��@6}��ۨٿ�Y�O��@�sw��3@�`L��!?�����@6}��ۨٿ�Y�O��@�sw��3@�`L��!?�����@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@���ٿ1y�p�K�@���r�3@x�+_��!?B��K�@-fe�ٿ��Fp�@t%��u 4@�`-�!?�&=u�@-fe�ٿ��Fp�@t%��u 4@�`-�!?�&=u�@T�kҞٿW����@���Q�4@�{ =�!?���\�@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@p��#�ٿa�"ً��@d�H�N 4@��K�ޏ!?2�O"��@�gC�;�ٿT�34��@��q�4@	E̏!?�
���@�gC�;�ٿT�34��@��q�4@	E̏!?�
���@�gC�;�ٿT�34��@��q�4@	E̏!?�
���@�gC�;�ٿT�34��@��q�4@	E̏!?�
���@��-M��ٿ�4Ǘ��@8�)� 4@����V�!?��O���@��-M��ٿ�4Ǘ��@8�)� 4@����V�!?��O���@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@92��˒ٿ� &e���@Wm�g� 4@��w�~�!?���f��@w��1��ٿ0��{�@�F>S 4@W_�[ڏ!?2�v�!��@w��1��ٿ0��{�@�F>S 4@W_�[ڏ!?2�v�!��@��+*�ٿVʦ�a-�@��h)4@%Fs�!?y���o�@��sJ��ٿo��C��@d�㫩 4@��n �!?Ϋ��uS�@�SED�ٿ���
�g�@�U��4@�_u��!?�Y>�{��@�SED�ٿ���
�g�@�U��4@�_u��!?�Y>�{��@�SED�ٿ���
�g�@�U��4@�_u��!?�Y>�{��@n�^�ٿV�}�X.�@.j��l4@���܏!?D����@n�^�ٿV�}�X.�@.j��l4@���܏!?D����@n�^�ٿV�}�X.�@.j��l4@���܏!?D����@n�^�ٿV�}�X.�@.j��l4@���܏!?D����@n�^�ٿV�}�X.�@.j��l4@���܏!?D����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@�87�C�ٿ���]7j�@��{1 4@�SV�!?V ����@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@Nb?��ٿ@��R��@���� 4@+�rJ��!?����g�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�MJ(�ٿ(M�<��@�F9$ 4@ޑ��i�!?�O}�@�+R�'�ٿcg�"��@à���3@��t'�!?���G��@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@3�ȣΡٿUۭxz��@��[� 4@��m6�!?Ʈ�� �@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@
�����ٿ(q[�@�@�3P�3@�c9[��!?�
s�@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@zCF��ٿT]���@�#���4@�3��x�!?��_���@sOHW��ٿ��,��@�/bSE 4@rb�!?�	�ͯ��@sOHW��ٿ��,��@�/bSE 4@rb�!?�	�ͯ��@�@X�ٿ��H�1��@�o"�4@��d��!?{<��}Q�@|�˯M�ٿ�������@�ӻc�4@�H�&��!?{��>i�@��#�P�ٿ�����@i�&) 4@����!?���Cd��@��#�P�ٿ�����@i�&) 4@����!?���Cd��@��#�P�ٿ�����@i�&) 4@����!?���Cd��@��#�P�ٿ�����@i�&) 4@����!?���Cd��@��#�P�ٿ�����@i�&) 4@����!?���Cd��@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@T�{$-�ٿ�a:@�7�@�a"�E�3@�<4��!?֛���[�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@������ٿS}��y.�@y��\G 4@��)iӏ!?K���3�@�5��J�ٿ'\�M6^�@$F�X4@9"ʎ�!?�3b�p�@�5��J�ٿ'\�M6^�@$F�X4@9"ʎ�!?�3b�p�@�5��J�ٿ'\�M6^�@$F�X4@9"ʎ�!?�3b�p�@P�*>�ٿ,�^"��@%�T�h4@��o��!?�,���@P�*>�ٿ,�^"��@%�T�h4@��o��!?�,���@P�*>�ٿ,�^"��@%�T�h4@��o��!?�,���@�Uz7��ٿ6<�J�^�@2J�Ռ4@�C�!?�{?^Ή�@�Uz7��ٿ6<�J�^�@2J�Ռ4@�C�!?�{?^Ή�@�Uz7��ٿ6<�J�^�@2J�Ռ4@�C�!?�{?^Ή�@�Uz7��ٿ6<�J�^�@2J�Ռ4@�C�!?�{?^Ή�@(�ǽ��ٿ�~[����@�"���4@	�K�!?���u���@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@8�����ٿƠ$�P	�@�NO���3@�u^ꪏ!?6�H��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@h0�Q�ٿז�(I��@��n�3@�
�ŏ!?�-��k��@f$��ٿ{�Cz%��@������3@&N�I��!?�O�<2��@f$��ٿ{�Cz%��@������3@&N�I��!?�O�<2��@f$��ٿ{�Cz%��@������3@&N�I��!?�O�<2��@f$��ٿ{�Cz%��@������3@&N�I��!?�O�<2��@f$��ٿ{�Cz%��@������3@&N�I��!?�O�<2��@�ēy�ٿW3�����@L��! 4@?���!?E�cG�@�ēy�ٿW3�����@L��! 4@?���!?E�cG�@8u�6��ٿk�Ph��@Q��7� 4@���ah�!?������@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@���̜ٿ�Ӽ�F~�@�FO� 4@�R݃�!?PIG�n��@��\rǥٿ�0�J�@��N��3@�'G⪏!?ZI?�@)��ٿ�������@� ����3@ݤb�!?�GI����@a�G�D�ٿ�XO��6�@u�����3@!�x���!?Ժ#̹�@a�G�D�ٿ�XO��6�@u�����3@!�x���!?Ժ#̹�@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�g���ٿ����ޙ�@R8$��3@�t�!?�0L2���@�y��ٿ��W�m�@�,�&�3@�!%뛏!?��/���@�y��ٿ��W�m�@�,�&�3@�!%뛏!?��/���@�y��ٿ��W�m�@�,�&�3@�!%뛏!?��/���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@h|)���ٿ��!1X�@ @�S��3@���!�!?�0�s���@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@�U��ٿb����@��՗�4@�u��!?rh����@��у��ٿ|D�_,��@�6���4@zR�冏!?����^�@��у��ٿ|D�_,��@�6���4@zR�冏!?����^�@�S���ٿ�\�C��@���r�3@����!?�E�Q�@�S���ٿ�\�C��@���r�3@����!?�E�Q�@ J7C�ٿhb)��@�G�U��3@G�J(ˏ!?jcKI�@o�vv�ٿ~��a��@=Ú4@mo��!?i���@o�vv�ٿ~��a��@=Ú4@mo��!?i���@.�avȸٿ#�yf��@��97g 4@���P׏!?�aR=� �@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@ :g���ٿ=ܹG�&�@{���� 4@E���n�!?�s�F���@�&���ٿw�w����@5	%s�4@��
s��!?5�U�@�&���ٿw�w����@5	%s�4@��
s��!?5�U�@�&���ٿw�w����@5	%s�4@��
s��!?5�U�@�&���ٿw�w����@5	%s�4@��
s��!?5�U�@��R�ٿ�O�����@<�X � 4@�9�Ԗ�!?*��l
�@�Ý���ٿ������@~��X��3@�c�܌�!?�܆��o�@�Ý���ٿ������@~��X��3@�c�܌�!?�܆��o�@ì�C�ٿ���!nQ�@��[�( 4@���U�!?C?V�b��@ì�C�ٿ���!nQ�@��[�( 4@���U�!?C?V�b��@ì�C�ٿ���!nQ�@��[�( 4@���U�!?C?V�b��@ì�C�ٿ���!nQ�@��[�( 4@���U�!?C?V�b��@�OV.�ٿW�l��@�Աڻ�3@a��_4�!?L��.�4�@ :[�W�ٿ�z�u���@����# 4@�E�o�!?���"3�@ :[�W�ٿ�z�u���@����# 4@�E�o�!?���"3�@����ٿ�Z��q�@=�H��3@s<�y�!?�l����@�A7��ٿ@N�H'l�@`�G� 4@���M�!?��m�Uc�@�A7��ٿ@N�H'l�@`�G� 4@���M�!?��m�Uc�@�A7��ٿ@N�H'l�@`�G� 4@���M�!?��m�Uc�@Tg|=�ٿ����P��@˦�@�4@�k���!?~�5g!��@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@��%��ٿ�1D�	�@­�&� 4@���ɏ!?�M��+�@���ٿLmz�V�@���g�3@���؏!?-6�LH��@���ٿLmz�V�@���g�3@���؏!?-6�LH��@���ٿLmz�V�@���g�3@���؏!?-6�LH��@��91ɡٿLM�u!>�@խ��e4@��Do�!?}�K��@��91ɡٿLM�u!>�@խ��e4@��Do�!?}�K��@��91ɡٿLM�u!>�@խ��e4@��Do�!?}�K��@��91ɡٿLM�u!>�@խ��e4@��Do�!?}�K��@D����ٿ0;�Q��@o`���4@m6�uf�!?4�4}��@D����ٿ0;�Q��@o`���4@m6�uf�!?4�4}��@D����ٿ0;�Q��@o`���4@m6�uf�!?4�4}��@D����ٿ0;�Q��@o`���4@m6�uf�!?4�4}��@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@�՞®ٿ��*R��@���v�4@��*���!?�4����@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��N_��ٿ��ǿ)�@����4@4+�ُ!?��*%5�@��D~��ٿ�o��A�@�١�4@��%��!?'�)!�@��D~��ٿ�o��A�@�١�4@��%��!?'�)!�@��D~��ٿ�o��A�@�١�4@��%��!?'�)!�@��D~��ٿ�o��A�@�١�4@��%��!?'�)!�@��D~��ٿ�o��A�@�١�4@��%��!?'�)!�@��|�ٿ�h���@�皺� 4@�����!?���t��@��|�ٿ�h���@�皺� 4@�����!?���t��@��|�ٿ�h���@�皺� 4@�����!?���t��@�T�3�ٿC��@v��@�F�� 4@��/厏!? �Z���@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�j�ѵٿ���m��@��� z 4@Q��S��!?0�Q�v�@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@�Ed�ٿ�?jq��@]$�7�4@-�����!?��?��@r���G�ٿ��f�M��@U)�	�4@��[�!?l�w�@�3��ٿ�X�g;�@�w|W4@[马k�!?O5Կ=w�@�3��ٿ�X�g;�@�w|W4@[马k�!?O5Կ=w�@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@��PZ�ٿ�L�k���@y,��4@�7�Z�!?lC����@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@b��ٿ�2���@Kr�շ 4@/��EG�!?������@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@����|�ٿ"�3|���@h�W� 4@�����!?_[��a�@���S~�ٿ�������@!Q�4@��K*I�!?Hu�>�S�@���\P�ٿ�935���@��^�> 4@��꩏!?���L&f�@%P�E�ٿ�զ�ɍ�@:��ܺ�3@�b����!?Pn�N�i�@	�`�ٿ�h�����@����� 4@i��ҏ!?�n{���@	�`�ٿ�h�����@����� 4@i��ҏ!?�n{���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@��ѢW�ٿ��g�b��@��M�� 4@z:�O��!?�+cb���@�m� �ٿ��_{b��@�Xg��3@���w�!?Ke�_���@�m� �ٿ��_{b��@�Xg��3@���w�!?Ke�_���@�)�鎭ٿw����@��;���3@	�hď!?��0�z�@;npk��ٿ& �_��@;����3@%�D��!?@'L����@;npk��ٿ& �_��@;����3@%�D��!?@'L����@;npk��ٿ& �_��@;����3@%�D��!?@'L����@;npk��ٿ& �_��@;����3@%�D��!?@'L����@;npk��ٿ& �_��@;����3@%�D��!?@'L����@;npk��ٿ& �_��@;����3@%�D��!?@'L����@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@�����ٿ��]��@����Z4@��Un�!?�-?�i��@9�}�f�ٿD0����@���� 4@��w���!?�l�?�@9�}�f�ٿD0����@���� 4@��w���!?�l�?�@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@A�Q��ٿ�Um`�(�@�����3@�;����!?���fW��@]\�,�ٿ� 2���@��A: 4@1f���!?����@]\�,�ٿ� 2���@��A: 4@1f���!?����@�哉{�ٿ�7D���@S^ټ�3@��9C��!?4q�鳱�@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@n���e�ٿ��H�j��@���4� 4@0�T���!?��]���@����ٿzjR���@у����3@"���!?�똬��@���ٿ��j���@OG����3@����!?��52�@���ٿ��j���@OG����3@����!?��52�@���ٿ��j���@OG����3@����!?��52�@���ٿ��j���@OG����3@����!?��52�@���ٿ��j���@OG����3@����!?��52�@���ٿ��j���@OG����3@����!?��52�@΢�ٿ�ٿ@B�	S�@�&亐�3@�����!?��'i���@΢�ٿ�ٿ@B�	S�@�&亐�3@�����!?��'i���@΢�ٿ�ٿ@B�	S�@�&亐�3@�����!?��'i���@΢�ٿ�ٿ@B�	S�@�&亐�3@�����!?��'i���@XT`�ٿ�?R��	�@6�>���3@H�h�ݏ!?���߆(�@XT`�ٿ�?R��	�@6�>���3@H�h�ݏ!?���߆(�@��Q�ٿ�B���M�@X��X�3@y�駏!?7�W�50�@��Q�ٿ�B���M�@X��X�3@y�駏!?7�W�50�@��Q�ٿ�B���M�@X��X�3@y�駏!?7�W�50�@��Q�ٿ�B���M�@X��X�3@y�駏!?7�W�50�@M�{���ٿS�5 ��@�Z���3@aP��Ώ!?�FP�[�@M�{���ٿS�5 ��@�Z���3@aP��Ώ!?�FP�[�@V� ,H�ٿ�z4y�b�@�ߢ9� 4@؀aO��!?K�e?F��@�(+��ٿM �_�@M�K�4@/�ď!?�V�����@�(+��ٿM �_�@M�K�4@/�ď!?�V�����@�(+��ٿM �_�@M�K�4@/�ď!?�V�����@�(+��ٿM �_�@M�K�4@/�ď!?�V�����@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@[���ٿ'(��~?�@Q���4@�'`��!?OI}'�8�@��2���ٿၸ�Af�@���B 4@0�Tܱ�!?����%�@��2���ٿၸ�Af�@���B 4@0�Tܱ�!?����%�@��2���ٿၸ�Af�@���B 4@0�Tܱ�!?����%�@��2���ٿၸ�Af�@���B 4@0�Tܱ�!?����%�@���yW�ٿ4N���_�@L3M84@3�܄r�!?�E<c�@���yW�ٿ4N���_�@L3M84@3�܄r�!?�E<c�@���yW�ٿ4N���_�@L3M84@3�܄r�!?�E<c�@���yW�ٿ4N���_�@L3M84@3�܄r�!?�E<c�@���yW�ٿ4N���_�@L3M84@3�܄r�!?�E<c�@f�,쑜ٿi�-(��@f��4@�͐��!?"����@f�,쑜ٿi�-(��@f��4@�͐��!?"����@f�,쑜ٿi�-(��@f��4@�͐��!?"����@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@��ѣx�ٿ��o@���@G:@�4@Gy#J׏!?<�xx��@�13N��ٿ��/��@�r�4@-��p�!?����@�13N��ٿ��/��@�r�4@-��p�!?����@�13N��ٿ��/��@�r�4@-��p�!?����@�13N��ٿ��/��@�r�4@-��p�!?����@��X�W�ٿbm!��@ש� 4@#�,��!?��Bn���@��X�W�ٿbm!��@ש� 4@#�,��!?��Bn���@Tr�>:�ٿ$�,A���@�����3@a����!?G�����@Tr�>:�ٿ$�,A���@�����3@a����!?G�����@Tr�>:�ٿ$�,A���@�����3@a����!?G�����@Tr�>:�ٿ$�,A���@�����3@a����!?G�����@Tr�>:�ٿ$�,A���@�����3@a����!?G�����@�*Ɓ�ٿRSS���@f`�g44@d�y��!?8�-^���@�*Ɓ�ٿRSS���@f`�g44@d�y��!?8�-^���@�*Ɓ�ٿRSS���@f`�g44@d�y��!?8�-^���@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@KF�}��ٿ@��?�@���U��3@Ld���!?����@)W�h��ٿg��tPk�@��94@2,|���!?�)�P��@�Nŉ��ٿC��5�8�@կ�. 4@C��N��!?"b�D��@�Nŉ��ٿC��5�8�@կ�. 4@C��N��!?"b�D��@�Nŉ��ٿC��5�8�@կ�. 4@C��N��!?"b�D��@i��'E�ٿC��?�j�@|�j 4@���K��!?�M����@�&Y^�ٿ��%�B0�@�Vm���3@�+�/��!?�H$��c�@���L��ٿv�?@%1�@|� ��3@)h�w��!?X�/V?��@�l�ZI�ٿ$뚧�)�@���5��3@2�����!?�u��T�@�l�ZI�ٿ$뚧�)�@���5��3@2�����!?�u��T�@�l�ZI�ٿ$뚧�)�@���5��3@2�����!?�u��T�@�l�ZI�ٿ$뚧�)�@���5��3@2�����!?�u��T�@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@��&7�ٿ[�TA�@���>@4@��)]t�!?���T��@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@�����ٿ :�� ��@l>�:4@�:��x�!?F�(�ĺ�@���ڥٿ1u�u���@U��h 4@�L����!?Tt�M���@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@fkf�ٿyg���N�@H�:�� 4@�o��͏!?(Bj��@[gx賩ٿ,*��p�@�H��V 4@A�S��!?�(����@[gx賩ٿ,*��p�@�H��V 4@A�S��!?�(����@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��m�D�ٿX��%�@�%k�4@�Wl���!?[ԩV�8�@��E6�ٿ�r)��@r�� 4@?W_Ϗ!?��Ì���@n����ٿ�E�E7Y�@�lR 4@F�s�u�!?��<L�@n����ٿ�E�E7Y�@�lR 4@F�s�u�!?��<L�@eZ�#�ٿ�{Ƌ?�@>��N��3@�Sϧy�!?'	m���@eZ�#�ٿ�{Ƌ?�@>��N��3@�Sϧy�!?'	m���@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@@�|��ٿ������@f�7��3@��~w�!?s>��/�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�^/�ٿ��_�7�@s3�B�3@�����!?��(rI$�@�KhU�ٿ��҈K�@���9@�3@��]��!?&.Z�>'�@�F��N�ٿ-�=�ye�@~�% 4@ߖ����!?��*�Y�@ރg�F�ٿ����k�@k��-� 4@E��Ǐ!?n"� hz�@ރg�F�ٿ����k�@k��-� 4@E��Ǐ!?n"� hz�@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@ӄ�R[�ٿ/�h3��@OUb���3@��$ʏ!??fԂn��@����ٿ*{"�lu�@W�3 ~ 4@��[v�!?������@����ٿ*{"�lu�@W�3 ~ 4@��[v�!?������@��L��ٿiI688t�@���;4@5���ӏ!?!p�8���@��L��ٿiI688t�@���;4@5���ӏ!?!p�8���@��L��ٿiI688t�@���;4@5���ӏ!?!p�8���@�#�W�ٿ)S����@���4@���䈏!?��p���@��g�ٿޱILp�@�t��4@�}:�!?34�{L �@��g�ٿޱILp�@�t��4@�}:�!?34�{L �@��g�ٿޱILp�@�t��4@�}:�!?34�{L �@��g�ٿޱILp�@�t��4@�}:�!?34�{L �@�^t�b�ٿ�bv>e�@���F�3@��lE�!?Uv�����@�^t�b�ٿ�bv>e�@���F�3@��lE�!?Uv�����@�wu	�ٿ�-�S�@���%�3@W}�!?��"%�:�@�^���ٿ���B�X�@�&��s�3@:r����!?�R��v�@�!�%I�ٿbz�.E�@���) 4@e
�%Ώ!?<�v���@�!�%I�ٿbz�.E�@���) 4@e
�%Ώ!?<�v���@�!�%I�ٿbz�.E�@���) 4@e
�%Ώ!?<�v���@�!�%I�ٿbz�.E�@���) 4@e
�%Ώ!?<�v���@�!�%I�ٿbz�.E�@���) 4@e
�%Ώ!?<�v���@�ߊLk�ٿ,�Tn�@>�w�� 4@ߡ�頏!?�{�9 ;�@�ߊLk�ٿ,�Tn�@>�w�� 4@ߡ�頏!?�{�9 ;�@�ߊLk�ٿ,�Tn�@>�w�� 4@ߡ�頏!?�{�9 ;�@p�Y6N�ٿ^-?�!��@���V 4@od�j�!?�D��]�@��6���ٿVT'�@�&�=[4@0L���!?����e�@���ٿr���N�@4�@�`�3@�v�.ˏ!?�#���+�@���ٿr���N�@4�@�`�3@�v�.ˏ!?�#���+�@Gi��֞ٿ"�U�R��@��	F4@�<D���!?wv�5-�@Gi��֞ٿ"�U�R��@��	F4@�<D���!?wv�5-�@Gi��֞ٿ"�U�R��@��	F4@�<D���!?wv�5-�@Gi��֞ٿ"�U�R��@��	F4@�<D���!?wv�5-�@Gi��֞ٿ"�U�R��@��	F4@�<D���!?wv�5-�@?�x�L�ٿinX�1��@�DS� 4@npT蒏!?�ecg��@�" ��ٿ��4!�s�@d��iJ4@rx�a��!?��Z�6�@|��g*�ٿp�)�P��@�|�P�3@� 8>�!?ۖ" ��@|��g*�ٿp�)�P��@�|�P�3@� 8>�!?ۖ" ��@|��g*�ٿp�)�P��@�|�P�3@� 8>�!?ۖ" ��@�*���ٿ�*����@=�_��3@<Zf<d�!?	Z��R��@�*���ٿ�*����@=�_��3@<Zf<d�!?	Z��R��@�*���ٿ�*����@=�_��3@<Zf<d�!?	Z��R��@aq�Y�ٿ>�v��@׿���3@� ֯t�!?�K
0���@aq�Y�ٿ>�v��@׿���3@� ֯t�!?�K
0���@aq�Y�ٿ>�v��@׿���3@� ֯t�!?�K
0���@2��'�ٿ����@ ��� 4@HⲎ��!?�^�d:E�@	m{J�ٿ��u* ��@g��HV�3@c�R��!?��0_|�@#�y�ٿ�-��zy�@p'��3@uN�WK�!?�V CW��@#�y�ٿ�-��zy�@p'��3@uN�WK�!?�V CW��@#�y�ٿ�-��zy�@p'��3@uN�WK�!?�V CW��@��r�ٿ�ٔ��@��J# 4@��҇��!?$_���@��yl*�ٿ�]Ad���@ ����3@�c���!?�&�i�N�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@�o��ٿ�/e��@;NF;� 4@\�����!?.F�㤁�@#��V�ٿ�����@�2xL?4@�����!?�+Jl2��@#��V�ٿ�����@�2xL?4@�����!?�+Jl2��@#��V�ٿ�����@�2xL?4@�����!?�+Jl2��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@��M��ٿ��C.�@;ω��4@Pm�]��!?Pm�ԥ��@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@�����ٿ�C�Y�@��@S4@v�׶�!?�lZ���@8?����ٿ�����@:� Js4@R�ɩ�!?��<���@M:��ٿ`+�XA�@�mTb� 4@�{"ǲ�!?6����@M:��ٿ`+�XA�@�mTb� 4@�{"ǲ�!?6����@M:��ٿ`+�XA�@�mTb� 4@�{"ǲ�!?6����@s�EFO�ٿt������@@�0{4@�=�Ϗ!?>�wN<4�@s�EFO�ٿt������@@�0{4@�=�Ϗ!?>�wN<4�@���X��ٿ��=�$��@w�wI�4@ݫCyȏ!?S� 
���@����ٿ�
�3�@��� 4@�}.\��!?V�����@i=gњ�ٿ�8V3�@��C� 4@��'O�!?�t	�2�@i=gњ�ٿ�8V3�@��C� 4@��'O�!?�t	�2�@i=gњ�ٿ�8V3�@��C� 4@��'O�!?�t	�2�@i=gњ�ٿ�8V3�@��C� 4@��'O�!?�t	�2�@i=gњ�ٿ�8V3�@��C� 4@��'O�!?�t	�2�@�X�7�ٿ���J,��@�AF�N 4@T���!?�@!4x�@�X�7�ٿ���J,��@�AF�N 4@T���!?�@!4x�@�X�7�ٿ���J,��@�AF�N 4@T���!?�@!4x�@�X�7�ٿ���J,��@�AF�N 4@T���!?�@!4x�@��2�6�ٿ�;�`~�@�?��4@ ��B��!?�س� �@��2�6�ٿ�;�`~�@�?��4@ ��B��!?�س� �@�����ٿ���Ȗ�@�\�'4@��6:̏!?�\����@�����ٿ���Ȗ�@�\�'4@��6:̏!?�\����@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@	/�]�ٿ+��}�F�@�G�4@�{7l��!?ѝB�?�@��#f�ٿ�#V�g�@��6�4@��޴��!?�P����@I{G��ٿ�κʴ�@8&�'4@M� R��!?T������@I{G��ٿ�κʴ�@8&�'4@M� R��!?T������@I{G��ٿ�κʴ�@8&�'4@M� R��!?T������@:d�[t�ٿ�*�����@T�R��4@�NN�n�!?�܂a���@:d�[t�ٿ�*�����@T�R��4@�NN�n�!?�܂a���@:d�[t�ٿ�*�����@T�R��4@�NN�n�!?�܂a���@:d�[t�ٿ�*�����@T�R��4@�NN�n�!?�܂a���@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@.�5�ٿ]�S&�@��D��4@�-x�r�!?N�S�'�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@ O�L�ٿ?��cA{�@e+�ƍ4@>26<�!?�#�ĶK�@�T��O�ٿ}����+�@��q'�4@&�,$��!?�:��+�@&w\Y��ٿ����$�@��9�4@�c�!?s�����@&w\Y��ٿ����$�@��9�4@�c�!?s�����@���Ωٿ���>8�@7"���3@�v�a��!?�c_�F�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@Ӈ"ሮٿ��ZG6�@O�xm+4@5 %��!?��!76�@���<S�ٿޕ[�J�@ܢ ^� 4@�D��!?�Tʇ��@���<S�ٿޕ[�J�@ܢ ^� 4@�D��!?�Tʇ��@���<S�ٿޕ[�J�@ܢ ^� 4@�D��!?�Tʇ��@Y�W��ٿќ>�z��@�����3@R~.�!?��9cnq�@Y�W��ٿќ>�z��@�����3@R~.�!?��9cnq�@Y�W��ٿќ>�z��@�����3@R~.�!?��9cnq�@@.����ٿ������@Y��Yg�3@�����!?�*�`��@@.����ٿ������@Y��Yg�3@�����!?�*�`��@���ٿ���*��@�5 ��4@��S,�!?Q��%�@!ګk�ٿ7_���@�-�f��3@*s�㻏!?ř|ˣ�@!ګk�ٿ7_���@�-�f��3@*s�㻏!?ř|ˣ�@}��`	�ٿ�܍Sk��@��\� 4@	IB��!?p��e�&�@}��`	�ٿ�܍Sk��@��\� 4@	IB��!?p��e�&�@��M[�ٿ��| bq�@Pݜb"�3@�W��ď!?����+�@��M[�ٿ��| bq�@Pݜb"�3@�W��ď!?����+�@�&d��ٿ�3I����@��y"�3@�����!?>�
0�i�@�&d��ٿ�3I����@��y"�3@�����!?>�
0�i�@��ER��ٿ��elf�@;[g��3@�>H��!?��2ǘ��@!��|�ٿ��B�E�@3{O�u 4@%�9[��!?��sa��@!��|�ٿ��B�E�@3{O�u 4@%�9[��!?��sa��@X���ٿ3�8���@`{��=4@�f?���!?iU��;�@L��ឤٿT����h�@�{B4@R��e��!?��o��\�@L��ឤٿT����h�@�{B4@R��e��!?��o��\�@G�ٿ��R�@ڡ�PG 4@�V����!?��y�e�@G�ٿ��R�@ڡ�PG 4@�V����!?��y�e�@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@��@��ٿ���Kjg�@7+-��3@X^뮸�!?k�Q����@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@�{FW�ٿ�\gV�@�~i	~�3@튌��!?���4)��@��u�ٿ�.<y��@�]�Q�3@D��/��!?�e�����@��u�ٿ�.<y��@�]�Q�3@D��/��!?�e�����@��u�ٿ�.<y��@�]�Q�3@D��/��!?�e�����@��u�ٿ�.<y��@�]�Q�3@D��/��!?�e�����@�|�夥ٿ��G74�@����3@[�65��!?X�Ȭ\Y�@�|�夥ٿ��G74�@����3@[�65��!?X�Ȭ\Y�@�|�夥ٿ��G74�@����3@[�65��!?X�Ȭ\Y�@������ٿ�-W��:�@Fs�u�3@��˱Ə!?;�ze;��@������ٿ�-W��:�@Fs�u�3@��˱Ə!?;�ze;��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@���PԚٿ͟�?��@�A�pR4@�{��ˏ!?v�S�E��@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@����ٿ#�i5R��@UY�%�4@t�L���!?=vW���@M�0w��ٿ�X����@�=09��3@�C�R�!?�l�|��@��>���ٿ�;�D��@�i1w 4@MP@7V�!?�}~�l�@��>���ٿ�;�D��@�i1w 4@MP@7V�!?�}~�l�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@�q�գٿ'�`�|��@%^n���3@�5_:��!?^��5k
�@U���]�ٿ����(�@���x�3@]�/�j�!?N��	;I�@U���]�ٿ����(�@���x�3@]�/�j�!?N��	;I�@U���]�ٿ����(�@���x�3@]�/�j�!?N��	;I�@U���]�ٿ����(�@���x�3@]�/�j�!?N��	;I�@��'
�ٿH+P�f�@�᭾ 4@]d!?� Hr��@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@���^�ٿ�dB5��@��ĕ�4@Ðv��!?F��\	8�@my��ܥٿ(�i��@{�gx\ 4@�IF�؏!?.���:��@my��ܥٿ(�i��@{�gx\ 4@�IF�؏!?.���:��@my��ܥٿ(�i��@{�gx\ 4@�IF�؏!?.���:��@my��ܥٿ(�i��@{�gx\ 4@�IF�؏!?.���:��@my��ܥٿ(�i��@{�gx\ 4@�IF�؏!?.���:��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@=8zC͡ٿ�W��N�@s� �
 4@��v;��!?�?�+��@����B�ٿ��>[e�@Z�B��3@>��d��!?�Z�����@����B�ٿ��>[e�@Z�B��3@>��d��!?�Z�����@����B�ٿ��>[e�@Z�B��3@>��d��!?�Z�����@����B�ٿ��>[e�@Z�B��3@>��d��!?�Z�����@����B�ٿ��>[e�@Z�B��3@>��d��!?�Z�����@.t8�ٿa�1E��@$޴� 4@v���!?M�8�6��@I\�7��ٿ����@d�q�4@�~jzӏ!?���'��@I\�7��ٿ����@d�q�4@�~jzӏ!?���'��@����Ϝٿd��V1��@@y9��4@�Q�ǳ�!?�4&�-�@����Ϝٿd��V1��@@y9��4@�Q�ǳ�!?�4&�-�@����Ϝٿd��V1��@@y9��4@�Q�ǳ�!?�4&�-�@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@��?ҫٿ&����@ON8�W 4@q^�1؏!?���5��@�\�"�ٿX��r��@,�@1�4@9�}�!?������@��w8E�ٿc�i��w�@����4@d���n�!?蒈��
�@�k�V�ٿ'��-���@�ޤ�24@��&[��!?Z#��ߺ�@�k�V�ٿ'��-���@�ޤ�24@��&[��!?Z#��ߺ�@�k�V�ٿ'��-���@�ޤ�24@��&[��!?Z#��ߺ�@�k�V�ٿ'��-���@�ޤ�24@��&[��!?Z#��ߺ�@�k�V�ٿ'��-���@�ޤ�24@��&[��!?Z#��ߺ�@�:����ٿ�i~"�	�@�@9�~4@��uw�!?zTH�56�@�:����ٿ�i~"�	�@�@9�~4@��uw�!?zTH�56�@�:����ٿ�i~"�	�@�@9�~4@��uw�!?zTH�56�@����w�ٿ�_�YX��@'wDу�3@�:�l�!?�c,��l�@����w�ٿ�_�YX��@'wDу�3@�:�l�!?�c,��l�@����w�ٿ�_�YX��@'wDу�3@�:�l�!?�c,��l�@����w�ٿ�_�YX��@'wDу�3@�:�l�!?�c,��l�@�e���ٿ:�=X��@y�_ � 4@(ʔ ��!?���ʋ�@%�[舥ٿ�u���@�ؾa��3@�΍��!?�G���@%�[舥ٿ�u���@�ؾa��3@�΍��!?�G���@%�[舥ٿ�u���@�ؾa��3@�΍��!?�G���@%�[舥ٿ�u���@�ؾa��3@�΍��!?�G���@P}`7�ٿ'���@X�4@�1��ڏ!?�l���G�@P}`7�ٿ'���@X�4@�1��ڏ!?�l���G�@P}`7�ٿ'���@X�4@�1��ڏ!?�l���G�@
V)��ٿo�XA��@���XL 4@�����!?�E�~oD�@
V)��ٿo�XA��@���XL 4@�����!?�E�~oD�@
V)��ٿo�XA��@���XL 4@�����!?�E�~oD�@
V)��ٿo�XA��@���XL 4@�����!?�E�~oD�@
V)��ٿo�XA��@���XL 4@�����!?�E�~oD�@.o�$�ٿ1K�Ȏ��@@f��v4@¶�!?��W���@5��k�ٿ���Z���@�<����3@��K�̏!?����^�@Y���ٿ�z�6O��@&3� 4@0�?���!?��7Z-J�@Y���ٿ�z�6O��@&3� 4@0�?���!?��7Z-J�@Y���ٿ�z�6O��@&3� 4@0�?���!?��7Z-J�@Y���ٿ�z�6O��@&3� 4@0�?���!?��7Z-J�@Y���ٿ�z�6O��@&3� 4@0�?���!?��7Z-J�@�[�z]�ٿ��ga�]�@�|z�� 4@�w�Kُ!?���3
�@�[�z]�ٿ��ga�]�@�|z�� 4@�w�Kُ!?���3
�@�[�z]�ٿ��ga�]�@�|z�� 4@�w�Kُ!?���3
�@�/�)�ٿM~<ц��@��O 4@G���ߏ!?��c�~w�@�/�)�ٿM~<ц��@��O 4@G���ߏ!?��c�~w�@�/�)�ٿM~<ц��@��O 4@G���ߏ!?��c�~w�@�/�)�ٿM~<ц��@��O 4@G���ߏ!?��c�~w�@/�a�ٿ��eˍ��@������3@�
%��!?qW)
��@�CQ�2�ٿɁ���@��u�G4@ {�!?�Q��+�@�CQ�2�ٿɁ���@��u�G4@ {�!?�Q��+�@҆z��ٿ��[/Q��@�m��>4@^�bSk�!?��_/%>�@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��M���ٿC�����@��� 4@�%��U�!?}��v[ �@��7��ٿ���aׂ�@2��GS4@"o/�,�!?2R"���@��7��ٿ���aׂ�@2��GS4@"o/�,�!?2R"���@��7��ٿ���aׂ�@2��GS4@"o/�,�!?2R"���@-[�!�ٿ�3g*��@Z��C4@'c��!?�"]Ϸ��@-[�!�ٿ�3g*��@Z��C4@'c��!?�"]Ϸ��@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@�ʗٿ��e+�?�@[��0� 4@"�!���!?���nϼ�@ղ{)�ٿ���1"�@a@�: 4@���AM�!?������@�e��֜ٿ1�}�Q3�@DHȁ�3@T_F]��!?u�����@��	�ٿ��j�/�@9��) 4@>�`�ߏ!?�Wwf߄�@��	�ٿ��j�/�@9��) 4@>�`�ߏ!?�Wwf߄�@��	�ٿ��j�/�@9��) 4@>�`�ߏ!?�Wwf߄�@��	�ٿ��j�/�@9��) 4@>�`�ߏ!?�Wwf߄�@T�?�ǣٿ,6�Sd��@V��A4@|[���!?d���f��@T�?�ǣٿ,6�Sd��@V��A4@|[���!?d���f��@T�?�ǣٿ,6�Sd��@V��A4@|[���!?d���f��@T�?�ǣٿ,6�Sd��@V��A4@|[���!?d���f��@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@å�ٿ���2��@�����3@�,����!?�}"���@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@e%�-�ٿMր*��@V�Q��3@�'O�ɏ!?�h����@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�)�懣ٿ�����@mD��: 4@_�߯��!?���e	6�@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@�ڛR�ٿz������@���r 4@5�{���!?N� ����@��Bu�ٿ+�h���@]�6Qw4@}yYȻ�!?���`
�@��Bu�ٿ+�h���@]�6Qw4@}yYȻ�!?���`
�@�z�.&�ٿ��\�@8=_ 4@[P��Ώ!?��VT�U�@�z�.&�ٿ��\�@8=_ 4@[P��Ώ!?��VT�U�@�z�.&�ٿ��\�@8=_ 4@[P��Ώ!?��VT�U�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@�>f��ٿ��)��@j'= � 4@�S��!?0¿��e�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@1u���ٿQ��:���@�~rG&4@��h��!?�B�{�@�Z80��ٿ�6=3���@7�:�� 4@��%[��!?%�p7+�@�Z80��ٿ�6=3���@7�:�� 4@��%[��!?%�p7+�@�z*Ơ�ٿK���@�㣚 4@+k�ۏ!?W���@�z*Ơ�ٿK���@�㣚 4@+k�ۏ!?W���@+(�ٿI�F��@%�{Y 4@t��fk�!?����8��@GM�28�ٿ5؆��@�\ng��3@p�͵�!?t/���=�@��e��ٿ��hҸ\�@���r��3@�ԥ�!?�4�]/�@��e��ٿ��hҸ\�@���r��3@�ԥ�!?�4�]/�@��bȯٿ\	Z���@ݕ���3@�uR�Ə!?�8����@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�n���ٿ-͒	���@-Ϊ$54@w�g%�!?+��A�s�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@�F��ٿ��g�z�@�{"� 4@��٥��!?�q�	�r�@~���g�ٿ�_ v�@�,�W� 4@�a��ߏ!?D�d�$_�@��|q�ٿ6�>q��@��٠�4@�*�w�!?C�M;��@��|q�ٿ6�>q��@��٠�4@�*�w�!?C�M;��@e+�cQ�ٿ�����@+�)f 4@����}�!?�)��4��@e+�cQ�ٿ�����@+�)f 4@����}�!?�)��4��@e+�cQ�ٿ�����@+�)f 4@����}�!?�)��4��@�-�"�ٿ��sR���@�����3@�^�Hy�!?ɖm,��@m�K �ٿ{���,��@}�f���3@�u��"�!?`B���@m�K �ٿ{���,��@}�f���3@�u��"�!?`B���@Z��Ҥٿ!���#S�@3�~���3@��x�*�!?21!�^��@Z��Ҥٿ!���#S�@3�~���3@��x�*�!?21!�^��@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@D�ig�ٿ�n}	'�@#wiq��3@q�!���!?��G���@�t��L�ٿ��|��@C��ſ�3@ �Z�!?R$6ͣ��@�t��L�ٿ��|��@C��ſ�3@ �Z�!?R$6ͣ��@�t��L�ٿ��|��@C��ſ�3@ �Z�!?R$6ͣ��@�t��L�ٿ��|��@C��ſ�3@ �Z�!?R$6ͣ��@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@lQ3�ۮٿ(6�(���@��; 4@��]��!?R��4!s�@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�8���ٿ�]]J)r�@
�ɋ�3@KS\}��!?kQ����@�d�V��ٿ&A܀2��@�b i��3@xB����!?G��	���@�1��;�ٿB�����@b�?E��3@�}݁ɏ!?�Xmn�&�@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@jSO�I�ٿ|�(���@]�Q 4@�L�.��!?��R���@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@ ��b�ٿj:B}*M�@�٘� 4@�%/��!?���f!I�@?t�Ħٿ��_{?�@?�� 4@*"����!?���9�@?t�Ħٿ��_{?�@?�� 4@*"����!?���9�@?t�Ħٿ��_{?�@?�� 4@*"����!?���9�@?t�Ħٿ��_{?�@?�� 4@*"����!?���9�@S_~��ٿ����8Z�@��:� 4@u�n��!?Qb���@S_~��ٿ����8Z�@��:� 4@u�n��!?Qb���@S_~��ٿ����8Z�@��:� 4@u�n��!?Qb���@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@V��,�ٿ�r׈�M�@��%�
4@���°�!?��D� �@��+!�ٿ�����@!<���3@@�}�!�!?o����@��+!�ٿ�����@!<���3@@�}�!�!?o����@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@��j��ٿ�,�<�@"�����3@�wȈ��!?R�])���@Ue9�ٿ�v}����@���74@RI�y��!?F �k���@Ue9�ٿ�v}����@���74@RI�y��!?F �k���@Ue9�ٿ�v}����@���74@RI�y��!?F �k���@Ue9�ٿ�v}����@���74@RI�y��!?F �k���@�#��Ʊٿ�jw�{&�@�󍹾4@�P�]̏!?��pqr�@�r��Էٿ\��˥�@��y�4@��9��!?�\�	19�@w��+Σٿ�.�
��@QJ��4@#��P��!?�nC�L��@ѫ��جٿv�d�R�@/�z�C4@�ǉ~�!?�8$���@ѫ��جٿv�d�R�@/�z�C4@�ǉ~�!?�8$���@x)�� �ٿ0��g��@�
Ϙ 4@g:�Q�!?�x^3���@금�#�ٿ���5���@l���3@���U�!?�� *n�@금�#�ٿ���5���@l���3@���U�!?�� *n�@n5�şٿ�|}r�@�(�4@rB�AU�!?z��d���@n5�şٿ�|}r�@�(�4@rB�AU�!?z��d���@n5�şٿ�|}r�@�(�4@rB�AU�!?z��d���@n5�şٿ�|}r�@�(�4@rB�AU�!?z��d���@n5�şٿ�|}r�@�(�4@rB�AU�!?z��d���@�{�˯�ٿ[--���@#�P�n4@ �;��!?b��ҥ(�@�{�˯�ٿ[--���@#�P�n4@ �;��!?b��ҥ(�@c���ٿÔb���@W�#��4@?g�*��!?էT���@c���ٿÔb���@W�#��4@?g�*��!?էT���@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@�I�\��ٿ�LT�r�@K�G�f4@7�Ц�!?�v߄�9�@~�jE�ٿ6�.�̯�@��2�4@1Wz{5�!?��y���@~�jE�ٿ6�.�̯�@��2�4@1Wz{5�!?��y���@~�jE�ٿ6�.�̯�@��2�4@1Wz{5�!?��y���@~�jE�ٿ6�.�̯�@��2�4@1Wz{5�!?��y���@��>�ٿ�5��>Y�@�k�@4@eT[�!?�����Z�@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@��t���ٿ���c�t�@/9�, 4@��U���!?�zQ�	��@4L'��ٿc��Lo�@w�]k� 4@��I��!?i��+���@]^Q.�ٿ���Q�@uGY1� 4@��K��!?��EL��@�B�B��ٿ����O�@��*/��3@�$Û��!?V�٫%�@�B�B��ٿ����O�@��*/��3@�$Û��!?V�٫%�@ÝY��ٿ'�B����@jvd9&4@��a��!?vZ���@��w⧤ٿ��G��@�K��T 4@�C����!?�V�i<�@��w⧤ٿ��G��@�K��T 4@�C����!?�V�i<�@��w⧤ٿ��G��@�K��T 4@�C����!?�V�i<�@��w⧤ٿ��G��@�K��T 4@�C����!?�V�i<�@��w⧤ٿ��G��@�K��T 4@�C����!?�V�i<�@Qb�ٿ;���x��@���;�4@�Zr�!?�?C����@Qb�ٿ;���x��@���;�4@�Zr�!?�?C����@Qb�ٿ;���x��@���;�4@�Zr�!?�?C����@Qb�ٿ;���x��@���;�4@�Zr�!?�?C����@�P�փ�ٿ��L��@O%�M� 4@�[E[`�!?�?*�5�@�P�փ�ٿ��L��@O%�M� 4@�[E[`�!?�?*�5�@�P�փ�ٿ��L��@O%�M� 4@�[E[`�!?�?*�5�@�[��ٿ_�Kՠ�@c\W���3@88ן/�!?�{��n��@�[��ٿ_�Kՠ�@c\W���3@88ן/�!?�{��n��@�[��ٿ_�Kՠ�@c\W���3@88ן/�!?�{��n��@�[��ٿ_�Kՠ�@c\W���3@88ן/�!?�{��n��@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@�
Xq�ٿr��Ֆs�@]I�X�3@٧õ��!?L3����@����̘ٿ:�J���@�Z*;4@xcy&ʏ!?��"��@����̘ٿ:�J���@�Z*;4@xcy&ʏ!?��"��@����̘ٿ:�J���@�Z*;4@xcy&ʏ!?��"��@����̘ٿ:�J���@�Z*;4@xcy&ʏ!?��"��@3����ٿ�w�ܲ��@pI��4@KC�4֏!?�{鱗y�@3����ٿ�w�ܲ��@pI��4@KC�4֏!?�{鱗y�@3����ٿ�w�ܲ��@pI��4@KC�4֏!?�{鱗y�@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@�5���ٿ���LT�@Lq��4@���u�!?����@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@m�,�ٿo����@�Rp�m4@ت�_ŏ!?�}%��@]�*2��ٿ������@�$!b4@�����!?�KV(wm�@]�*2��ٿ������@�$!b4@�����!?�KV(wm�@F�C��ٿD�=?��@(Y'4@\"�C��!?`=��_�@F�C��ٿD�=?��@(Y'4@\"�C��!?`=��_�@F�C��ٿD�=?��@(Y'4@\"�C��!?`=��_�@F�C��ٿD�=?��@(Y'4@\"�C��!?`=��_�@F�C��ٿD�=?��@(Y'4@\"�C��!?`=��_�@�!���ٿҢU�P��@�ו�c4@��U�!?��v�=�@�!���ٿҢU�P��@�ו�c4@��U�!?��v�=�@�!���ٿҢU�P��@�ו�c4@��U�!?��v�=�@�!���ٿҢU�P��@�ו�c4@��U�!?��v�=�@�!���ٿҢU�P��@�ו�c4@��U�!?��v�=�@�ږ�ٿ	F��@q��^ 4@K���L�!?~��'�@�ږ�ٿ	F��@q��^ 4@K���L�!?~��'�@�ږ�ٿ	F��@q��^ 4@K���L�!?~��'�@�ږ�ٿ	F��@q��^ 4@K���L�!?~��'�@�ږ�ٿ	F��@q��^ 4@K���L�!?~��'�@����ٿ�G�Kz��@��M�4@�3�/��!?�D��f��@Z�/�ٿ��y�� �@ ��� 4@���!?ށP��D�@Z�/�ٿ��y�� �@ ��� 4@���!?ށP��D�@Z�/�ٿ��y�� �@ ��� 4@���!?ށP��D�@Z�/�ٿ��y�� �@ ��� 4@���!?ށP��D�@Z�/�ٿ��y�� �@ ��� 4@���!?ށP��D�@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@?e�-�ٿ�g���@��w�; 4@(�@�!?��{���@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@��$�ٿ�֑�A�@8��r� 4@�S�]؏!?߰~�u�@���L�ٿo��v8�@�F�� 4@�}��!?�6"�@�}�wN�ٿ�M��j�@{w�S4@ܒ�:/�!?�l��u�@�}�wN�ٿ�M��j�@{w�S4@ܒ�:/�!?�l��u�@��Z��ٿ�f! �(�@��/uK4@$'�P�!?��M���@��Z��ٿ�f! �(�@��/uK4@$'�P�!?��M���@��Z��ٿ�f! �(�@��/uK4@$'�P�!?��M���@��i��ٿ�nĘ���@��uBl4@�����!?^	����@��i��ٿ�nĘ���@��uBl4@�����!?^	����@��i��ٿ�nĘ���@��uBl4@�����!?^	����@��i��ٿ�nĘ���@��uBl4@�����!?^	����@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@ �o�ٿ�G0Հ��@�"�@4@Y�Q�h�!?��	���@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@r��^�ٿ �[u�(�@�)֗4@�׬f��!?-�����@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@�+);�ٿ�]S,v�@o�� 4@�V�m��!?�w��@y<L��ٿ���e��@�Y�G� 4@7�|��!?W�Ua��@y<L��ٿ���e��@�Y�G� 4@7�|��!?W�Ua��@y<L��ٿ���e��@�Y�G� 4@7�|��!?W�Ua��@y<L��ٿ���e��@�Y�G� 4@7�|��!?W�Ua��@8(&�ٿ�s�6]�@����3@�>nO�!?�:/����@8(&�ٿ�s�6]�@����3@�>nO�!?�:/����@8(&�ٿ�s�6]�@����3@�>nO�!?�:/����@8(&�ٿ�s�6]�@����3@�>nO�!?�:/����@��E��ٿ��M��F�@��$�f4@�'�|�!?����&�@��E��ٿ��M��F�@��$�f4@�'�|�!?����&�@��E��ٿ��M��F�@��$�f4@�'�|�!?����&�@��E��ٿ��M��F�@��$�f4@�'�|�!?����&�@��E��ٿ��M��F�@��$�f4@�'�|�!?����&�@�߷�R�ٿ4�r���@d�74@Q���!?�*��.�@d< B8�ٿnվ����@$�b>4@�L���!?�eC`��@d< B8�ٿnվ����@$�b>4@�L���!?�eC`��@�U?Wҫٿ��CۉZ�@��7�?4@9Tt�!?]�J���@�U?Wҫٿ��CۉZ�@��7�?4@9Tt�!?]�J���@�U?Wҫٿ��CۉZ�@��7�?4@9Tt�!?]�J���@�U?Wҫٿ��CۉZ�@��7�?4@9Tt�!?]�J���@2ÂLy�ٿu;xna�@lBԢ$4@)��"�!?�S��Bx�@2ÂLy�ٿu;xna�@lBԢ$4@)��"�!?�S��Bx�@�s�;�ٿx���7�@$�`��4@�1�x�!?��R2F��@�s�;�ٿx���7�@$�`��4@�1�x�!?��R2F��@�s�;�ٿx���7�@$�`��4@�1�x�!?��R2F��@�s�;�ٿx���7�@$�`��4@�1�x�!?��R2F��@�z�u�ٿ�Z/���@��I~4@*HY�!?τb����@�z�u�ٿ�Z/���@��I~4@*HY�!?τb����@�z�u�ٿ�Z/���@��I~4@*HY�!?τb����@��Z�ٛٿ��3 ��@Ba��[ 4@�Mn��!?��.j���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@���F��ٿ��L���@���4@�_�*Y�!?�Դ5���@npA^Y�ٿ��ֱ���@�n�4��3@�d;�@�!?�+����@npA^Y�ٿ��ֱ���@�n�4��3@�d;�@�!?�+����@npA^Y�ٿ��ֱ���@�n�4��3@�d;�@�!?�+����@npA^Y�ٿ��ֱ���@�n�4��3@�d;�@�!?�+����@}r=*K�ٿ7��#�@�Xt�E�3@��D*��!?s�d���@}r=*K�ٿ7��#�@�Xt�E�3@��D*��!?s�d���@Fjq.�ٿ�8ww��@�&� 4@$���Ə!?�UД��@Fjq.�ٿ�8ww��@�&� 4@$���Ə!?�UД��@Fjq.�ٿ�8ww��@�&� 4@$���Ə!?�UД��@M/e��ٿ��|��1�@\��4@�p��!?:���@M/e��ٿ��|��1�@\��4@�p��!?:���@��Zb�ٿ���+"z�@����4@=��ݲ�!?*6�R��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@���I�ٿh��+���@����4@Y�-\Ï!?�g��@d����ٿ�?b��@�W�� 4@_<�͏!?�A�:X?�@d����ٿ�?b��@�W�� 4@_<�͏!?�A�:X?�@���eO�ٿ95K����@��L4@jkbf!?�^�s�@-i:��ٿ+�����@߂�Z 4@�q�<��!?�$���@-i:��ٿ+�����@߂�Z 4@�q�<��!?�$���@-i:��ٿ+�����@߂�Z 4@�q�<��!?�$���@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@H>�D�ٿ38�
ٹ�@�#u*a4@G��6��!?��lb%��@]�ځ�ٿD�f�a��@�ٖ�4@�lŢ�!?�)�(�U�@K����ٿ���34��@w�u�4@� ���!?�hk�q�@ua8��ٿ�_�E��@� ��-4@	ϫg��!?�Eif�J�@ua8��ٿ�_�E��@� ��-4@	ϫg��!?�Eif�J�@ua8��ٿ�_�E��@� ��-4@	ϫg��!?�Eif�J�@ua8��ٿ�_�E��@� ��-4@	ϫg��!?�Eif�J�@�캟ٿ0i�a���@V�� 4@�L�u��!?�Q��,�@�캟ٿ0i�a���@V�� 4@�L�u��!?�Q��,�@�Uw�ٿMG|���@LRB�	4@w�"�֏!?Q����@�{�`ԫٿ:*�b���@��'֊4@�z�G��!?��� y��@�{�`ԫٿ:*�b���@��'֊4@�z�G��!?��� y��@�{�`ԫٿ:*�b���@��'֊4@�z�G��!?��� y��@��z;r�ٿ�Lw���@l��4@��ଏ!?���J��@�%�ɞٿ���-�@2q�� 4@܎�'��!?	,���`�@�%�ɞٿ���-�@2q�� 4@܎�'��!?	,���`�@�%�ɞٿ���-�@2q�� 4@܎�'��!?	,���`�@�%�ɞٿ���-�@2q�� 4@܎�'��!?	,���`�@��	�P�ٿ$ay���@�8� 4@��&:�!?�����@��	�P�ٿ$ay���@�8� 4@��&:�!?�����@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@�%�)�ٿ^��_���@)��V��3@P2 P�!?�^h�9��@o�����ٿ��L��G�@v����4@�$*h�!?������@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@yW��5�ٿ�����@�J��4@1��U�!?�z��N��@��hp��ٿ�qW;��@Z��o��3@�_+R��!?jz�˲��@�j+��ٿ]��ڲW�@ RO��3@�!ԏ!?��f����@�j+��ٿ]��ڲW�@ RO��3@�!ԏ!?��f����@�j+��ٿ]��ڲW�@ RO��3@�!ԏ!?��f����@�j+��ٿ]��ڲW�@ RO��3@�!ԏ!?��f����@�j+��ٿ]��ڲW�@ RO��3@�!ԏ!?��f����@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@^N-ƥ�ٿ���D��@��)��3@�d�4��!?_*i ���@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@�0y�ƞٿ�+I�f��@����� 4@�<����!? ��?��@8:�)��ٿ���.φ�@����3@�;^9��!?[q�-�@8:�)��ٿ���.φ�@����3@�;^9��!?[q�-�@8:�)��ٿ���.φ�@����3@�;^9��!?[q�-�@8:�)��ٿ���.φ�@����3@�;^9��!?[q�-�@�-�c�ٿ����<��@��1��3@�Y����!?�~;���@�-�c�ٿ����<��@��1��3@�Y����!?�~;���@�-�c�ٿ����<��@��1��3@�Y����!?�~;���@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@�!�2|�ٿ��	q�7�@|�z�4@8�u��!?$;�V ��@C�����ٿ�
����@�TP�4@��3�͏!?U~��p�@C�����ٿ�
����@�TP�4@��3�͏!?U~��p�@C�����ٿ�
����@�TP�4@��3�͏!?U~��p�@�=o�b�ٿ;�`//$�@i�^4@vss�z�!?E��M-"�@�=o�b�ٿ;�`//$�@i�^4@vss�z�!?E��M-"�@���U|�ٿ�J�t��@�k��4@�$���!?Q�)-j��@���U|�ٿ�J�t��@�k��4@�$���!?Q�)-j��@^�X<��ٿ�Pi�n��@��ą
4@�)Y�}�!?�q�\'��@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@" ��ٿ�t� J��@?�f |4@r����!?�F,�7�@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@k���ٿX��~S��@��-�h4@�f�C�!?f0��f��@��y(J�ٿ>N��5��@�_���3@A(�ek�!?�7ߋ��@�}��8�ٿ��p�@S���3@��m�~�!?�r����@A	�-�ٿF�ѧ���@^_\��4@����!?���c��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@V���L�ٿ����@K\�c4@�����!?�᥽]��@��i�ٿ�GS,v�@�8����3@fzC�!?����:��@��i�ٿ�GS,v�@�8����3@fzC�!?����:��@��i�ٿ�GS,v�@�8����3@fzC�!?����:��@c�
u�ٿl�yM�W�@}�Z��3@\����!?�	����@c�
u�ٿl�yM�W�@}�Z��3@\����!?�	����@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@+����ٿ_�8\;�@���I�3@;���!?3��P��@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@S���ٿy��ʐ$�@����3@B��!?�>���P�@�g��Ұٿvwbи��@,ř��3@��_?��!?p�X<J��@�g��Ұٿvwbи��@,ř��3@��_?��!?p�X<J��@�g��Ұٿvwbи��@,ř��3@��_?��!?p�X<J��@�g��Ұٿvwbи��@,ř��3@��_?��!?p�X<J��@�c�i�ٿ+dm���@�K^���3@�H�N��!?j��2B��@9�W�ƫٿ�4�[L��@��1�=�3@@󲄖�!?�?�ޛ-�@9�W�ƫٿ�4�[L��@��1�=�3@@󲄖�!?�?�ޛ-�@9�W�ƫٿ�4�[L��@��1�=�3@@󲄖�!?�?�ޛ-�@��o|-�ٿiAo+�@*�xٿ�3@5�'���!?������@��o|-�ٿiAo+�@*�xٿ�3@5�'���!?������@��o|-�ٿiAo+�@*�xٿ�3@5�'���!?������@��o|-�ٿiAo+�@*�xٿ�3@5�'���!?������@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@��4��ٿYT �A5�@�P�p 4@mS�囏!?Cф2���@Yܧ�ٿ�+g&��@Y�*�4@�jInz�!?���T��@Yܧ�ٿ�+g&��@Y�*�4@�jInz�!?���T��@Yܧ�ٿ�+g&��@Y�*�4@�jInz�!?���T��@Yܧ�ٿ�+g&��@Y�*�4@�jInz�!?���T��@Yܧ�ٿ�+g&��@Y�*�4@�jInz�!?���T��@t�?��ٿ~T��E��@@��� 4@��!?J���1�@t�?��ٿ~T��E��@@��� 4@��!?J���1�@t�?��ٿ~T��E��@@��� 4@��!?J���1�@t�?��ٿ~T��E��@@��� 4@��!?J���1�@A�ݝٿ��%�@@�&�v�3@������!?'GN:�T�@�I�V�ٿ��֬��@_ܩ�� 4@-��ň�!?�ٜ�
k�@/���s�ٿ'R�"K��@AAi�4@��2�!?ȃ���K�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@>�r�ٿ;Y[��r�@4lW��4@9�[X�!?:V�he'�@�6��ٿ��B�S��@Y��i4@��n�!?CS�f0��@�Y�4ҟٿ����WA�@�k�)�4@d�>ȏ!?v�C���@�Y�4ҟٿ����WA�@�k�)�4@d�>ȏ!?v�C���@�Y�4ҟٿ����WA�@�k�)�4@d�>ȏ!?v�C���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@kn-�P�ٿ�&N#c��@@%+4@(0f&��!?���$���@�;��O�ٿ�J�E��@�(��� 4@�9��Ώ!?N����@�;��O�ٿ�J�E��@�(��� 4@�9��Ώ!?N����@�;��O�ٿ�J�E��@�(��� 4@�9��Ώ!?N����@�;��O�ٿ�J�E��@�(��� 4@�9��Ώ!?N����@�;��O�ٿ�J�E��@�(��� 4@�9��Ώ!?N����@'����ٿSQ���@����� 4@l�A��!?�o�]�k�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@u'ϯٿ��8j���@�J���3@X��^ԏ!?�YF�
�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@`�PVg�ٿ�M��'�@�MX�~ 4@����!?��cb�Q�@�PP+�ٿ>>qg�Q�@�^� 4@o���!?����/�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@�D��8�ٿ	/:���@��!'� 4@����!?v9���G�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@ ��Üٿ"�Z�!��@!�g��3@�)k��!?|2��h�@��E��ٿ�.��#i�@�Z���3@�xŖo�!?Ǐ��@��E��ٿ�.��#i�@�Z���3@�xŖo�!?Ǐ��@�(P�h�ٿ�u\e
��@h��4�4@N�����!?�ʌ����@�(P�h�ٿ�u\e
��@h��4�4@N�����!?�ʌ����@�(P�h�ٿ�u\e
��@h��4�4@N�����!?�ʌ����@�(P�h�ٿ�u\e
��@h��4�4@N�����!?�ʌ����@A����ٿ�c���@������3@bP���!?�\����@A����ٿ�c���@������3@bP���!?�\����@A����ٿ�c���@������3@bP���!?�\����@A����ٿ�c���@������3@bP���!?�\����@A����ٿ�c���@������3@bP���!?�\����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@@5��/�ٿ�a0}Q��@�	"2��3@���я!?j����@^(��ٿ���:�t�@��-�(�3@,�@��!?���*��@^(��ٿ���:�t�@��-�(�3@,�@��!?���*��@��1��ٿ��u�v�@t$�� �3@ਥ��!?ŉɏ��@�j�Y0�ٿU ��
��@�� �� 4@mb&�!?"W����@�j�Y0�ٿU ��
��@�� �� 4@mb&�!?"W����@�j�Y0�ٿU ��
��@�� �� 4@mb&�!?"W����@ \��s�ٿXʧ�u�@�MYb�3@>�i�؏!?!k�m&��@���ٯٿ�_��w��@�Q����3@�]�B��!?sMwng�@$�d��ٿ�����E�@f5��q 4@1�l!?�u� T�@$�d��ٿ�����E�@f5��q 4@1�l!?�u� T�@$�d��ٿ�����E�@f5��q 4@1�l!?�u� T�@���\h�ٿ+2*4��@k1�`� 4@��,�U�!? �ڹ�@���\h�ٿ+2*4��@k1�`� 4@��,�U�!? �ڹ�@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@y�c�ٿ�����@���$ 4@j�nW��!?�F�	 ��@h֩�ٿ��ӗ���@�A=��4@BM�f��!?��"K���@h֩�ٿ��ӗ���@�A=��4@BM�f��!?��"K���@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@��@ؙٿ<�{��=�@TV�B)4@#��{��!?������@�]�_��ٿ�<Ȃ�@.D����3@n�Qr��!?��<��@�]�_��ٿ�<Ȃ�@.D����3@n�Qr��!?��<��@�]�_��ٿ�<Ȃ�@.D����3@n�Qr��!?��<��@�]�_��ٿ�<Ȃ�@.D����3@n�Qr��!?��<��@PB�m��ٿV�D��l�@��K�4@q��:��!?,m����@PB�m��ٿV�D��l�@��K�4@q��:��!?,m����@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@�Sݼ�ٿ	�+�y�@�/lS#4@���=�!?7���>�@����6�ٿ�u ��#�@�vɷ� 4@*��;�!?Y�-��L�@����6�ٿ�u ��#�@�vɷ� 4@*��;�!?Y�-��L�@����6�ٿ�u ��#�@�vɷ� 4@*��;�!?Y�-��L�@�(#Ur�ٿ��A���@�����3@��W��!?��<�@�(#Ur�ٿ��A���@�����3@��W��!?��<�@�(#Ur�ٿ��A���@�����3@��W��!?��<�@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@�0�fL�ٿ:�9�O�@y���4@P�ݤ�!?=ETN���@L���ٿ$�Bsm^�@N���"4@��}Kf�!?��7����@L���ٿ$�Bsm^�@N���"4@��}Kf�!?��7����@
��r�ٿJ,kH�n�@K�&�4@@#"Y�!?(��X�@^p|B�ٿ�m�.���@��_��3@Ϯ:�n�!?e2Hc�@^p|B�ٿ�m�.���@��_��3@Ϯ:�n�!?e2Hc�@^p|B�ٿ�m�.���@��_��3@Ϯ:�n�!?e2Hc�@��λc�ٿ�v��s �@9�A�3@�OV�e�!?�����I�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@��O��ٿ~�=K��@�*Pp��3@M0���!?��2ҕr�@���ٿ���t�~�@�괎 4@��Oل�!?�t��.�@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@�]vb �ٿ�Ce��S�@-HM^��3@��u���!?�9����@/�c.�ٿ��>?y�@��ΠH4@�˘ᙏ!?��,!��@/�c.�ٿ��>?y�@��ΠH4@�˘ᙏ!?��,!��@/�c.�ٿ��>?y�@��ΠH4@�˘ᙏ!?��,!��@/�c.�ٿ��>?y�@��ΠH4@�˘ᙏ!?��,!��@/�c.�ٿ��>?y�@��ΠH4@�˘ᙏ!?��,!��@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@����e�ٿ3�,^���@����,4@)I,���!?�>!@	,�@�&����ٿ��tT���@�J, 4@g�U��!?2$6�y�@�&����ٿ��tT���@�J, 4@g�U��!?2$6�y�@�&����ٿ��tT���@�J, 4@g�U��!?2$6�y�@�&����ٿ��tT���@�J, 4@g�U��!?2$6�y�@����ٿD���i��@^�1�� 4@��)��!?�����@����ٿD���i��@^�1�� 4@��)��!?�����@M<�F��ٿ��A���@�"դ�3@ N�b�!?�����@'��$#�ٿ�㼵���@d�*���3@�G��S�!?~�$
!�@'��$#�ٿ�㼵���@d�*���3@�G��S�!?~�$
!�@�MC�ٿ�9�V[�@̭�94@���z�!?F�gJ�@�MC�ٿ�9�V[�@̭�94@���z�!?F�gJ�@ %Sd��ٿ��i[���@<��d@ 4@���e�!?��A�C�@ %Sd��ٿ��i[���@<��d@ 4@���e�!?��A�C�@ %Sd��ٿ��i[���@<��d@ 4@���e�!?��A�C�@ %Sd��ٿ��i[���@<��d@ 4@���e�!?��A�C�@ %Sd��ٿ��i[���@<��d@ 4@���e�!?��A�C�@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@*p@MD�ٿ<��VG��@�ͭ�� 4@��B��!?�b���@gzv�ٿ��5i��@u���3@0�Wg�!?��b�r�@gzv�ٿ��5i��@u���3@0�Wg�!?��b�r�@gzv�ٿ��5i��@u���3@0�Wg�!?��b�r�@gzv�ٿ��5i��@u���3@0�Wg�!?��b�r�@���x��ٿm`����@������3@H���S�!?��D�A�@ﱇM#�ٿ�hS�@���r�3@�&��!?�� ܵ�@ﱇM#�ٿ�hS�@���r�3@�&��!?�� ܵ�@ﱇM#�ٿ�hS�@���r�3@�&��!?�� ܵ�@QNe�^�ٿ�j3T���@������3@���,��!?��f�6r�@r�����ٿg��,I�@�n�y� 4@N�Hя!?ͨf��@r�����ٿg��,I�@�n�y� 4@N�Hя!?ͨf��@3M�;צٿ��D�]$�@�xv�� 4@ETJ���!?�#܍8��@3M�;צٿ��D�]$�@�xv�� 4@ETJ���!?�#܍8��@3M�;צٿ��D�]$�@�xv�� 4@ETJ���!?�#܍8��@�`�Gx�ٿ���>܆�@ث��q4@e��y�!?�R8]h�@�`�Gx�ٿ���>܆�@ث��q4@e��y�!?�R8]h�@�`�Gx�ٿ���>܆�@ث��q4@e��y�!?�R8]h�@�`�Gx�ٿ���>܆�@ث��q4@e��y�!?�R8]h�@�`�Gx�ٿ���>܆�@ث��q4@e��y�!?�R8]h�@�~ĩ�ٿ�9�7�@�!h��4@_I���!?�aT0;�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��/�ٿ*f�A<��@�@���3@�D�m�!?�OC�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@��+�ȣٿc;���@��W��3@%_hk�!?_�#��!�@�bl�ǧٿ�9����@�{��1 4@*���]�!?1���@�bl�ǧٿ�9����@�{��1 4@*���]�!?1���@�bl�ǧٿ�9����@�{��1 4@*���]�!?1���@��U��ٿk��;���@W�{�4@bQ콏!?��T6Vn�@��U��ٿk��;���@W�{�4@bQ콏!?��T6Vn�@�bb��ٿ/d' 	��@r��4@��f;��!?~�f�F��@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@f5GWD�ٿ��_]3��@��eΓ 4@^����!?zA�z���@L�#���ٿb{�`��@ϗ�$o4@���!?�����@L�#���ٿb{�`��@ϗ�$o4@���!?�����@L�#���ٿb{�`��@ϗ�$o4@���!?�����@L�#���ٿb{�`��@ϗ�$o4@���!?�����@L�#���ٿb{�`��@ϗ�$o4@���!?�����@O�z��ٿ�Y�ZA�@`�狣4@[��6ߏ!?�K��uH�@������ٿ1 �'+:�@��4@ũ+Џ!?r���@������ٿ1 �'+:�@��4@ũ+Џ!?r���@������ٿ1 �'+:�@��4@ũ+Џ!?r���@������ٿ1 �'+:�@��4@ũ+Џ!?r���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@¶��+�ٿ�=l�d�@���z4@��}9��!?�n;i���@��� �ٿS$U���@𜴜� 4@,jps�!?�3>n`f�@��L�W�ٿ��3���@.KT� 4@OT�As�!?Z�ŋz�@��L�W�ٿ��3���@.KT� 4@OT�As�!?Z�ŋz�@nGL���ٿ���u��@Z?�� 4@����y�!?|E�b��@nGL���ٿ���u��@Z?�� 4@����y�!?|E�b��@nGL���ٿ���u��@Z?�� 4@����y�!?|E�b��@nGL���ٿ���u��@Z?�� 4@����y�!?|E�b��@����s�ٿ�ΘW��@S� `4@����Z�!?L�D-
�@��fj�ٿ���j��@��e|4@1��U�!?Sa~����@��fj�ٿ���j��@��e|4@1��U�!?Sa~����@��fj�ٿ���j��@��e|4@1��U�!?Sa~����@Tg�ٿ�>�l�t�@'4���3@u���ُ!?K��x+�@Tg�ٿ�>�l�t�@'4���3@u���ُ!?K��x+�@Tg�ٿ�>�l�t�@'4���3@u���ُ!?K��x+�@v�e�ٿ�޻��@��v|�3@���U_�!?�7��7g�@j�_��ٿ{܊\�o�@J��-a 4@�S��:�!?� q:�~�@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@4�r�ٿ��I|��@Ɂ$�)4@}��bw�!?�W�b���@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@��3[�ٿ���� �@�<�'n 4@��7��!?PZ�
�@�?�Ԉ�ٿ���Fp5�@�ĕ{4@7�7��!?�l�H�@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@Q�y_�ٿ�����@]����3@����!?W6��T��@��F���ٿ^ἃI��@} $ҳ�3@��@ܕ�!?�h��@��F���ٿ^ἃI��@} $ҳ�3@��@ܕ�!?�h��@�y�ޞٿ$���$��@�H#1?4@̌�f��!?�ώ�Ǹ�@�RЎ�ٿ���B�@k���> 4@�����!?j�1�m��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@Z��q�ٿ��B��@�ӆ ��3@�g�9��!?F��h"��@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@����ٿ�N�[��@�*�T 4@LM��ŏ!?���u�@>�땈�ٿ�z�E�@%o
��3@�y����!?}�O�O��@>�땈�ٿ�z�E�@%o
��3@�y����!?}�O�O��@��r��ٿ��?Z�m�@>)�4@Lo��!?B����@��r��ٿ��?Z�m�@>)�4@Lo��!?B����@�;
��ٿ0"+��p�@��Ә}4@����!?���r��@�;
��ٿ0"+��p�@��Ә}4@����!?���r��@�;
��ٿ0"+��p�@��Ә}4@����!?���r��@�;
��ٿ0"+��p�@��Ә}4@����!?���r��@�;
��ٿ0"+��p�@��Ә}4@����!?���r��@�"�e��ٿ	�~��@(Ԭ��4@܍ˏ!?&�d���@�"�e��ٿ	�~��@(Ԭ��4@܍ˏ!?&�d���@hS5��ٿ��e��@����Z4@3��!?�����@hS5��ٿ��e��@����Z4@3��!?�����@hS5��ٿ��e��@����Z4@3��!?�����@"���f�ٿG�D����@��i\4@�9SeЏ!?�b���@"���f�ٿG�D����@��i\4@�9SeЏ!?�b���@����ٿpRI���@��%� 4@<v���!?v�=C�@����ٿpRI���@��%� 4@<v���!?v�=C�@����ٿpRI���@��%� 4@<v���!?v�=C�@����ٿpRI���@��%� 4@<v���!?v�=C�@����ٿpRI���@��%� 4@<v���!?v�=C�@�)����ٿ|D� ��@�T�"��3@ĳ0:��!?x��$��@�)����ٿ|D� ��@�T�"��3@ĳ0:��!?x��$��@��X2��ٿ��A-E��@�Xv�4@�'���!?b�u ��@�uçٿ#��&g��@UrP� 4@8����!?Q�d���@�uçٿ#��&g��@UrP� 4@8����!?Q�d���@�uçٿ#��&g��@UrP� 4@8����!?Q�d���@�uçٿ#��&g��@UrP� 4@8����!?Q�d���@�uçٿ#��&g��@UrP� 4@8����!?Q�d���@$��4�ٿǐʜ9��@���r.�3@^w�{f�!?��X���@$��4�ٿǐʜ9��@���r.�3@^w�{f�!?��X���@6lP1�ٿ��x�.��@��#� 4@(�G�0�!?6������@F�ů�ٿ5�n[*��@1����3@��h�P�!?�X#�z��@���
��ٿM�����@4����3@�����!?M�Rx��@���
��ٿM�����@4����3@�����!?M�Rx��@���
��ٿM�����@4����3@�����!?M�Rx��@б��n�ٿ�
�5�@P�H4@f�E�̏!?<ToUA�@б��n�ٿ�
�5�@P�H4@f�E�̏!?<ToUA�@б��n�ٿ�
�5�@P�H4@f�E�̏!?<ToUA�@б��n�ٿ�
�5�@P�H4@f�E�̏!?<ToUA�@б��n�ٿ�
�5�@P�H4@f�E�̏!?<ToUA�@�/.�ٿ��b$�@�ZI�4@6� %p�!?c�Y~��@�*,)ʙٿk��9�@�iɳ 4@�ん��!?(:��H�@�*,)ʙٿk��9�@�iɳ 4@�ん��!?(:��H�@�ԃ��ٿ�q ��@�/��A4@���\�!?G�?'�P�@�ԃ��ٿ�q ��@�/��A4@���\�!?G�?'�P�@�ԃ��ٿ�q ��@�/��A4@���\�!?G�?'�P�@����ٿ��3W,�@=��� 4@�Cbm�!?n}�@����ٿ��3W,�@=��� 4@�Cbm�!?n}�@����ٿ��3W,�@=��� 4@�Cbm�!?n}�@����ٿ��3W,�@=��� 4@�Cbm�!?n}�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@9�1a�ٿ�6�ģz�@ ���[ 4@m����!?��{\.�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�ꎗ��ٿ|��'77�@�R�� 4@(�s�ӏ!?4�]�@�A8[S�ٿ	u�5�@�Ob�p4@��0ŏ!?2�|�l�@�A8[S�ٿ	u�5�@�Ob�p4@��0ŏ!?2�|�l�@�A8[S�ٿ	u�5�@�Ob�p4@��0ŏ!?2�|�l�@�A8[S�ٿ	u�5�@�Ob�p4@��0ŏ!?2�|�l�@�A8[S�ٿ	u�5�@�Ob�p4@��0ŏ!?2�|�l�@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@I��*��ٿ�/$����@m�Hq�4@�(O ��!?W��bF��@��	��ٿ3H^fΞ�@]���3@�����!?��'�w��@��	��ٿ3H^fΞ�@]���3@�����!?��'�w��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@���cp�ٿ�ư�I��@�58i 4@^�G��!?��K��@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@�z��ٿ����N��@F�r� 4@)�^���!?25��7�@���
*�ٿ�^��d�@1t�Z� 4@m�z��!?������@��y�ٿr~I�@{��4@���!?s�Tl��@��y�ٿr~I�@{��4@���!?s�Tl��@��y�ٿr~I�@{��4@���!?s�Tl��@��y�ٿr~I�@{��4@���!?s�Tl��@��y�ٿr~I�@{��4@���!?s�Tl��@��y�ٿr~I�@{��4@���!?s�Tl��@-�`��ٿ�aRwW��@��h< 4@�����!? �()٩�@��Mv�ٿ�K��@���c4@�Xꆏ!?Y�h ���@��Mv�ٿ�K��@���c4@�Xꆏ!?Y�h ���@��Mv�ٿ�K��@���c4@�Xꆏ!?Y�h ���@�%";Ƨٿ����O�@��yWX4@�l�$��!?�SM�4�@�%";Ƨٿ����O�@��yWX4@�l�$��!?�SM�4�@?��ڥٿ/ߑ��@\J')� 4@��{�T�!?��B)�@\M^¤ٿn�M��@� �J4@������!?�E��V��@\M^¤ٿn�M��@� �J4@������!?�E��V��@�˲ڶ�ٿAŉx���@m�:-4@�1�>p�!?�J�v���@:�����ٿ�sp&�@���44@�<9Y@�!?��-���@:�����ٿ�sp&�@���44@�<9Y@�!?��-���@:�����ٿ�sp&�@���44@�<9Y@�!?��-���@�mn� �ٿ9w����@e�o�E 4@�|R�!?�d��L�@��&ڠٿF��bU�@�,h� 4@3Mr	S�!?�sʌ�@��&ڠٿF��bU�@�,h� 4@3Mr	S�!?�sʌ�@�ym/�ٿ��E8��@u�$�4@��4r�!?vv��@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@�*�v&�ٿqvk��^�@<��C4@�K�!?�Ý����@83M4�ٿ��/T��@�c�I� 4@G�I��!?f#\]@c�@83M4�ٿ��/T��@�c�I� 4@G�I��!?f#\]@c�@83M4�ٿ��/T��@�c�I� 4@G�I��!?f#\]@c�@83M4�ٿ��/T��@�c�I� 4@G�I��!?f#\]@c�@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@B�}军ٿ�ݨ?��@���^� 4@�MUv�!?�u-2m��@��H�B�ٿs��|��@���zW4@�5g�|�!?EN�D��@(��ml�ٿt1%��@O��J4@�=Oq�!?x�/&��@(��ml�ٿt1%��@O��J4@�=Oq�!?x�/&��@(��ml�ٿt1%��@O��J4@�=Oq�!?x�/&��@(��ml�ٿt1%��@O��J4@�=Oq�!?x�/&��@YEKh��ٿ���I�+�@Spz� 4@���!?n����@YEKh��ٿ���I�+�@Spz� 4@���!?n����@YEKh��ٿ���I�+�@Spz� 4@���!?n����@YEKh��ٿ���I�+�@Spz� 4@���!?n����@YEKh��ٿ���I�+�@Spz� 4@���!?n����@YEKh��ٿ���I�+�@Spz� 4@���!?n����@G0=ӗٿK�����@���4@���2^�!?�N���@G0=ӗٿK�����@���4@���2^�!?�N���@<��]Y�ٿ�Z�&�@��nq4@k��v�!?T}`��@<��]Y�ٿ�Z�&�@��nq4@k��v�!?T}`��@H]Yڿ�ٿ��ܒ�@Y��i4@��ס��!?g��a��@H]Yڿ�ٿ��ܒ�@Y��i4@��ס��!?g��a��@H]Yڿ�ٿ��ܒ�@Y��i4@��ס��!?g��a��@Lma��ٿA��d��@t��,4@�xh"P�!?s� ��t�@?��.έٿMO����@�i$�4@
R�!?��lL�4�@���}��ٿ*�eN�>�@�^��4@�����!?�0�@��(�	�ٿe�g�$��@����4@�W�Q`�!?.��/��@��(�	�ٿe�g�$��@����4@�W�Q`�!?.��/��@��(�	�ٿe�g�$��@����4@�W�Q`�!?.��/��@��(�	�ٿe�g�$��@����4@�W�Q`�!?.��/��@��(�	�ٿe�g�$��@����4@�W�Q`�!?.��/��@�ȣxǖٿN����@,F�Zr4@�g@h�!?�p߀���@c`�1�ٿ˧^��@�_R�4@�S��]�!?p��n��@c`�1�ٿ˧^��@�_R�4@�S��]�!?p��n��@c`�1�ٿ˧^��@�_R�4@�S��]�!?p��n��@c`�1�ٿ˧^��@�_R�4@�S��]�!?p��n��@L�u�ٿ^�����@��Ư� 4@K�Wc`�!?�c���@L�u�ٿ^�����@��Ư� 4@K�Wc`�!?�c���@L�u�ٿ^�����@��Ư� 4@K�Wc`�!?�c���@�ҙ�K�ٿB���/��@���4@�Շ�s�!?=صHJ�@0W�?�ٿ��ya[�@�G���3@W�r*܏!?8y��@��@C>_�ٿ8�e�;��@n�%t��3@ͮ�6��!?tw�-��@C>_�ٿ8�e�;��@n�%t��3@ͮ�6��!?tw�-��@C>_�ٿ8�e�;��@n�%t��3@ͮ�6��!?tw�-��@��9��ٿ�i��@�V��� 4@��P�!?wȹi�u�@�T'�ۓٿ	C9Be��@�:��g4@m�-��!?���<}�@�T'�ۓٿ	C9Be��@�:��g4@m�-��!?���<}�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@b��/��ٿ߲A�6�@#5?�F4@$'���!?�����{�@ie�s�ٿ[�A��@=A�� 4@��zp�!?�����^�@ie�s�ٿ[�A��@=A�� 4@��zp�!?�����^�@ie�s�ٿ[�A��@=A�� 4@��zp�!?�����^�@�j�#��ٿ�.8���@�3�i4@v�j��!?���:�X�@�j�#��ٿ�.8���@�3�i4@v�j��!?���:�X�@tѶ���ٿ'����@7�.6 4@u�D���!?I��˝��@tѶ���ٿ'����@7�.6 4@u�D���!?I��˝��@�5��w�ٿP�#3��@�j�;�3@�<#��!?<�d��u�@q����ٿ��N��@�`Ss 4@_��Ǐ!?A�1t'�@q����ٿ��N��@�`Ss 4@_��Ǐ!?A�1t'�@q����ٿ��N��@�`Ss 4@_��Ǐ!?A�1t'�@q����ٿ��N��@�`Ss 4@_��Ǐ!?A�1t'�@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�ɚխٿ����~��@�~�}��3@pV�׏!?����h��@�	7Jv�ٿG��k�@I�9�`4@z��`��!?
�8{q�@�	7Jv�ٿG��k�@I�9�`4@z��`��!?
�8{q�@��k,�ٿ��7�_��@w�:J%4@ӣ/@�!?F�ٯ}�@��k,�ٿ��7�_��@w�:J%4@ӣ/@�!?F�ٯ}�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@���`ߣٿ$��)��@޵;�O 4@�{�F�!?��zꎬ�@������ٿ�����@o��z�3@)K'�؏!?��?91�@������ٿ�����@o��z�3@)K'�؏!?��?91�@��&�ٿ����J�@�!!z�3@j/�F��!?Z+�RX��@��&�ٿ����J�@�!!z�3@j/�F��!?Z+�RX��@��&�ٿ����J�@�!!z�3@j/�F��!?Z+�RX��@!<�T�ٿ��JTy�@��W;��3@����!?E�QQ��@!<�T�ٿ��JTy�@��W;��3@����!?E�QQ��@�o��>�ٿ��`��W�@Jh%P�3@1��ŷ�!?�B>|f�@�o��>�ٿ��`��W�@Jh%P�3@1��ŷ�!?�B>|f�@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@^�҅��ٿ�N���-�@�j4@v9E�!?�Я����@ǳ�j��ٿ�M=8�.�@a���4@��PR�!?�)���B�@ǳ�j��ٿ�M=8�.�@a���4@��PR�!?�)���B�@ǳ�j��ٿ�M=8�.�@a���4@��PR�!?�)���B�@ǳ�j��ٿ�M=8�.�@a���4@��PR�!?�)���B�@ǳ�j��ٿ�M=8�.�@a���4@��PR�!?�)���B�@A�^�k�ٿ���q���@P?8h4@6N�V�!?�'T�_�@A�^�k�ٿ���q���@P?8h4@6N�V�!?�'T�_�@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@ѥLӹ�ٿ�k�����@ӥ�� 4@��u�!?5�/.��@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@��#M��ٿ��{���@���*��3@��)���!?���ߦ
�@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@�[��*�ٿ0%V���@�ˍ 4@%g��!?���,��@u_���ٿ��ך�@���4@%P��!?g:�ֱ��@Ե��*�ٿ�i��]��@�t[&e4@{l�d�!?TDc<�1�@Ե��*�ٿ�i��]��@�t[&e4@{l�d�!?TDc<�1�@�,Rf��ٿ}t�e�@?�Ҽ� 4@��m'ԏ!?����@�aq�׭ٿ�����@���+� 4@Tt1!Џ!?�;@��j�@�aq�׭ٿ�����@���+� 4@Tt1!Џ!?�;@��j�@�aq�׭ٿ�����@���+� 4@Tt1!Џ!?�;@��j�@�aq�׭ٿ�����@���+� 4@Tt1!Џ!?�;@��j�@�W���ٿc�_D��@�vЏ4@X~sU�!?HI�Z^[�@�W���ٿc�_D��@�vЏ4@X~sU�!?HI�Z^[�@�W���ٿc�_D��@�vЏ4@X~sU�!?HI�Z^[�@�W���ٿc�_D��@�vЏ4@X~sU�!?HI�Z^[�@�6?J�ٿ��1���@)��z� 4@&`Y���!?�T�B��@�/�.�ٿC:�2��@�ԉ4@���Տ!?�� ��@Z�Nnx�ٿ%%����@�K��14@���C��!?/&�%�@Z�Nnx�ٿ%%����@�K��14@���C��!?/&�%�@Z�Nnx�ٿ%%����@�K��14@���C��!?/&�%�@Z�Nnx�ٿ%%����@�K��14@���C��!?/&�%�@n�NɮٿO.xy���@�3�w4@{��Џ!?22
o��@n�NɮٿO.xy���@�3�w4@{��Џ!?22
o��@n�NɮٿO.xy���@�3�w4@{��Џ!?22
o��@Ѧ��@�ٿ�&�����@B�[�\4@8PϏ!?�֋����@F��&�ٿ�Y�J��@5���4@ƻ�J��!?*M��@F��&�ٿ�Y�J��@5���4@ƻ�J��!?*M��@��:�ٿŗ	���@ۋ��#4@w��!?�����@��:�ٿŗ	���@ۋ��#4@w��!?�����@��:�ٿŗ	���@ۋ��#4@w��!?�����@��:�ٿŗ	���@ۋ��#4@w��!?�����@�T�엱ٿ��^\T�@γ]�� 4@���r��!?/��q��@w�^x��ٿY�g�FO�@&/�C�4@c[�S��!?qk����@^H>m�ٿ�;��=�@ñb~��3@��1˯�!?��}q��@^H>m�ٿ�;��=�@ñb~��3@��1˯�!?��}q��@��Q�ٿe�^XX��@ EQ���3@N.&�я!?�Z[���@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�Ëg�ٿ^#���@���GH4@�Dl���!?�:հ-.�@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@�@G���ٿ�sQ9"��@L�a4@fKzZ�!?�6_���@@9���ٿNf�j��@���B4@��0u�!?~��}#�@@9���ٿNf�j��@���B4@��0u�!?~��}#�@@9���ٿNf�j��@���B4@��0u�!?~��}#�@@9���ٿNf�j��@���B4@��0u�!?~��}#�@@9���ٿNf�j��@���B4@��0u�!?~��}#�@t&E��ٿ���>�@��.� 4@wj+���!?`��2E�@t&E��ٿ���>�@��.� 4@wj+���!?`��2E�@t&E��ٿ���>�@��.� 4@wj+���!?`��2E�@t&E��ٿ���>�@��.� 4@wj+���!?`��2E�@t&E��ٿ���>�@��.� 4@wj+���!?`��2E�@9�cq]�ٿA5����@:ذ�*4@lǲ��!?81���@����ٿ�ϩ����@Õ'�� 4@���^�!?�hJ���@����ٿ�ϩ����@Õ'�� 4@���^�!?�hJ���@����ٿ�ϩ����@Õ'�� 4@���^�!?�hJ���@���BO�ٿ��k���@g!��� 4@sZj��!?�w�2��@���BO�ٿ��k���@g!��� 4@sZj��!?�w�2��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@zBL*��ٿvK��s�@�4hP�3@2?2���!?�Fs�R��@({��ٿ�n.����@��|�i�3@ʬ����!? ߨhS*�@({��ٿ�n.����@��|�i�3@ʬ����!? ߨhS*�@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@����ͧٿ�.���d�@ߏ�IY�3@}�ɏ!?��mH��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@�И�ٿO�˄��@+�2E�4@��%?ُ!?s�w�}��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@h�{���ٿ�g�J���@�t�`4@d�����!?�p�T��@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@���a��ٿ���q���@$��<4@p����!?����]�@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@;�qR�ٿ�S��1��@��7 4@$�&�ԏ!?|u$b`��@0��Sٝٿ��j%���@`F��� 4@"Ù
�!?�eK���@0��Sٝٿ��j%���@`F��� 4@"Ù
�!?�eK���@0��Sٝٿ��j%���@`F��� 4@"Ù
�!?�eK���@0��Sٝٿ��j%���@`F��� 4@"Ù
�!?�eK���@0��Sٝٿ��j%���@`F��� 4@"Ù
�!?�eK���@�H�r�ٿhg����@�����3@I����!?
���
N�@�H�r�ٿhg����@�����3@I����!?
���
N�@��ޮٿ� �i�@�����3@X��Џ!?�!->���@��ޮٿ� �i�@�����3@X��Џ!?�!->���@��ޮٿ� �i�@�����3@X��Џ!?�!->���@v����ٿhn��yk�@VxRǳ4@jEл�!?�%�P��@v����ٿhn��yk�@VxRǳ4@jEл�!?�%�P��@v����ٿhn��yk�@VxRǳ4@jEл�!?�%�P��@v����ٿhn��yk�@VxRǳ4@jEл�!?�%�P��@k-o�ٿERV�N�@�a����3@�П�!?�;b��h�@k�֡ٿu,��
��@�J���4@�u뇏!?$:����@N�\�ޞٿk�<en��@"�J|�4@$!|���!?�4	#��@�Oe��ٿ�Z�Ut_�@"��4@uw��g�!?Z����@�Oe��ٿ�Z�Ut_�@"��4@uw��g�!?Z����@�Oe��ٿ�Z�Ut_�@"��4@uw��g�!?Z����@�(LiԚٿ��a֏8�@j��V 4@�槮��!?IÒ��@�(LiԚٿ��a֏8�@j��V 4@�槮��!?IÒ��@�(LiԚٿ��a֏8�@j��V 4@�槮��!?IÒ��@�(LiԚٿ��a֏8�@j��V 4@�槮��!?IÒ��@�(LiԚٿ��a֏8�@j��V 4@�槮��!?IÒ��@s��lʕٿρ�-^�@%n�44@�u����!?y��l|��@s��lʕٿρ�-^�@%n�44@�u����!?y��l|��@s��lʕٿρ�-^�@%n�44@�u����!?y��l|��@�F�u��ٿՀ�-o��@����4@ṗ���!?xP�b�@�F�u��ٿՀ�-o��@����4@ṗ���!?xP�b�@�(WG8�ٿ�ǌ����@B�O��4@��.d��!?	E��.�@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@��œ3�ٿn^�\���@��� 4@�P<���!?���(��@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@D��{�ٿ�:�@���@9h*wx 4@FS�tb�!?�,����@����ٿV'����@j�>_.4@�]ڛW�!?��_$3�@����ٿV'����@j�>_.4@�]ڛW�!?��_$3�@����ٿV'����@j�>_.4@�]ڛW�!?��_$3�@����ٿV'����@j�>_.4@�]ڛW�!?��_$3�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@��?�ٿUͶ����@� J� 4@�즃x�!?T�b$U�@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@=-���ٿ�ћ㤕�@c�	� 4@\���a�!?�y�2��@S�5�ٿ�o���[�@W�;�b4@�KZ�7�!?��P��T�@S�5�ٿ�o���[�@W�;�b4@�KZ�7�!?��P��T�@r�0�חٿ+��St~�@���� 4@߈J��!? |����@r�0�חٿ+��St~�@���� 4@߈J��!? |����@r�0�חٿ+��St~�@���� 4@߈J��!? |����@
�j��ٿ�@J,�@�"u 4@�A�v�!?��^�7�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@�ᯍ��ٿֈ�:kN�@��0�;4@�M3�!?��Na�!�@%�J���ٿ�B�1��@��EH 4@����Џ!?�Ԩ+��@%�J���ٿ�B�1��@��EH 4@����Џ!?�Ԩ+��@���bQ�ٿm�3١��@��;���3@�~d��!?�!DK���@���bQ�ٿm�3١��@��;���3@�~d��!?�!DK���@���bQ�ٿm�3١��@��;���3@�~d��!?�!DK���@3锌�ٿ�|�I��@yc 4@�d��	�!?�"��W�@�~h͟ٿ�n�v��@L�{]E�3@�8�V��!?�e�2��@� Bہ�ٿ�r�����@����v�3@�\�e��!?	��Vd�@� Bہ�ٿ�r�����@����v�3@�\�e��!?	��Vd�@� Bہ�ٿ�r�����@����v�3@�\�e��!?	��Vd�@� Bہ�ٿ�r�����@����v�3@�\�e��!?	��Vd�@��Ѵ��ٿ��J���@t62٨�3@��Ï!?ʇ&F��@@��-��ٿr�Yg3��@�y�$4@+�e�Ώ!?Tnk2�E�@@��-��ٿr�Yg3��@�y�$4@+�e�Ώ!?Tnk2�E�@@��-��ٿr�Yg3��@�y�$4@+�e�Ώ!?Tnk2�E�@՝�ٛٿ&h�@d���4@U��Dۏ!?��Ǉ��@՝�ٛٿ&h�@d���4@U��Dۏ!?��Ǉ��@՝�ٛٿ&h�@d���4@U��Dۏ!?��Ǉ��@��"�ڠٿ��mXa�@ݯ�ݚ 4@q�p.��!?��Y��@��"�ڠٿ��mXa�@ݯ�ݚ 4@q�p.��!?��Y��@��"�ڠٿ��mXa�@ݯ�ݚ 4@q�p.��!?��Y��@��"�ڠٿ��mXa�@ݯ�ݚ 4@q�p.��!?��Y��@B�d�ٿ���@��@�'��H�3@�I櫉�!?k��7qz�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�]���ٿ'��Γ��@@Դ� 4@<P���!?���e�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@�e���ٿ� ��E`�@0�xh4@�Dg�^�!?��_J-l�@F�+Q@�ٿ��vW_9�@����4@hp�咏!?�qκ*��@F�+Q@�ٿ��vW_9�@����4@hp�咏!?�qκ*��@F�+Q@�ٿ��vW_9�@����4@hp�咏!?�qκ*��@F�+Q@�ٿ��vW_9�@����4@hp�咏!?�qκ*��@F�+Q@�ٿ��vW_9�@����4@hp�咏!?�qκ*��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@v�0W��ٿ�'�m��@�"4@v�.e�!?@c&��@o�..ڥٿ-ӽ����@ڞ�e`4@9T�71�!?�leў��@o�..ڥٿ-ӽ����@ڞ�e`4@9T�71�!?�leў��@o�..ڥٿ-ӽ����@ڞ�e`4@9T�71�!?�leў��@�Ct	I�ٿ�|�<�@/N�^� 4@2��4�!?G��%.�@�����ٿ����"�@��&�)4@*E�/8�!?cAm�I�@�h,y�ٿ��T�xP�@V���]4@�/�3��!?w��1d�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@ ���ٿX�L���@�Y&N 4@�-؏!?��f�@e�p�ٿ�S��g��@#��nm 4@����Џ!?�t��S�@e�p�ٿ�S��g��@#��nm 4@����Џ!?�t��S�@e�p�ٿ�S��g��@#��nm 4@����Џ!?�t��S�@��]�بٿf;
�p��@R"�N 4@'K{�Ï!?ζ�&��@��]�بٿf;
�p��@R"�N 4@'K{�Ï!?ζ�&��@i�p�6�ٿo�qz��@�n�� 4@�]�Y��!?U���8�@i�p�6�ٿo�qz��@�n�� 4@�]�Y��!?U���8�@i�p�6�ٿo�qz��@�n�� 4@�]�Y��!?U���8�@i�p�6�ٿo�qz��@�n�� 4@�]�Y��!?U���8�@��<}��ٿC��uZ{�@���Y� 4@�Q�x��!?�-h'k�@&���|�ٿ>ˍ����@km6�4@�5�H��!?q{�VV*�@&���|�ٿ>ˍ����@km6�4@�5�H��!?q{�VV*�@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@1u��ٿi�m��@�� 4@���׏!?p 
���@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@��ȥg�ٿ����@��H��4@3�ۡ��!?/�ư߰�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@�
��ٿ�0�Z��@Z�{(� 4@^c[��!?V`=�*�@��W�ٿsLn�E�@F�4@�C��!?e��p�c�@��W�ٿsLn�E�@F�4@�C��!?e��p�c�@[��ٿp=&Ʀ�@]N�(:4@�
g��!?��W궜�@[��ٿp=&Ʀ�@]N�(:4@�
g��!?��W궜�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@V�rӢٿk�Ҷ�R�@��U4@�_��!?e���K�@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@n<���ٿ�y}��@h6ti�4@y*V�p�!?;"���@`�B���ٿ�Ħ��@JvW��4@J�fg�!?^�ym)_�@�5�u�ٿXEYdۇ�@�/�S�4@޽��z�!?3��)\�@�5�u�ٿXEYdۇ�@�/�S�4@޽��z�!?3��)\�@�5�u�ٿXEYdۇ�@�/�S�4@޽��z�!?3��)\�@�mO��ٿ��8�\�@W-P8m 4@�b�{ُ!?�����@�mO��ٿ��8�\�@W-P8m 4@�b�{ُ!?�����@�mO��ٿ��8�\�@W-P8m 4@�b�{ُ!?�����@�mO��ٿ��8�\�@W-P8m 4@�b�{ُ!?�����@=$Z�ٿ�"�~�@��qE4@1�mЏ!?FP�r��@=$Z�ٿ�"�~�@��qE4@1�mЏ!?FP�r��@��o��ٿT?2�-�@�+��� 4@�o��ڏ!?`�[����@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@�pB�ٿ���ʷ�@�f 4@ق$��!?�9��{�@� C�G�ٿ�� �,�@�vV�=4@v����!?l`V�Js�@� C�G�ٿ�� �,�@�vV�=4@v����!?l`V�Js�@�sLē�ٿ��8M���@�
��- 4@�@��!?56w2��@�sLē�ٿ��8M���@�
��- 4@�@��!?56w2��@�sLē�ٿ��8M���@�
��- 4@�@��!?56w2��@�sLē�ٿ��8M���@�
��- 4@�@��!?56w2��@�sLē�ٿ��8M���@�
��- 4@�@��!?56w2��@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@ G�[S�ٿŀ�j��@�t��F 4@��o)��!?�
���@!�K�T�ٿ����N�@/$%WX 4@wTS���!?-k,O
�@���ٿwFU)[��@t0�� 4@9���!?#',�|�@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�ͮ֜ٿ�~&���@8�c6��3@,&��!?�͎� �@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@�л7�ٿ)ԁ@���@T�|I4@ʙǍt�!?Q�tHJ�@SGW�M�ٿ�A��@$p��(4@���Ώ!?�\��_��@�n}$��ٿ록�>�@��sS� 4@!S��$�!?Z�h��@�n}$��ٿ록�>�@��sS� 4@!S��$�!?Z�h��@��-�ٿS���c��@��B�x�3@�7й��!?٩V�x�@��-�ٿS���c��@��B�x�3@�7й��!?٩V�x�@1�  y�ٿ;퍵z�@d8C���3@��:噏!?C��+{��@�S�Q�ٿf�LԠ�@��BJT 4@?p��D�!?�Eg^mt�@E���ٿAӟM��@�k��? 4@����A�!?�?H���@E���ٿAӟM��@�k��? 4@����A�!?�?H���@�YG�ٿ��8N�V�@�/�L 4@z��^�!?�U�E`�@�YG�ٿ��8N�V�@�/�L 4@z��^�!?�U�E`�@&K�ٿ��>7w�@�����3@��}���!?��c�W�@&K�ٿ��>7w�@�����3@��}���!?��c�W�@&K�ٿ��>7w�@�����3@��}���!?��c�W�@&K�ٿ��>7w�@�����3@��}���!?��c�W�@�i����ٿ�%����@g�1h@4@���A�!?O<x�d^�@�7ڤٿ���i��@`����4@�1�`�!?����zJ�@�7ڤٿ���i��@`����4@�1�`�!?����zJ�@�7ڤٿ���i��@`����4@�1�`�!?����zJ�@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@��Ȍf�ٿ�J�В�@P��'\4@i`�'g�!?�I����@4�Y�ٿшގ��@��Za�4@�����!?i Nv.��@�.�L��ٿ�2X���@�eת 4@ɷw���!?�:����@�.�L��ٿ�2X���@�eת 4@ɷw���!?�:����@�.�L��ٿ�2X���@�eת 4@ɷw���!?�:����@�.�L��ٿ�2X���@�eת 4@ɷw���!?�:����@��u�ٿd�d���@���E4@fC���!?A�2����@]\�(\�ٿv�o��@r�t3j4@ѥk'V�!?��l��m�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@�z+{��ٿ� �@'�$4@R�.�2�!?aQz�)�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@!;>�r�ٿ
lԕ���@��R� 4@�A 5�!?��y>�Q�@����ٿh���c�@Iu�w4@�آ&9�!?���.]u�@����ٿh���c�@Iu�w4@�آ&9�!?���.]u�@����ٿh���c�@Iu�w4@�آ&9�!?���.]u�@����ٿh���c�@Iu�w4@�آ&9�!?���.]u�@����ٿh���c�@Iu�w4@�آ&9�!?���.]u�@�#@=��ٿZ�d� ��@�ň�4@�,b��!? 'D�ei�@�#@=��ٿZ�d� ��@�ň�4@�,b��!? 'D�ei�@�#@=��ٿZ�d� ��@�ň�4@�,b��!? 'D�ei�@!�	�ٿ8�&P�k�@��01� 4@�>0�!?j��,��@!�	�ٿ8�&P�k�@��01� 4@�>0�!?j��,��@!�	�ٿ8�&P�k�@��01� 4@�>0�!?j��,��@!�	�ٿ8�&P�k�@��01� 4@�>0�!?j��,��@��9䬢ٿӂ�w�@�����3@��`�)�!?f�T\��@��9䬢ٿӂ�w�@�����3@��`�)�!?f�T\��@��9䬢ٿӂ�w�@�����3@��`�)�!?f�T\��@��9䬢ٿӂ�w�@�����3@��`�)�!?f�T\��@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@봃TÝٿ�8���@z��C 4@�;$�ˏ!?{��(�;�@��
�ٿa�𦳙�@p�Uv��3@_����!?�%�?���@��
�ٿa�𦳙�@p�Uv��3@_����!?�%�?���@��
�ٿa�𦳙�@p�Uv��3@_����!?�%�?���@��
�ٿa�𦳙�@p�Uv��3@_����!?�%�?���@��
�ٿa�𦳙�@p�Uv��3@_����!?�%�?���@넉/��ٿ�'i�C��@1?��% 4@1���=�!?�v��Z��@U�
�O�ٿY�Hs�@U4�0 4@�DDS�!?n����@U�
�O�ٿY�Hs�@U4�0 4@�DDS�!?n����@�x'ߠٿI����@wY�M 4@f��US�!?�Ћ8g�@�x'ߠٿI����@wY�M 4@f��US�!?�Ћ8g�@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@��U�q�ٿ���\��@vu[���3@�'	>w�!?�,�ƺ��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@���O\�ٿ"Z�&�@ ?�� 4@i�^��!?C�\��@��aLi�ٿt������@�JO�^4@O��!?�M�I��@��aLi�ٿt������@�JO�^4@O��!?�M�I��@��aLi�ٿt������@�JO�^4@O��!?�M�I��@6���S�ٿ��M��@KI��(4@hX��!?��F�)�@6���S�ٿ��M��@KI��(4@hX��!?��F�)�@FGL���ٿ>Q
�d��@�*�?L4@�"ȿ�!?t6`Mߔ�@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@Xz[D$�ٿĚ���@j��Q�4@@]ӏ!?��U��@]ʖ�A�ٿK�P;���@V 9� 4@0Y@N�!?�u�H�@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@k��G�ٿ���T!��@R���q 4@����W�!?w5�֛��@s�eB�ٿ�A��_�@sd���3@�)�E�!?�`���@���)i�ٿZ�=,�@��v�3@�m���!?j�	�6?�@���)i�ٿZ�=,�@��v�3@�m���!?j�	�6?�@���)i�ٿZ�=,�@��v�3@�m���!?j�	�6?�@���)i�ٿZ�=,�@��v�3@�m���!?j�	�6?�@���)i�ٿZ�=,�@��v�3@�m���!?j�	�6?�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@��|�ٿ�,ՠ��@]�r��3@��o�Ǐ!?����/�@�0��ٿ��^F��@dK5k�3@a�����!?�Ʈ�\�@�0��ٿ��^F��@dK5k�3@a�����!?�Ʈ�\�@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@*����ٿEr5���@^�{4� 4@P�yCo�!?Z������@OUC
��ٿp3���@����4@CE���!?p(6!E�@��sٿh4����@¯���3@��5׏!?k\?����@��sٿh4����@¯���3@��5׏!?k\?����@�6��ɞٿ�>z��@싍��3@Ǯ�jˏ!?��T����@�6��ɞٿ�>z��@싍��3@Ǯ�jˏ!?��T����@�-[Ԡٿq�(���@-$��3@����я!?��kD���@�-[Ԡٿq�(���@-$��3@����я!?��kD���@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@�s�	�ٿ{w'�t��@���r�3@I<�ޏ!?TsUͽ�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��|vm�ٿ�a<� �@�	����3@�+ZC��!?����$�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@��Л�ٿ[B�?���@_K?� 4@j�����!?�&|�o�@ޓ��ٿ�:�J�@.m
�4@�ځ���!?#�+q�@���oz�ٿ��@�Cu�@��t�$4@=?OR�!?���g�u�@���oz�ٿ��@�Cu�@��t�$4@=?OR�!?���g�u�@���oz�ٿ��@�Cu�@��t�$4@=?OR�!?���g�u�@���oz�ٿ��@�Cu�@��t�$4@=?OR�!?���g�u�@���oz�ٿ��@�Cu�@��t�$4@=?OR�!?���g�u�@$
��ٿ�&&QFm�@��z5�4@��Mi#�!?��Z�nU�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@$�	�R�ٿW��b�j�@$�O�'�3@��B5G�!?�����A�@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@ql�*�ٿӆ�P4��@3����4@0�%'��!?����@t����ٿ�p��@Q�\���3@_��Cȏ!?g��UhM�@t����ٿ�p��@Q�\���3@_��Cȏ!?g��UhM�@t����ٿ�p��@Q�\���3@_��Cȏ!?g��UhM�@t����ٿ�p��@Q�\���3@_��Cȏ!?g��UhM�@t����ٿ�p��@Q�\���3@_��Cȏ!?g��UhM�@����ٿ��vQ�@z�jF�3@DL��!?���zH��@����ٿ��vQ�@z�jF�3@DL��!?���zH��@����ٿ��vQ�@z�jF�3@DL��!?���zH��@��?�3�ٿ��lm�6�@�+�[�3@�P�Y�!?ǝ5K1��@��?�3�ٿ��lm�6�@�+�[�3@�P�Y�!?ǝ5K1��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@�{ƃ7�ٿ�ޏ��@��Y��3@�r��q�!?/��77��@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@
W��ٿ�[�܋�@��� 4@u�n�a�!?���()�@��_ܢٿ���?���@�%�
4@�Z�R�!?�<���@��_ܢٿ���?���@�%�
4@�Z�R�!?�<���@u��4�ٿ_	o�t�@9D�#��3@�[�M�!?u�~��n�@u��4�ٿ_	o�t�@9D�#��3@�[�M�!?u�~��n�@u��4�ٿ_	o�t�@9D�#��3@�[�M�!?u�~��n�@�����ٿq�j�n�@HR)�C�3@�~�yY�!?O��iH�@�����ٿq�j�n�@HR)�C�3@�~�yY�!?O��iH�@�����ٿq�j�n�@HR)�C�3@�~�yY�!?O��iH�@�����ٿq�j�n�@HR)�C�3@�~�yY�!?O��iH�@�����ٿq�j�n�@HR)�C�3@�~�yY�!?O��iH�@n��&8�ٿ̏7��@�@$>���3@n��K�!?��2�r�@n��&8�ٿ̏7��@�@$>���3@n��K�!?��2�r�@n��&8�ٿ̏7��@�@$>���3@n��K�!?��2�r�@n��&8�ٿ̏7��@�@$>���3@n��K�!?��2�r�@�3B�ٿ ��O�o�@�|�a 4@�g�V�!?�6�0�@�3B�ٿ ��O�o�@�|�a 4@�g�V�!?�6�0�@�3B�ٿ ��O�o�@�|�a 4@�g�V�!?�6�0�@�3B�ٿ ��O�o�@�|�a 4@�g�V�!?�6�0�@�#�~�ٿI�Q�^�@BdZ���3@K�Ǐ!?e�M٘�@�#�~�ٿI�Q�^�@BdZ���3@K�Ǐ!?e�M٘�@c~i�ٿ�������@M��lS4@�<*'ُ!?�����?�@�1��'�ٿ�n��+z�@3�]�4@q8"��!?E���@�1��'�ٿ�n��+z�@3�]�4@q8"��!?E���@�1��'�ٿ�n��+z�@3�]�4@q8"��!?E���@�1��'�ٿ�n��+z�@3�]�4@q8"��!?E���@��� �ٿ+|a�v�@���% 4@ j3f�!?�bC
CX�@�Q:�ٿ��b7+��@)YQ4@DzU!��!?Wf�bX�@�Q:�ٿ��b7+��@)YQ4@DzU!��!?Wf�bX�@�Q:�ٿ��b7+��@)YQ4@DzU!��!?Wf�bX�@�Q:�ٿ��b7+��@)YQ4@DzU!��!?Wf�bX�@𘏖V�ٿ���=���@O��� 4@\N���!?3f �~��@𘏖V�ٿ���=���@O��� 4@\N���!?3f �~��@��6N�ٿJuA��,�@Ὼ6 4@�J{g�!?5���[��@��6N�ٿJuA��,�@Ὼ6 4@�J{g�!?5���[��@��6N�ٿJuA��,�@Ὼ6 4@�J{g�!?5���[��@��6N�ٿJuA��,�@Ὼ6 4@�J{g�!?5���[��@�>V�#�ٿ"0?0��@m�)�N 4@g��ў�!?q`c�m�@�>V�#�ٿ"0?0��@m�)�N 4@g��ў�!?q`c�m�@�>V�#�ٿ"0?0��@m�)�N 4@g��ў�!?q`c�m�@J��,�ٿ>L�&���@��a�\ 4@w�ᎏ!?�1�].T�@J��,�ٿ>L�&���@��a�\ 4@w�ᎏ!?�1�].T�@J��,�ٿ>L�&���@��a�\ 4@w�ᎏ!?�1�].T�@J��,�ٿ>L�&���@��a�\ 4@w�ᎏ!?�1�].T�@Et�J��ٿ4�%q�@G�*"e�3@v��a�!?&������@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@6��&I�ٿ��/v%�@�M���4@t���ŏ!?C�s��@Zd�샮ٿ��|�0��@���� 4@��!���!?�x�!jC�@���ٿ�Q[����@A��0�4@���ʏ!?�s'!��@���ٿ�Q[����@A��0�4@���ʏ!?�s'!��@���ٿ�Q[����@A��0�4@���ʏ!?�s'!��@���ٿ�Q[����@A��0�4@���ʏ!?�s'!��@j"Ix1�ٿ�������@�p�о4@�$ug��!?��@h��@j"Ix1�ٿ�������@�p�о4@�$ug��!?��@h��@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@�p}��ٿA�J���@����4@=���!?-OH�b�@��SIS�ٿ7!���@U��� 4@� ~�ޏ!?J.nwm�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�PcΣٿ�,�U��@�� 4@������!?.XP��C�@�N�[��ٿ~iP�W�@Z%��� 4@�� �ԏ!?��;��q�@�N�[��ٿ~iP�W�@Z%��� 4@�� �ԏ!?��;��q�@�N�[��ٿ~iP�W�@Z%��� 4@�� �ԏ!?��;��q�@�g3���ٿ�!��4�@#�g94@��f��!?�kR=�@�g3���ٿ�!��4�@#�g94@��f��!?�kR=�@�g3���ٿ�!��4�@#�g94@��f��!?�kR=�@�g3���ٿ�!��4�@#�g94@��f��!?�kR=�@�g3���ٿ�!��4�@#�g94@��f��!?�kR=�@���)ڛٿ��v+���@�޷m��3@ �5�!?L#��3]�@���)ڛٿ��v+���@�޷m��3@ �5�!?L#��3]�@�Uu�ٿ�+Z�D�@�����3@�����!?��>LC��@�Uu�ٿ�+Z�D�@�����3@�����!?��>LC��@�Uu�ٿ�+Z�D�@�����3@�����!?��>LC��@�Uu�ٿ�+Z�D�@�����3@�����!?��>LC��@�Uu�ٿ�+Z�D�@�����3@�����!?��>LC��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@(9 ���ٿ�Vo�4��@vQ�4@����!?�۠z��@�[��ٿ�����@�c�34@3���!?^�ܦp��@�[��ٿ�����@�c�34@3���!?^�ܦp��@�[��ٿ�����@�c�34@3���!?^�ܦp��@�[��ٿ�����@�c�34@3���!?^�ܦp��@�[��ٿ�����@�c�34@3���!?^�ܦp��@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@bE�|�ٿ8k���@�M��54@������!?X��E=[�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@(���ٿ�H��@߃�� 4@,��؏!?�Q��F�@lz���ٿ���\k��@QY�� 4@�F���!?6��pǙ�@lz���ٿ���\k��@QY�� 4@�F���!?6��pǙ�@l�ws�ٿ��O���@��,T�4@�>���!?{w�Ǆ��@l�ws�ٿ��O���@��,T�4@�>���!?{w�Ǆ��@l�ws�ٿ��O���@��,T�4@�>���!?{w�Ǆ��@i�;^��ٿ�cu�?�@����" 4@:\�k�!?�8h��N�@i�;^��ٿ�cu�?�@����" 4@:\�k�!?�8h��N�@�j��ٿ����L�@_l�� 4@6|a̏!?�
d���@�j��ٿ����L�@_l�� 4@6|a̏!?�
d���@)Z�
�ٿa�{S�@�@�o&# 4@�N��!?�{��@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@Bc֬�ٿ؆��I�@X02-?4@��,�ȏ!?�/��Kj�@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@)�e��ٿq�rs���@z?�J� 4@�cۏ!?&Y���@�W����ٿ�<�,��@�����4@�NE�Տ!?ޱ����@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@c�4`̢ٿ�%����@*�W>W4@���x�!?�eH�>�@��pgA�ٿ-��ݴ��@�<cF�4@�!ӏ!?-�z�@`�@�Q��g�ٿ2���p�@��*&� 4@f��(��!?����-�@�Q��g�ٿ2���p�@��*&� 4@f��(��!?����-�@�Q��g�ٿ2���p�@��*&� 4@f��(��!?����-�@�Q��g�ٿ2���p�@��*&� 4@f��(��!?����-�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@������ٿG;����@
�?34@ɽ�!?f!~I�@��}�ٿy����@a���B4@�16��!?X�SCй�@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@8� ���ٿ�6�����@�ͽ�D4@{�
��!?��R}r��@�ٲ4I�ٿ	�6��@�R��4@-�V\��!?D�!-I��@�ٲ4I�ٿ	�6��@�R��4@-�V\��!?D�!-I��@;����ٿL�����@�X�Ea 4@r�9�t�!?l��<�@�@;����ٿL�����@�X�Ea 4@r�9�t�!?l��<�@�@;����ٿL�����@�X�Ea 4@r�9�t�!?l��<�@�@;����ٿL�����@�X�Ea 4@r�9�t�!?l��<�@�@;����ٿL�����@�X�Ea 4@r�9�t�!?l��<�@�@����6�ٿ�k�d��@@ '4@�<�Y�!?0��E�e�@����6�ٿ�k�d��@@ '4@�<�Y�!?0��E�e�@���[�ٿ>vRJ���@}v�я 4@�k�3O�!?�Yz��@B?�!�ٿ��%6���@<���4@h�x�!?��k0D�@B?�!�ٿ��%6���@<���4@h�x�!?��k0D�@B?�!�ٿ��%6���@<���4@h�x�!?��k0D�@B?�!�ٿ��%6���@<���4@h�x�!?��k0D�@/����ٿq-�.)��@!�L	v4@ؾW��!?�����@/����ٿq-�.)��@!�L	v4@ؾW��!?�����@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@�~	�ٿ�y>h=��@-�Iz� 4@�7�!?�H�v��@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@ٟ��<�ٿ�T�����@��9�4@ �	w��!?8�_V���@|yߵٿ�}G�B��@���� 4@ϒ�̏!?��Vt\�@|yߵٿ�}G�B��@���� 4@ϒ�̏!?��Vt\�@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@ڤ���ٿ��PX ��@f8�x�4@7M��!?��ha���@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�s��ٿL���iy�@�8�u�4@�;���!?�3ʿ��@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�,���ٿ���E`��@6c&+4@�5��Y�!?8Z��\v�@�v����ٿ+�]���@Ė�c� 4@l ;���!?�3�_ �@�v����ٿ+�]���@Ė�c� 4@l ;���!?�3�_ �@�v����ٿ+�]���@Ė�c� 4@l ;���!?�3�_ �@�v����ٿ+�]���@Ė�c� 4@l ;���!?�3�_ �@�v����ٿ+�]���@Ė�c� 4@l ;���!?�3�_ �@���J��ٿP�Qzl��@3�]��4@g�	��!?�����@���J��ٿP�Qzl��@3�]��4@g�	��!?�����@^�J@k�ٿi�F��@�U���3@�:L��!?%/� ��@^�J@k�ٿi�F��@�U���3@�:L��!?%/� ��@^�J@k�ٿi�F��@�U���3@�:L��!?%/� ��@^�J@k�ٿi�F��@�U���3@�:L��!?%/� ��@XyƐ�ٿ�j�sH��@B��4@�Pd��!?��/!1�@XyƐ�ٿ�j�sH��@B��4@�Pd��!?��/!1�@��oL��ٿ�~���@����4@���ҏ!?�|��E�@��oL��ٿ�~���@����4@���ҏ!?�|��E�@��oL��ٿ�~���@����4@���ҏ!?�|��E�@��oL��ٿ�~���@����4@���ҏ!?�|��E�@��oL��ٿ�~���@����4@���ҏ!?�|��E�@*ao��ٿI����&�@�A|�N4@(爄�!?�Y��@��@*ao��ٿI����&�@�A|�N4@(爄�!?�Y��@��@��R9��ٿmy�s��@w�l.s�3@q�3�!?ΥTi��@��R9��ٿmy�s��@w�l.s�3@q�3�!?ΥTi��@�a;��ٿ�eh5:b�@��O��3@�/$c�!?�7�!2r�@�a;��ٿ�eh5:b�@��O��3@�/$c�!?�7�!2r�@�a;��ٿ�eh5:b�@��O��3@�/$c�!?�7�!2r�@�a;��ٿ�eh5:b�@��O��3@�/$c�!?�7�!2r�@��?��ٿYH��B��@Wd�8��3@9�Q]��!?�a�����@��?��ٿYH��B��@Wd�8��3@9�Q]��!?�a�����@��?��ٿYH��B��@Wd�8��3@9�Q]��!?�a�����@��?��ٿYH��B��@Wd�8��3@9�Q]��!?�a�����@��?��ٿYH��B��@Wd�8��3@9�Q]��!?�a�����@���#�ٿ�/ ���@d���4@cVM\I�!?�	(��S�@���#�ٿ�/ ���@d���4@cVM\I�!?�	(��S�@���#�ٿ�/ ���@d���4@cVM\I�!?�	(��S�@���#�ٿ�/ ���@d���4@cVM\I�!?�	(��S�@���#�ٿ��"���@���n4@?�6}��!?$��@$`�ƭٿ&6��Z��@�T��4@'=��]�!?�=i+ ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@׻s���ٿ�k�)*�@�� � 4@l��=!�!?��� ��@&����ٿO���
z�@�!\��4@��5J�!?�]����@b�����ٿ<�A���@��� $4@�w��=�!?�ζp�@�z�p��ٿn�?^�a�@�� 4@�,֥Y�!?�O7T5k�@�z�p��ٿn�?^�a�@�� 4@�,֥Y�!?�O7T5k�@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@W�����ٿU�@RV�@*`�i$4@79G���!?P��Ȱ��@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@)Gc���ٿH%[)Ԁ�@I';��4@��	˺�!?+������@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�:2�Q�ٿ�ֳB�@{ą�4@I�� ��!?�M�OT��@�;����ٿ�K1�@�w	���3@��z��!?3�VA�I�@�;����ٿ�K1�@�w	���3@��z��!?3�VA�I�@�;����ٿ�K1�@�w	���3@��z��!?3�VA�I�@�;����ٿ�K1�@�w	���3@��z��!?3�VA�I�@�b�q	�ٿ�H���@f�ew 4@�Q���!?�?9�i�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@t)ϡٿ �ł�t�@��H�7 4@x䨅��!?>�	�G�@�-�K]�ٿ^�[�ڷ�@�Zax��3@���ȏ!?dCR!���@�-�K]�ٿ^�[�ڷ�@�Zax��3@���ȏ!?dCR!���@�-�K]�ٿ^�[�ڷ�@�Zax��3@���ȏ!?dCR!���@�-�K]�ٿ^�[�ڷ�@�Zax��3@���ȏ!?dCR!���@�NU�W�ٿ_؃���@/�A<� 4@8@%X��!?�6�T��@�NU�W�ٿ_؃���@/�A<� 4@8@%X��!?�6�T��@�NU�W�ٿ_؃���@/�A<� 4@8@%X��!?�6�T��@�NU�W�ٿ_؃���@/�A<� 4@8@%X��!?�6�T��@�NU�W�ٿ_؃���@/�A<� 4@8@%X��!?�6�T��@�]d�:�ٿ��	@��@E�	�) 4@q�Ͱ�!?ȏĊ���@�]d�:�ٿ��	@��@E�	�) 4@q�Ͱ�!?ȏĊ���@�]d�:�ٿ��	@��@E�	�) 4@q�Ͱ�!?ȏĊ���@�]d�:�ٿ��	@��@E�	�) 4@q�Ͱ�!?ȏĊ���@�]d�:�ٿ��	@��@E�	�) 4@q�Ͱ�!?ȏĊ���@�n}�3�ٿ����@q4/J;4@�%�sS�!?`[��O�@�n}�3�ٿ����@q4/J;4@�%�sS�!?`[��O�@�n}�3�ٿ����@q4/J;4@�%�sS�!?`[��O�@�n}�3�ٿ����@q4/J;4@�%�sS�!?`[��O�@�n}�3�ٿ����@q4/J;4@�%�sS�!?`[��O�@�ņ�}�ٿ���n��@hO�:�4@�(8�N�!?����%�@D��l/�ٿ�`����@爙�� 4@�f�H�!?IT�W4�@D��l/�ٿ�`����@爙�� 4@�f�H�!?IT�W4�@D��l/�ٿ�`����@爙�� 4@�f�H�!?IT�W4�@�{���ٿc:,��&�@�%{;� 4@ȟ��\�!?����(�@�{���ٿc:,��&�@�%{;� 4@ȟ��\�!?����(�@�{���ٿc:,��&�@�%{;� 4@ȟ��\�!?����(�@�Nx�ٿb�16�@�u�4@Ӷ&R�!?��M�@�Nx�ٿb�16�@�u�4@Ӷ&R�!?��M�@�Nx�ٿb�16�@�u�4@Ӷ&R�!?��M�@�Nx�ٿb�16�@�u�4@Ӷ&R�!?��M�@�Nx�ٿb�16�@�u�4@Ӷ&R�!?��M�@!���ٿ�C����@����4@�l�j�!?B��O{��@|�P�ͨٿE�8�'��@;��E4@�~}�!?_��@�M�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@77
��ٿ܄7�C�@_�-?4@i򙥶�!?���4l�@�LA��ٿ[IwPX��@F��~��3@��ya�!?����D��@�LA��ٿ[IwPX��@F��~��3@��ya�!?����D��@�LA��ٿ[IwPX��@F��~��3@��ya�!?����D��@U�t ��ٿ��b���@���'�3@���]��!?�!����@U�t ��ٿ��b���@���'�3@���]��!?�!����@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@�f����ٿ�ٌh���@)H� 4@�>�7��!?㽫ET�@!��%�ٿ��/L��@���H	4@֒�C^�!?=d([���@!��%�ٿ��/L��@���H	4@֒�C^�!?=d([���@!��%�ٿ��/L��@���H	4@֒�C^�!?=d([���@!��%�ٿ��/L��@���H	4@֒�C^�!?=d([���@!��%�ٿ��/L��@���H	4@֒�C^�!?=d([���@����ͣٿ�/�z���@��:<G4@��ډď!?{�	RE�@����ͣٿ�/�z���@��:<G4@��ډď!?{�	RE�@����ͣٿ�/�z���@��:<G4@��ډď!?{�	RE�@@�Ow<�ٿ��yg*�@�'��4@K����!?�Q���@@�Ow<�ٿ��yg*�@�'��4@K����!?�Q���@@�Ow<�ٿ��yg*�@�'��4@K����!?�Q���@@�Ow<�ٿ��yg*�@�'��4@K����!?�Q���@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@����ٿ׵L���@*�]� 4@���O��!?��3�Cx�@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@�ACa
�ٿC�^��@YDF&g 4@l�&|ȏ!?�k!X���@݆ɨ�ٿH�q�	h�@�ԕ� 4@t#F���!?�ؿ8�6�@݆ɨ�ٿH�q�	h�@�ԕ� 4@t#F���!?�ؿ8�6�@cE�b�ٿ���(�@]�U^@�3@���w�!?�u����@cE�b�ٿ���(�@]�U^@�3@���w�!?�u����@cE�b�ٿ���(�@]�U^@�3@���w�!?�u����@cE�b�ٿ���(�@]�U^@�3@���w�!?�u����@cE�b�ٿ���(�@]�U^@�3@���w�!?�u����@s�G��ٿؘt����@9B���3@\�W�!?��7���@s�G��ٿؘt����@9B���3@\�W�!?��7���@	�s��ٿX���NZ�@��;� 4@.9�`�!?4B�?b�@	�s��ٿX���NZ�@��;� 4@.9�`�!?4B�?b�@	�s��ٿX���NZ�@��;� 4@.9�`�!?4B�?b�@�b�0��ٿ���>`a�@'	���3@��A:�!?b5T�@�b�0��ٿ���>`a�@'	���3@��A:�!?b5T�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@9�F���ٿ������@�҃�y 4@����!?ޒ�w_U�@�chR?�ٿ�\0Scc�@����3@Yh�UϏ!?�6�-N�@� ��Ơٿx�}���@�����3@]�b�ŏ!?v!�!��@� ��Ơٿx�}���@�����3@]�b�ŏ!?v!�!��@� ��Ơٿx�}���@�����3@]�b�ŏ!?v!�!��@� ��Ơٿx�}���@�����3@]�b�ŏ!?v!�!��@� ��Ơٿx�}���@�����3@]�b�ŏ!?v!�!��@Ax�R��ٿ V�"q��@*�[ 4@���i�!?�y�W���@Ax�R��ٿ V�"q��@*�[ 4@���i�!?�y�W���@��gG�ٿ�.b���@�k�� 4@ݨ�ϋ�!?j��ԇN�@��gG�ٿ�.b���@�k�� 4@ݨ�ϋ�!?j��ԇN�@��M��ٿ�������@A��,�4@K����!?y!��s�@��M��ٿ�������@A��,�4@K����!?y!��s�@��M��ٿ�������@A��,�4@K����!?y!��s�@��zsu�ٿ�~����@��&��3@����<�!?�sf���@��zsu�ٿ�~����@��&��3@����<�!?�sf���@�jv��ٿ��b��@[��ä�3@ײ;�r�!?�	���d�@�jv��ٿ��b��@[��ä�3@ײ;�r�!?�	���d�@�jv��ٿ��b��@[��ä�3@ײ;�r�!?�	���d�@!�#�o�ٿ%l*:���@�ÝT��3@	�kڍ�!?�"訜g�@!�#�o�ٿ%l*:���@�ÝT��3@	�kڍ�!?�"訜g�@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@1�+��ٿ��%=�@\ ����3@)���c�!?jJ{��@S���ٿ�=�
�@l�� ��3@{N�bW�!?��}�,�@��Y���ٿ�ޠ�`��@҃���3@~��pO�!?&�]�1k�@�,<�ٿ�3�Ѵ=�@�h�V��3@Qe�M!�!?�L�y�@�,<�ٿ�3�Ѵ=�@�h�V��3@Qe�M!�!?�L�y�@�,<�ٿ�3�Ѵ=�@�h�V��3@Qe�M!�!?�L�y�@A ��9�ٿ����'X�@�eF��3@m1i-"�!?I~H� �@r�Lf>�ٿ���=ݔ�@�jY 4@F����!?Y[ 7��@8R���ٿF�9v5�@�� 4@����!?u�� �h�@8R���ٿF�9v5�@�� 4@����!?u�� �h�@淓	,�ٿ�C��%�@z|ƞ�4@J�tq��!?�_��>�@����ٿ�#����@�Bf�4@βEB��!?���0�E�@����ٿ�#����@�Bf�4@βEB��!?���0�E�@����ٿ�#����@�Bf�4@βEB��!?���0�E�@Q2(��ٿ� �+X^�@o� (�4@�ծ��!?a�$��@Q2(��ٿ� �+X^�@o� (�4@�ծ��!?a�$��@Q2(��ٿ� �+X^�@o� (�4@�ծ��!?a�$��@Q2(��ٿ� �+X^�@o� (�4@�ծ��!?a�$��@2��?�ٿ6E�/�@l�,M4@Gd'�F�!?�z�)��@2��?�ٿ6E�/�@l�,M4@Gd'�F�!?�z�)��@2��?�ٿ6E�/�@l�,M4@Gd'�F�!?�z�)��@2��?�ٿ6E�/�@l�,M4@Gd'�F�!?�z�)��@��ӂ��ٿ�����@�h�4@L	B6+�!?J���1�@E����ٿ����@3�;4@���|i�!?Z]>� ��@E����ٿ����@3�;4@���|i�!?Z]>� ��@E����ٿ����@3�;4@���|i�!?Z]>� ��@,�Ĺ�ٿ��VeX��@��O,y�3@��xat�!?8�p��@,�Ĺ�ٿ��VeX��@��O,y�3@��xat�!?8�p��@,�Ĺ�ٿ��VeX��@��O,y�3@��xat�!?8�p��@,�Ĺ�ٿ��VeX��@��O,y�3@��xat�!?8�p��@��ܢٿ���Il�@�]&�&4@�N���!?�)Q�@��ܢٿ���Il�@�]&�&4@�N���!?�)Q�@�<�B�ٿ+j'$s��@��F�j4@���x�!?���;�@�<�B�ٿ+j'$s��@��F�j4@���x�!?���;�@�<�B�ٿ+j'$s��@��F�j4@���x�!?���;�@�e���ٿ���ƶ��@��nQ�4@�z����!?5"k4�O�@�e���ٿ���ƶ��@��nQ�4@�z����!?5"k4�O�@�e���ٿ���ƶ��@��nQ�4@�z����!?5"k4�O�@�e���ٿ���ƶ��@��nQ�4@�z����!?5"k4�O�@����ٿl��1���@\`�x4@	�a��!?u��Vn�@X�d�áٿU*���Q�@&�fW��3@K/�š�!?��&&��@X�d�áٿU*���Q�@&�fW��3@K/�š�!?��&&��@X�d�áٿU*���Q�@&�fW��3@K/�š�!?��&&��@X�d�áٿU*���Q�@&�fW��3@K/�š�!?��&&��@X�d�áٿU*���Q�@&�fW��3@K/�š�!?��&&��@�B��_�ٿV��N�~�@�� � 4@��ٴ�!?�3޴�N�@��'9��ٿ������@ *��4@!���!?���.��@��'9��ٿ������@ *��4@!���!?���.��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@����ٿ��*����@.�I�k 4@c��h�!?Y�J��@0i0xҬٿܘ����@�\��84@�nM�׏!?�
��4�@0i0xҬٿܘ����@�\��84@�nM�׏!?�
��4�@0i0xҬٿܘ����@�\��84@�nM�׏!?�
��4�@���Ë�ٿ#�����@Xs7��4@��C�!?m{�F�c�@�)���ٿ35��}��@+&�!4@����!?D��}�@�)���ٿ35��}��@+&�!4@����!?D��}�@�JQN�ٿ�>�ŀY�@��^�_ 4@;���ޏ!?�ZR����@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@X#r��ٿ%���t�@��C�4@�7	dޏ!?��&�4�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@�-���ٿ�`Q�@=�h])4@��3�_�!?���C)�@4�$M�ٿ��I�fy�@N�y��4@0R�P�!?X�T&ا�@4�$M�ٿ��I�fy�@N�y��4@0R�P�!?X�T&ا�@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��\>�ٿX����@y&��^4@�U�tP�!?���f��@��(��ٿ��d���@�M���3@O�K˝�!?P�h.2�@��(��ٿ��d���@�M���3@O�K˝�!?P�h.2�@��(��ٿ��d���@�M���3@O�K˝�!?P�h.2�@��(��ٿ��d���@�M���3@O�K˝�!?P�h.2�@��(��ٿ��d���@�M���3@O�K˝�!?P�h.2�@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@Ե)!�ٿ�[>�}�@�$����3@O��ϑ�!?�%�
��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@o�l�n�ٿ���+e(�@Aj����3@����!?� ��#��@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@tM|��ٿq��t���@ʛ����3@j�/���!?��.ay�@$r�p��ٿVDv��@�i�� 4@k�׬��!?����p�@$r�p��ٿVDv��@�i�� 4@k�׬��!?����p�@$r�p��ٿVDv��@�i�� 4@k�׬��!?����p�@$r�p��ٿVDv��@�i�� 4@k�׬��!?����p�@eq0�4�ٿ�g����@/Mۿ 4@��6�!?B\ki?�@:e/��ٿ�z�ւ�@c	�N�4@>��ϫ�!?`���چ�@��P�ٿB��P-�@<'��4@�	����!?�M��k�@��P�ٿB��P-�@<'��4@�	����!?�M��k�@��P�ٿB��P-�@<'��4@�	����!?�M��k�@��P�ٿB��P-�@<'��4@�	����!?�M��k�@��P�ٿB��P-�@<'��4@�	����!?�M��k�@�fXqX�ٿ���B,r�@N��4@�[��Ə!?�����@�fXqX�ٿ���B,r�@N��4@�[��Ə!?�����@�fXqX�ٿ���B,r�@N��4@�[��Ə!?�����@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@!�7��ٿ# ����@y/ld�4@G�nr�!?��\�C��@F!W�ٿ��t7__�@�v��4@G33$��!?��8z���@F!W�ٿ��t7__�@�v��4@G33$��!?��8z���@F!W�ٿ��t7__�@�v��4@G33$��!?��8z���@F!W�ٿ��t7__�@�v��4@G33$��!?��8z���@�S�ӭٿ���\P�@���� 4@f�GF
�!?֯x�v�@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@4=�E�ٿH�t�&��@\�Kn� 4@�>ް��!?*v"����@՞�L�ٿl@�:�@/S/4@���[��!?�iJ���@��"T�ٿ��D��@W��Y�4@�0ݕ�!?�
����@��"T�ٿ��D��@W��Y�4@�0ݕ�!?�
����@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@��~ţٿQ�~Q�@ĹrY4@(��ɥ�!?ђ��#A�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@�a,��ٿj스(��@m�I$4@,��w͏!?#Uq^�\�@k���K�ٿ�pI����@��ʄC 4@�G�&��!?�5��Y.�@k���K�ٿ�pI����@��ʄC 4@�G�&��!?�5��Y.�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@{�D�:�ٿh�2���@/�V� 4@UU�?y�!?@j�#nf�@�RsR%�ٿ��[4���@
��d 4@Y��̏!?;�o��@�RsR%�ٿ��[4���@
��d 4@Y��̏!?;�o��@�RsR%�ٿ��[4���@
��d 4@Y��̏!?;�o��@�RsR%�ٿ��[4���@
��d 4@Y��̏!?;�o��@�RsR%�ٿ��[4���@
��d 4@Y��̏!?;�o��@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@����ٿ�'�r�@�r��[ 4@t�H�!?¾���@�, `�ٿ}$t� �@�J�)4@�si༏!?0��;��@�, `�ٿ}$t� �@�J�)4@�si༏!?0��;��@��n�ٿ0�Q���@���<t 4@.h�I��!?(�W�-�@��n�ٿ0�Q���@���<t 4@.h�I��!?(�W�-�@��n�ٿ0�Q���@���<t 4@.h�I��!?(�W�-�@��n�ٿ0�Q���@���<t 4@.h�I��!?(�W�-�@X=�Tšٿ@7�\�@�Q;�04@�!\�֏!?PK)��@X=�Tšٿ@7�\�@�Q;�04@�!\�֏!?PK)��@���7�ٿ���+#�@R}u! 4@����!?9N����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@�u��n�ٿ��T���@a��ie 4@0b ��!?0H����@b���ըٿL,��[4�@vp4���3@ė�沏!?Y�=��@b���ըٿL,��[4�@vp4���3@ė�沏!?Y�=��@�@k�9�ٿ���ܟ�@�����3@�S����!?���m�@�@k�9�ٿ���ܟ�@�����3@�S����!?���m�@Ö4���ٿ?b�x,�@*�%��3@�Z��!?���x@|�@Ö4���ٿ?b�x,�@*�%��3@�Z��!?���x@|�@Ö4���ٿ?b�x,�@*�%��3@�Z��!?���x@|�@����C�ٿ�"c.��@�PC�3@�&aݏ!?zU�	��@W�
��ٿ����@�M��3@���>6�!?~�uvc.�@W�
��ٿ����@�M��3@���>6�!?~�uvc.�@W�
��ٿ����@�M��3@���>6�!?~�uvc.�@W�
��ٿ����@�M��3@���>6�!?~�uvc.�@���;�ٿ�DNI�@��1J�3@*��꬏!?w��l��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@k5��Z�ٿjc�g��@�C�'4@mG�҃�!?�8Z��@d�����ٿsN�A��@U�K�4@MQ��!? B 8��@>+8��ٿ��i͋�@���4@kJ� ��!?y�����@��N�ٿ�P��@^�+W 4@�/�ӏ!?�b ��@o���ٿ4���ƪ�@��t��3@�gd�!?�^;AJ��@˷��Тٿ����\�@�R�5�3@���1�!?����D�@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@= +��ٿT��U���@uV"4@���ڏ!?�����@�ê��ٿ�	_�<��@>�h1n 4@�ʙ��!?H��~���@�ê��ٿ�	_�<��@>�h1n 4@�ʙ��!?H��~���@�ê��ٿ�	_�<��@>�h1n 4@�ʙ��!?H��~���@�ê��ٿ�	_�<��@>�h1n 4@�ʙ��!?H��~���@�ê��ٿ�	_�<��@>�h1n 4@�ʙ��!?H��~���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@E_裣�ٿao�����@���� 4@�俏�!?.�a���@�0[�!�ٿV�'b�@Swg�4@�����!?K�m�r�@�0[�!�ٿV�'b�@Swg�4@�����!?K�m�r�@��!��ٿ%yy=���@�H�� 4@á�5��!?P�V����@��!��ٿ%yy=���@�H�� 4@á�5��!?P�V����@��!��ٿ%yy=���@�H�� 4@á�5��!?P�V����@z�uͧ�ٿ��� n�@�\<� 4@jX��x�!?�v��2?�@z�uͧ�ٿ��� n�@�\<� 4@jX��x�!?�v��2?�@z�uͧ�ٿ��� n�@�\<� 4@jX��x�!?�v��2?�@T]����ٿ�� ��|�@y�@>:�3@UNCi�!?'̥[�@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@M�Ӵ�ٿÆ�̀��@,'H���3@�T�t�!?DSc���@�;��%�ٿD3z�/n�@>�ݟ��3@����!?�w���%�@�;��%�ٿD3z�/n�@>�ݟ��3@����!?�w���%�@�;��%�ٿD3z�/n�@>�ݟ��3@����!?�w���%�@���s��ٿz��Qg3�@�� � 4@���Տ!?�0D�y^�@���s��ٿz��Qg3�@�� � 4@���Տ!?�0D�y^�@���s��ٿz��Qg3�@�� � 4@���Տ!?�0D�y^�@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@�N���ٿ.(��v�@f��x�3@v���{�!?�?����@��΋�ٿ�	/	�Y�@>��{�3@�ȸ�5�!?d�h����@��΋�ٿ�	/	�Y�@>��{�3@�ȸ�5�!?d�h����@��΋�ٿ�	/	�Y�@>��{�3@�ȸ�5�!?d�h����@��΋�ٿ�	/	�Y�@>��{�3@�ȸ�5�!?d�h����@��΋�ٿ�	/	�Y�@>��{�3@�ȸ�5�!?d�h����@���'�ٿ�����@ ��{4@�I3~�!?��v��Y�@���'�ٿ�����@ ��{4@�I3~�!?��v��Y�@���'�ٿ�����@ ��{4@�I3~�!?��v��Y�@���H��ٿ�,��.G�@��p 4@�*���!?�TF����@q����ٿo)F�@>0pUs4@:�8累!?h�$�@����ٿ��5���@��E;W4@S�^�Ϗ!?;��k�@�٪���ٿ��Q� Y�@뢅d4@�r�F��!?2��OQ�@�٪���ٿ��Q� Y�@뢅d4@�r�F��!?2��OQ�@��7�v�ٿ��Oo��@|��0�4@�Y{��!?Ѹ$�$�@��7�v�ٿ��Oo��@|��0�4@�Y{��!?Ѹ$�$�@��7�v�ٿ��Oo��@|��0�4@�Y{��!?Ѹ$�$�@��7�v�ٿ��Oo��@|��0�4@�Y{��!?Ѹ$�$�@��7�v�ٿ��Oo��@|��0�4@�Y{��!?Ѹ$�$�@E�2s�ٿ�#��g7�@i
��4@qP܏!?���"�@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�쀴��ٿ���/�@�P4@��",�!?�Ɣ&t��@�%�߳�ٿbxv�0�@QD�+�4@P��8��!?9,�n�J�@��Ǎ�ٿ��6H@�@+:*��3@9)���!?~Z ��@��Ǎ�ٿ��6H@�@+:*��3@9)���!?~Z ��@c�sެٿ����5�@ 3� 4@T����!?u}~�@c�sެٿ����5�@ 3� 4@T����!?u}~�@c�sެٿ����5�@ 3� 4@T����!?u}~�@c�sެٿ����5�@ 3� 4@T����!?u}~�@c�sެٿ����5�@ 3� 4@T����!?u}~�@�}9\��ٿ@��[s�@)X���4@(����!?M^u3t�@�}9\��ٿ@��[s�@)X���4@(����!?M^u3t�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@a�cm��ٿ�)���;�@I��#T 4@�����!?��f�@��嘮�ٿ�
d FV�@���54@�5����!?)޽b	��@��嘮�ٿ�
d FV�@���54@�5����!?)޽b	��@�aΤٿ��Z1g�@ŕ,�c4@D�oc�!?		ߣ�@�aΤٿ��Z1g�@ŕ,�c4@D�oc�!?		ߣ�@�aΤٿ��Z1g�@ŕ,�c4@D�oc�!?		ߣ�@�aΤٿ��Z1g�@ŕ,�c4@D�oc�!?		ߣ�@�aΤٿ��Z1g�@ŕ,�c4@D�oc�!?		ߣ�@9�����ٿߑ�:��@H�N 4@� y�2�!?��I��{�@9�����ٿߑ�:��@H�N 4@� y�2�!?��I��{�@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@��	�@�ٿ�C7��@;�0��3@�a�:�!?�i&H��@�DM�ߩٿᝒ�r��@��d]%�3@,q5���!?�z)��@L.b�ٿ,+��!�@*�#�:4@�vr�!?J	��i�@L.b�ٿ,+��!�@*�#�:4@�vr�!?J	��i�@L.b�ٿ,+��!�@*�#�:4@�vr�!?J	��i�@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@i�$��ٿ�@��h2�@,���4@oarU�!?K\�>7��@/� 3�ٿO����@\�4@�LR���!?�[��:@�@/� 3�ٿO����@\�4@�LR���!?�[��:@�@/� 3�ٿO����@\�4@�LR���!?�[��:@�@�|��h�ٿǤ��מ�@�<�w�4@�@�w�!?�D)�`��@�^���ٿ�W[
�@W���A 4@��׏!?G�j��+�@�^���ٿ�W[
�@W���A 4@��׏!?G�j��+�@�^���ٿ�W[
�@W���A 4@��׏!?G�j��+�@�^���ٿ�W[
�@W���A 4@��׏!?G�j��+�@l�eΰٿ)-7���@��B@ 4@��C�܏!?46��8�@l�eΰٿ)-7���@��B@ 4@��C�܏!?46��8�@l�eΰٿ)-7���@��B@ 4@��C�܏!?46��8�@l�eΰٿ)-7���@��B@ 4@��C�܏!?46��8�@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@1s��ˬٿ����|��@*eD�� 4@N*{��!?b�E_���@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@"��/��ٿj�����@'��9�4@���%��!?"a�f��@��=�f�ٿ�^�1�@�>uI4@۠��!?.G�����@��=�f�ٿ�^�1�@�>uI4@۠��!?.G�����@��=�f�ٿ�^�1�@�>uI4@۠��!?.G�����@��=�f�ٿ�^�1�@�>uI4@۠��!?.G�����@��=�f�ٿ�^�1�@�>uI4@۠��!?.G�����@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@@�U��ٿ�c���@[ar�W 4@I#���!?��̠RA�@��+�ȟٿ+��@�@(�7�4@��dOǏ!?�V���@��+�ȟٿ+��@�@(�7�4@��dOǏ!?�V���@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@����ٿ��t���@�/�4@�j�]��!?T4�� ��@*"�̝ٿ�ɷ���@I�Y�4@(���!?A�	���@*"�̝ٿ�ɷ���@I�Y�4@(���!?A�	���@*"�̝ٿ�ɷ���@I�Y�4@(���!?A�	���@*"�̝ٿ�ɷ���@I�Y�4@(���!?A�	���@*"�̝ٿ�ɷ���@I�Y�4@(���!?A�	���@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@�L���ٿ[�o�`��@֕I�4@'�9`ޏ!?h�g�o�@��x�ٿar�/Y��@1ѥE�4@�"��ُ!?�a��z��@��x�ٿar�/Y��@1ѥE�4@�"��ُ!?�a��z��@��x�ٿar�/Y��@1ѥE�4@�"��ُ!?�a��z��@��x�ٿar�/Y��@1ѥE�4@�"��ُ!?�a��z��@R�]dI�ٿе�]���@gu�.4@�r�!?��:;�@R�]dI�ٿе�]���@gu�.4@�r�!?��:;�@R�]dI�ٿе�]���@gu�.4@�r�!?��:;�@R�]dI�ٿе�]���@gu�.4@�r�!?��:;�@R�]dI�ٿе�]���@gu�.4@�r�!?��:;�@��(��ٿ@8^���@��k4@�B��!?M'�U�@��(��ٿ@8^���@��k4@�B��!?M'�U�@��(��ٿ@8^���@��k4@�B��!?M'�U�@�M�ٿ�y�� ��@��@r�4@����ӏ!?G"��_��@�M�ٿ�y�� ��@��@r�4@����ӏ!?G"��_��@{s�ǟ�ٿ��a.��@�x�D�4@���"�!?�S����@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@L�N��ٿ1�ǂN�@# 4@����Տ!?|�ᒻ��@�ܯ��ٿ�n�9��@#XW� 4@�i���!?IfJ�h��@�^v^6�ٿ�O�Ԍ9�@�<��o 4@�f��Տ!?�F��@�^v^6�ٿ�O�Ԍ9�@�<��o 4@�f��Տ!?�F��@�^v^6�ٿ�O�Ԍ9�@�<��o 4@�f��Տ!?�F��@�^v^6�ٿ�O�Ԍ9�@�<��o 4@�f��Տ!?�F��@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�6��y�ٿ������@0Kl{�3@�/έ�!?�:���@�[�娤ٿ"?^�8�@��� 4@e[��֏!?c�s9&�@�[�娤ٿ"?^�8�@��� 4@e[��֏!?c�s9&�@�[�娤ٿ"?^�8�@��� 4@e[��֏!?c�s9&�@�V��ٿ�ٖ=�@�
ٝ��3@�-���!?�h2|�m�@�V��ٿ�ٖ=�@�
ٝ��3@�-���!?�h2|�m�@�V��ٿ�ٖ=�@�
ٝ��3@�-���!?�h2|�m�@t؜�ٿ��$Q���@��M�9 4@���}��!?W�-:�U�@t؜�ٿ��$Q���@��M�9 4@���}��!?W�-:�U�@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@����k�ٿ;13����@�X.4@�ͤ �!?�l�0��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@z0SO��ٿ��A*��@mڥ& 4@v�7���!?5
�@��@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@
:��#�ٿ�����@���6g�3@�$K�!?OW�����@�$���ٿ��W�,��@5�����3@pw"�h�!?��w���@�$���ٿ��W�,��@5�����3@pw"�h�!?��w���@�$���ٿ��W�,��@5�����3@pw"�h�!?��w���@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@#y��ǚٿՓ"����@��ɛ' 4@h��妏!?<���1�@6�x��ٿ�K-��r�@%ҁ��3@yŨƏ!?�*6�D^�@6�x��ٿ�K-��r�@%ҁ��3@yŨƏ!?�*6�D^�@�n
��ٿv��H�@�]A�N4@���H��!?/��a-$�@hB��Y�ٿF�Gy�1�@���'4@�rvj��!?�$�F޴�@Hܷ�ٿ[�9�+�@g��9�4@f��!?�[}�$��@Hܷ�ٿ[�9�+�@g��9�4@f��!?�[}�$��@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@'S��M�ٿ�_Sc��@�j�c� 4@��t��!?t��Zh�@N��ٿI�@Z�	�@4�C��4@��R1��!?ScO~�x�@���Y��ٿ���$��@��vS��3@���I�!?*!�[���@���Y��ٿ���$��@��vS��3@���I�!?*!�[���@���Y��ٿ���$��@��vS��3@���I�!?*!�[���@���Y��ٿ���$��@��vS��3@���I�!?*!�[���@�D�J��ٿ�j@e�~�@����+�3@@�]))�!?#K&>[��@`����ٿ��14�@3%/F��3@,�7�>�!?�]_
I��@�5���ٿ]7zK��@� ���3@D�*^�!?C�M�t�@�5���ٿ]7zK��@� ���3@D�*^�!?C�M�t�@�5���ٿ]7zK��@� ���3@D�*^�!?C�M�t�@�5���ٿ]7zK��@� ���3@D�*^�!?C�M�t�@�5���ٿ]7zK��@� ���3@D�*^�!?C�M�t�@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@h9r7�ٿ��>K��@�5� 4@���a�!?x��.���@Xop�ٿ��;c�@�r�$4@[3��!?HGغ�K�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@u����ٿ�]r/��@����4@�I��ޏ!?M.Y6�9�@�d��ٿ�W5���@��f4@������!?j���@�d��ٿ�W5���@��f4@������!?j���@�d��ٿ�W5���@��f4@������!?j���@r�BA�ٿ�AOv�w�@aF�04@�!��!?��I_TV�@7�F6��ٿ�U�H�x�@�|��4@�(�Ə!?��`,-�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@�ۄ}�ٿc5:�\�@����H4@�.-��!?�>�BU�@��z+�ٿ^�	1w�@�KE��4@��S3��!?��D�@��z+�ٿ^�	1w�@�KE��4@��S3��!?��D�@��z+�ٿ^�	1w�@�KE��4@��S3��!?��D�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@�3��ٿ��9���@;z���3@������!?�&�ϡ�@u�,y�ٿ�G	��@	=1�� 4@j�я!?���2-�@u�,y�ٿ�G	��@	=1�� 4@j�я!?���2-�@u�,y�ٿ�G	��@	=1�� 4@j�я!?���2-�@u�,y�ٿ�G	��@	=1�� 4@j�я!?���2-�@I`[q�ٿ{�,i4��@߅����3@�=��!?i(L<o�@I`[q�ٿ{�,i4��@߅����3@�=��!?i(L<o�@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@AAg#�ٿ�" �{��@��q��3@,}z���!?�6��x��@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@�v�f��ٿ�M���y�@������3@A'����!?�ßseb�@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@+�t��ٿ����_O�@���4n�3@Fr����!?L��\���@E�����ٿ�]�L��@�z�� 4@�S,��!?`����a�@E�����ٿ�]�L��@�z�� 4@�S,��!?`����a�@E�����ٿ�]�L��@�z�� 4@�S,��!?`����a�@E�����ٿ�]�L��@�z�� 4@�S,��!?`����a�@E�����ٿ�]�L��@�z�� 4@�S,��!?`����a�@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@ϵ�V,�ٿ�S���@���9o 4@b3�ʏ!?A��=���@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@��D9�ٿ�刔��@�^��� 4@!�.ߗ�!?_7�(��@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@���ݟٿ����I�@4�U'��3@�Mi��!?��!����@j����ٿ�ۯf��@[~�ܒ�3@��	���!?������@j����ٿ�ۯf��@[~�ܒ�3@��	���!?������@j����ٿ�ۯf��@[~�ܒ�3@��	���!?������@j����ٿ�ۯf��@[~�ܒ�3@��	���!?������@[�vқٿg!;���@U�E�l4@	N��e�!?T'��D�@[�vқٿg!;���@U�E�l4@	N��e�!?T'��D�@[�vқٿg!;���@U�E�l4@	N��e�!?T'��D�@[�vқٿg!;���@U�E�l4@	N��e�!?T'��D�@[�vқٿg!;���@U�E�l4@	N��e�!?T'��D�@%��̞�ٿ��!B�w�@��p(4@��'��!?��.��@%��̞�ٿ��!B�w�@��p(4@��'��!?��.��@%��̞�ٿ��!B�w�@��p(4@��'��!?��.��@%��̞�ٿ��!B�w�@��p(4@��'��!?��.��@ˣ}.��ٿ�%�E\�@ 84��4@ waj�!?�*:�2�@��L4��ٿ�A�/��@ˁt@a�3@����]�!?@Q{���@��L4��ٿ�A�/��@ˁt@a�3@����]�!?@Q{���@��L4��ٿ�A�/��@ˁt@a�3@����]�!?@Q{���@��'�E�ٿ��fe��@�i�� 4@)d�'��!?���I��@��'�E�ٿ��fe��@�i�� 4@)d�'��!?���I��@��'�E�ٿ��fe��@�i�� 4@)d�'��!?���I��@�"a�ٿ�xS�Q�@�*t���3@��]�!?�A�{�@�"a�ٿ�xS�Q�@�*t���3@��]�!?�A�{�@�"a�ٿ�xS�Q�@�*t���3@��]�!?�A�{�@�"a�ٿ�xS�Q�@�*t���3@��]�!?�A�{�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@��Ĭٿ��q��@x��`H4@l~�5��!?,Lx�@3pM&��ٿ\��3�@Ƒ�D�4@�SO��!?$�c�V��@3pM&��ٿ\��3�@Ƒ�D�4@�SO��!?$�c�V��@3pM&��ٿ\��3�@Ƒ�D�4@�SO��!?$�c�V��@3pM&��ٿ\��3�@Ƒ�D�4@�SO��!?$�c�V��@3pM&��ٿ\��3�@Ƒ�D�4@�SO��!?$�c�V��@T7�?b�ٿ�t�e�@�ɤ 4@lnv���!?��(�@T7�?b�ٿ�t�e�@�ɤ 4@lnv���!?��(�@T7�?b�ٿ�t�e�@�ɤ 4@lnv���!?��(�@�Q��ٿ�WQ�/	�@P@+
4@�ϤUN�!?�ƕ�{��@�Q��ٿ�WQ�/	�@P@+
4@�ϤUN�!?�ƕ�{��@�Q��ٿ�WQ�/	�@P@+
4@�ϤUN�!?�ƕ�{��@��`��ٿ�����F�@��g	�4@�;46��!?�>��b�@�cW��ٿr����C�@�y�:4@U��0��!?8��ү(�@�cW��ٿr����C�@�y�:4@U��0��!?8��ү(�@�cW��ٿr����C�@�y�:4@U��0��!?8��ү(�@�cW��ٿr����C�@�y�:4@U��0��!?8��ү(�@�cW��ٿr����C�@�y�:4@U��0��!?8��ү(�@>���ٿ���/��@��mP4@��4&��!?�$ʫ?�@p�a���ٿs� ���@v���4@�Q=λ�!?(ӑ�v�@p�a���ٿs� ���@v���4@�Q=λ�!?(ӑ�v�@p�a���ٿs� ���@v���4@�Q=λ�!?(ӑ�v�@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@�X���ٿ���O���@6��4@<�oK�!?f��k��@&��@z�ٿ$%`��@"�5�4@9�����!?��9�e�@k�H�,�ٿ�q���@Ea��J4@,�����!?���-��@k�H�,�ٿ�q���@Ea��J4@,�����!?���-��@��՚ɰٿz)�����@)R� 4@��^��!?N�,�߸�@��՚ɰٿz)�����@)R� 4@��^��!?N�,�߸�@�eπ��ٿY���	`�@��n�� 4@
��F��!?��B�q��@�q
�5�ٿ�=�.Q�@�e8��4@��Տ!?4�<z$A�@ȭǇ�ٿLDVB\��@pa�F4@����ȏ!?ۤ�8��@ȭǇ�ٿLDVB\��@pa�F4@����ȏ!?ۤ�8��@ȭǇ�ٿLDVB\��@pa�F4@����ȏ!?ۤ�8��@ȭǇ�ٿLDVB\��@pa�F4@����ȏ!?ۤ�8��@��9jȟٿ
�sل��@3F��� 4@��ivʏ!?���f��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@!$'�ٿй�r��@��(�3@Z��2��!?m�T�x��@�r�3�ٿq�D+x�@��qZ�3@��#ջ�!?�����@�r�3�ٿq�D+x�@��qZ�3@��#ջ�!?�����@����,�ٿ�H�F��@Ӎ�)��3@�#�؏!?Ĩj�Y�@����,�ٿ�H�F��@Ӎ�)��3@�#�؏!?Ĩj�Y�@L�ȧ�ٿ(���	��@����3@,����!?�Y���L�@L�ȧ�ٿ(���	��@����3@,����!?�Y���L�@Ջ��ٿN�W����@������3@ 0&�ޏ!?I�T�"��@^��0�ٿ�=��Cj�@e���!�3@x�>D��!?ޤ��7�@^��0�ٿ�=��Cj�@e���!�3@x�>D��!?ޤ��7�@^��0�ٿ�=��Cj�@e���!�3@x�>D��!?ޤ��7�@^��0�ٿ�=��Cj�@e���!�3@x�>D��!?ޤ��7�@�����ٿמJ�+Y�@�ݸ�3@:mA�!?���(�@�����ٿמJ�+Y�@�ݸ�3@:mA�!?���(�@�����ٿמJ�+Y�@�ݸ�3@:mA�!?���(�@�����ٿמJ�+Y�@�ݸ�3@:mA�!?���(�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@&�����ٿ�M��0�@s�Mr@ 4@V�ϳ�!? ��$ S�@R�ңX�ٿ���`�@��1Z��3@�g�̏!?��Km��@]�?�ٿ��yÀ�@�{9� 4@GW���!?eOr��@]�?�ٿ��yÀ�@�{9� 4@GW���!?eOr��@]�?�ٿ��yÀ�@�{9� 4@GW���!?eOr��@]�?�ٿ��yÀ�@�{9� 4@GW���!?eOr��@kĺ݊�ٿh��I���@��j�%4@8'L���!?R�z����@������ٿRf���@)��v4@������!?m<|�I��@������ٿRf���@)��v4@������!?m<|�I��@������ٿRf���@)��v4@������!?m<|�I��@N�_'��ٿ7������@u����4@��l��!?��@�w�@N�_'��ٿ7������@u����4@��l��!?��@�w�@N�_'��ٿ7������@u����4@��l��!?��@�w�@N�_'��ٿ7������@u����4@��l��!?��@�w�@N�_'��ٿ7������@u����4@��l��!?��@�w�@\Qt�[�ٿ�"ZO�@�$T�n 4@N")V%�!?&�>g��@\Qt�[�ٿ�"ZO�@�$T�n 4@N")V%�!?&�>g��@\Qt�[�ٿ�"ZO�@�$T�n 4@N")V%�!?&�>g��@\Qt�[�ٿ�"ZO�@�$T�n 4@N")V%�!?&�>g��@�/N�ٿ���B�@B�П� 4@��n��!?�-\����@�/N�ٿ���B�@B�П� 4@��n��!?�-\����@�/N�ٿ���B�@B�П� 4@��n��!?�-\����@�/N�ٿ���B�@B�П� 4@��n��!?�-\����@e�N:4�ٿE\?{K�@C/�#4@-�#g�!?q�7W�F�@e�N:4�ٿE\?{K�@C/�#4@-�#g�!?q�7W�F�@e�N:4�ٿE\?{K�@C/�#4@-�#g�!?q�7W�F�@e�N:4�ٿE\?{K�@C/�#4@-�#g�!?q�7W�F�@e�N:4�ٿE\?{K�@C/�#4@-�#g�!?q�7W�F�@ͳvC��ٿ���$��@ 1�J4@�M.�ӏ!?��h����@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@P�Y2�ٿ�Y`��'�@���TJ4@�@c�!?��Z���@97=p�ٿ�VF��@Ui���3@�}?dۏ!?�0p6�@97=p�ٿ�VF��@Ui���3@�}?dۏ!?�0p6�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@uա�J�ٿ$�mq�@���ؼ 4@s�z���!?0��1zc�@���L��ٿ8���@b�@����� 4@������!?���w0�@���L��ٿ8���@b�@����� 4@������!?���w0�@�{bʨٿʆ�k���@5y�
[ 4@60���!?�6ME�P�@�{bʨٿʆ�k���@5y�
[ 4@60���!?�6ME�P�@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@�Z)bn�ٿ��YkY��@2.W� 4@]*�"y�!?:�I��@z6�8Ŭٿ����B�@P��d 4@���!��!?jR`*Dg�@z6�8Ŭٿ����B�@P��d 4@���!��!?jR`*Dg�@z6�8Ŭٿ����B�@P��d 4@���!��!?jR`*Dg�@ռaՓ�ٿ�A��]��@Hj|P��3@S
�]ҏ!?�w�'�@ռaՓ�ٿ�A��]��@Hj|P��3@S
�]ҏ!?�w�'�@�`��a�ٿ�:�nإ�@p*W�4@�2|Vp�!?L���.#�@�`��a�ٿ�:�nإ�@p*W�4@�2|Vp�!?L���.#�@�`��a�ٿ�:�nإ�@p*W�4@�2|Vp�!?L���.#�@�`��a�ٿ�:�nإ�@p*W�4@�2|Vp�!?L���.#�@�`��a�ٿ�:�nإ�@p*W�4@�2|Vp�!?L���.#�@5����ٿox�S�@6�њ�4@Yy4�M�!?�X ,3��@��5n֩ٿe���Z�@��d'_ 4@�{�Q�!?���	p��@��5n֩ٿe���Z�@��d'_ 4@�{�Q�!?���	p��@��5n֩ٿe���Z�@��d'_ 4@�{�Q�!?���	p��@�#�,ڝٿ���O�@��p�3@4���!?��&�}�@�L��W�ٿJ����@wߡsK4@^��!?Y���@�L��W�ٿJ����@wߡsK4@^��!?Y���@�L��W�ٿJ����@wߡsK4@^��!?Y���@�L��W�ٿJ����@wߡsK4@^��!?Y���@�L��W�ٿJ����@wߡsK4@^��!?Y���@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@%X��s�ٿ�?��L��@X�}�3@�M84}�!?���Q�@~�a��ٿ�E: �4�@ ϒ�<4@�s���!?���n��@U(�[v�ٿ�c�$�@�9�w�4@�{�7v�!?�
�K��@U(�[v�ٿ�c�$�@�9�w�4@�{�7v�!?�
�K��@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@ny�gL�ٿ �����@�����4@�Iq��!?E4�d;,�@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@�,����ٿ�N1x�+�@��T�94@wSdr��!?[׌����@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@%��e�ٿ��Cp�q�@J:;��4@���Y��!?̦�Z)�@�4SFm�ٿ�H�W��@7{���4@+����!?v5q��d�@�4SFm�ٿ�H�W��@7{���4@+����!?v5q��d�@�4SFm�ٿ�H�W��@7{���4@+����!?v5q��d�@6 vg�ٿVjt�9
�@�|�~��3@>��Ï!?�qX��u�@6 vg�ٿVjt�9
�@�|�~��3@>��Ï!?�qX��u�@6 vg�ٿVjt�9
�@�|�~��3@>��Ï!?�qX��u�@����y�ٿv�0���@H�t�3@t����!?x�skLI�@����y�ٿv�0���@H�t�3@t����!?x�skLI�@qDy�ٿ�k�*�@����3@�����!?�km
���@qDy�ٿ�k�*�@����3@�����!?�km
���@qDy�ٿ�k�*�@����3@�����!?�km
���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�vM��ٿ��q]��@B���3@SuZJ��!?�22C���@�fg_X�ٿ�Z�����@z�	" 4@��w"ۏ!?�ӟ����@�fg_X�ٿ�Z�����@z�	" 4@��w"ۏ!?�ӟ����@�fg_X�ٿ�Z�����@z�	" 4@��w"ۏ!?�ӟ����@�fg_X�ٿ�Z�����@z�	" 4@��w"ۏ!?�ӟ����@�fg_X�ٿ�Z�����@z�	" 4@��w"ۏ!?�ӟ����@�6`�ٿ��'��@�;>��3@��%ڏ!?�����[�@�6`�ٿ��'��@�;>��3@��%ڏ!?�����[�@�6`�ٿ��'��@�;>��3@��%ڏ!?�����[�@����Ŝٿ(�����@w�)ر4@������!?b�V��@��6��ٿjIe9Ux�@&����4@�>�"��!?eg|q�@��6��ٿjIe9Ux�@&����4@�>�"��!?eg|q�@h����ٿ���+���@���_ 4@#�\���!?|I�t�@h����ٿ���+���@���_ 4@#�\���!?|I�t�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@ %���ٿ�{�c^��@f���{ 4@�E��ȏ!?Uw���`�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@/F����ٿ�J[j��@`>w�j4@�⟏!?����R�@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@Y� Z�ٿ��ݐ���@�\�n� 4@ן��͏!?	I����@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@8{���ٿ��֫�K�@�W�4@'�&���!?޳~}T�@���ٿDCM�@�@� ��3@ZI�N�!?��]z	��@���ٿDCM�@�@� ��3@ZI�N�!?��]z	��@���ٿDCM�@�@� ��3@ZI�N�!?��]z	��@���ٿDCM�@�@� ��3@ZI�N�!?��]z	��@���ٿDCM�@�@� ��3@ZI�N�!?��]z	��@/=�E��ٿ������@Fb���3@���*,�!?Tn����@>�2v�ٿ��>a ��@K�Q�4@`�7�1�!?ŸO6k��@AYU�8�ٿ�_��0��@�f�� 4@��$�T�!?�����F�@�H�f�ٿ���L5��@Yg�L 4@�Ta�g�!?e50���@)'�&­ٿ�{"�Rq�@?���4@�r3���!?�igE���@)'�&­ٿ�{"�Rq�@?���4@�r3���!?�igE���@)'�&­ٿ�{"�Rq�@?���4@�r3���!?�igE���@�h6g�ٿ!�4��@pj!���3@XkK��!?���+�@�h6g�ٿ!�4��@pj!���3@XkK��!?���+�@�h6g�ٿ!�4��@pj!���3@XkK��!?���+�@�h6g�ٿ!�4��@pj!���3@XkK��!?���+�@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@���٫ٿ;��$j�@aAYR+�3@�uҥ�!?�(y��@�Nc;9�ٿ�H�����@�f����3@-xO,ҏ!?Y� ���@�Nc;9�ٿ�H�����@�f����3@-xO,ҏ!?Y� ���@�Nc;9�ٿ�H�����@�f����3@-xO,ҏ!?Y� ���@�Nc;9�ٿ�H�����@�f����3@-xO,ҏ!?Y� ���@>?#ѳٿ`H\_�@�ڏ�7 4@Y"+��!?�<dc��@>?#ѳٿ`H\_�@�ڏ�7 4@Y"+��!?�<dc��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@��uI�ٿ��5���@tH��4@Zd���!?��Yc*��@�ԇ�٨ٿL�jZ�@���7 4@�Rcs��!?���nͽ�@�ԇ�٨ٿL�jZ�@���7 4@�Rcs��!?���nͽ�@�o=�ۢٿ��9��@���p4@J%��i�!?��i^ˇ�@�o=�ۢٿ��9��@���p4@J%��i�!?��i^ˇ�@�o=�ۢٿ��9��@���p4@J%��i�!?��i^ˇ�@�o=�ۢٿ��9��@���p4@J%��i�!?��i^ˇ�@�c$�ٿ��G��@"W�j��3@�B�ӷ�!?C�"����@��E�ٿ<{�?��@k��d��3@��	�!?�ncA���@��E�ٿ<{�?��@k��d��3@��	�!?�ncA���@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@?��'�ٿ�x���@u���j4@�h�VϏ!?cV�����@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@��З�ٿK�6)��@�ND�4@��<3��!?/���	1�@GA�'�ٿ�|�5���@���4@�Ѣ�!?S�|���@T�}�ٿ�|��*�@[�~��4@@/�U��!? ��߼�@px��t�ٿ�h�&r0�@懝Y�3@����U�!?Z��D�P�@px��t�ٿ�h�&r0�@懝Y�3@����U�!?Z��D�P�@px��t�ٿ�h�&r0�@懝Y�3@����U�!?Z��D�P�@��F`�ٿ��O�j��@1n�V<�3@$�GR�!?g��#�@��F`�ٿ��O�j��@1n�V<�3@$�GR�!?g��#�@��F`�ٿ��O�j��@1n�V<�3@$�GR�!?g��#�@o�?<�ٿ�CG�,�@�{�s�3@ ��rM�!?4&K��i�@o�?<�ٿ�CG�,�@�{�s�3@ ��rM�!?4&K��i�@o�?<�ٿ�CG�,�@�{�s�3@ ��rM�!?4&K��i�@o�?<�ٿ�CG�,�@�{�s�3@ ��rM�!?4&K��i�@� ̛�ٿ�.����@��d 4@�x�ɟ�!?L_�C(�@� ̛�ٿ�.����@��d 4@�x�ɟ�!?L_�C(�@� ̛�ٿ�.����@��d 4@�x�ɟ�!?L_�C(�@� ̛�ٿ�.����@��d 4@�x�ɟ�!?L_�C(�@t� Y/�ٿY��[��@��E 4@#����!?P��%;��@t� Y/�ٿY��[��@��E 4@#����!?P��%;��@t� Y/�ٿY��[��@��E 4@#����!?P��%;��@t� Y/�ٿY��[��@��E 4@#����!?P��%;��@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@�O��	�ٿ���a�@��~�
 4@�bcEȏ!?��9�\S�@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@v�y���ٿ�ᾈ���@r��lr 4@*�(��!? �S���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@�Q\,��ٿ�ş!��@]B4�N�3@F�{.5�!?��n���@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@��D� �ٿm 9��g�@��l� 4@���A��!?�Îi��@z��}ڥٿ���^F�@�yO�+�3@����!?�qU����@z��}ڥٿ���^F�@�yO�+�3@����!?�qU����@�t.�r�ٿ�s�.p�@.��4@�'g���!?����@g��f�ٿ~:{�^�@�wfK�4@Z�\N��!?"8M5���@g��f�ٿ~:{�^�@�wfK�4@Z�\N��!?"8M5���@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@+��;�ٿ*�����@=��% 4@)_&U��!?F��>��@����ٿ':�x��@�~��h�3@	=�z��!?�c�����@����ٿ':�x��@�~��h�3@	=�z��!?�c�����@��g(��ٿ��[N��@��_R�3@V�Xˏ!?m��U�@
��19�ٿJ~���@eJg*&4@�x���!?��$,�Z�@
��19�ٿJ~���@eJg*&4@�x���!?��$,�Z�@
��19�ٿJ~���@eJg*&4@�x���!?��$,�Z�@��鐃�ٿ��$�&*�@`$�� 4@����u�!?P��m�@��o���ٿJ��@��@�v�04@<Uh!?|GʑO}�@��o���ٿJ��@��@�v�04@<Uh!?|GʑO}�@a�^�ٿ"��w���@YkC�4@�W���!?��× ��@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@ֈae�ٿ΄��Pp�@Ҙ�С 4@�i�'��!?�e�'�l�@|WO�ٿ��s��z�@K����3@�4�5!?��};���@u9hK9�ٿ=`��4��@�����3@�o���!?�Ļ]���@u9hK9�ٿ=`��4��@�����3@�o���!?�Ļ]���@u9hK9�ٿ=`��4��@�����3@�o���!?�Ļ]���@1�>��ٿ��k����@�`q�c�3@��)���!?7,`G"�@1�>��ٿ��k����@�`q�c�3@��)���!?7,`G"�@1�>��ٿ��k����@�`q�c�3@��)���!?7,`G"�@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@6�L1:�ٿ�o�����@tx̊�4@B$H�!?c#j*��@�
�l�ٿ����.I�@.�j%4@��lԏ!?�MZ�u�@�
�l�ٿ����.I�@.�j%4@��lԏ!?�MZ�u�@�
�l�ٿ����.I�@.�j%4@��lԏ!?�MZ�u�@	B�(`�ٿ�����C�@Ũ�"�4@3\�T�!?��ͼ��@	B�(`�ٿ�����C�@Ũ�"�4@3\�T�!?��ͼ��@	B�(`�ٿ�����C�@Ũ�"�4@3\�T�!?��ͼ��@ݰ�A��ٿ)PB��6�@��A�4@�uZ���!?5Vd�~�@ݰ�A��ٿ)PB��6�@��A�4@�uZ���!?5Vd�~�@ݰ�A��ٿ)PB��6�@��A�4@�uZ���!?5Vd�~�@�ixjU�ٿA�U�]��@���24@u�Xl��!?�# <��@�ixjU�ٿA�U�]��@���24@u�Xl��!?�# <��@�ixjU�ٿA�U�]��@���24@u�Xl��!?�# <��@�ixjU�ٿA�U�]��@���24@u�Xl��!?�# <��@�ߦ�7�ٿ���g�@� �Ը 4@|��{�!?��.���@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@w�]d�ٿZ�QT2�@����� 4@S�*L�!?��$�F��@5�n�k�ٿ4}��)��@�vnE� 4@�)��!?�����@S��_g�ٿ��?4���@aH�r4@�5����!?@�%'��@S��_g�ٿ��?4���@aH�r4@�5����!?@�%'��@S��_g�ٿ��?4���@aH�r4@�5����!?@�%'��@���È�ٿ7RM�d��@J']P�4@�v!x�!?�&��Yt�@���È�ٿ7RM�d��@J']P�4@�v!x�!?�&��Yt�@��`�ٿ�/�#>�@K�(�b4@ma�ُ!?'�DY�@��`�ٿ�/�#>�@K�(�b4@ma�ُ!?'�DY�@RP�ٿ��䆳�@gVl�3@i��뷏!?�VO�H�@RP�ٿ��䆳�@gVl�3@i��뷏!?�VO�H�@RP�ٿ��䆳�@gVl�3@i��뷏!?�VO�H�@T��-�ٿN;�����@��x�4@����!?�؅Hu=�@T��-�ٿN;�����@��x�4@����!?�؅Hu=�@sVќ�ٿ<���l��@<�b4@�{=��!?v�sT(��@�����ٿ��+��@�����4@Yka.��!?����7��@�����ٿ��+��@�����4@Yka.��!?����7��@�����ٿ��+��@�����4@Yka.��!?����7��@��2�G�ٿ�����@[�Ƌ 4@E7�Ui�!?�A��M�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@�/��I�ٿu�2n���@���K4@�4���!?��,�=�@t��\A�ٿ{�P�b��@X0�+�3@�MLƏ!?��(o���@t��\A�ٿ{�P�b��@X0�+�3@�MLƏ!?��(o���@t��\A�ٿ{�P�b��@X0�+�3@�MLƏ!?��(o���@&�h�M�ٿ�Y�6��@"��`��3@�=\ì�!?M��q���@&�h�M�ٿ�Y�6��@"��`��3@�=\ì�!?M��q���@&�h�M�ٿ�Y�6��@"��`��3@�=\ì�!?M��q���@&�h�M�ٿ�Y�6��@"��`��3@�=\ì�!?M��q���@*�\5��ٿx�삛�@��' 4@r\���!?���:���@*�\5��ٿx�삛�@��' 4@r\���!?���:���@ݾ��Ǟٿ�C�E��@vɤp�4@����!?�P.>��@ݾ��Ǟٿ�C�E��@vɤp�4@����!?�P.>��@ݾ��Ǟٿ�C�E��@vɤp�4@����!?�P.>��@ݾ��Ǟٿ�C�E��@vɤp�4@����!?�P.>��@�*L�ޣٿ������@�\!� 4@��4lΏ!?���|��@�*L�ޣٿ������@�\!� 4@��4lΏ!?���|��@�( "�ٿvQ:�&�@�3���4@���!?�U�5��@�( "�ٿvQ:�&�@�3���4@���!?�U�5��@���ٿ�\3�'��@8���4@�L�!?���	�@���ٿ�\3�'��@8���4@�L�!?���	�@���ٿ�\3�'��@8���4@�L�!?���	�@��p�ٿ�X���W�@m��$4@�7�!Ï!?/aJ��k�@��p�ٿ�X���W�@m��$4@�7�!Ï!?/aJ��k�@��p�ٿ�X���W�@m��$4@�7�!Ï!?/aJ��k�@� ���ٿ�@�i���@O��(�4@��Є�!?�����@� ���ٿ�@�i���@O��(�4@��Є�!?�����@cN��ٿc]���@���u4@/#-g��!?����A�@cN��ٿc]���@���u4@/#-g��!?����A�@cN��ٿc]���@���u4@/#-g��!?����A�@cN��ٿc]���@���u4@/#-g��!?����A�@cN��ٿc]���@���u4@/#-g��!?����A�@cN��ٿc]���@���u4@/#-g��!?����A�@�˪�ٿb�k�_�@G_$��4@��G�ӏ!?f���t��@�KJg�ٿPN.����@�*��D4@C�Gp��!?�8u��@�KJg�ٿPN.����@�*��D4@C�Gp��!?�8u��@�KJg�ٿPN.����@�*��D4@C�Gp��!?�8u��@�KJg�ٿPN.����@�*��D4@C�Gp��!?�8u��@�����ٿ���>�@��n��4@b����!?at<&�X�@�(s�8�ٿ]cV���@L9�JN4@��Y��!?����wy�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@3(��ٿ:���o�@y��. 4@ٷ���!?q1�Ld�@��h�ٿ9$Q�/�@���24@�J���!?!t(p���@��h�ٿ9$Q�/�@���24@�J���!?!t(p���@�ҫcp�ٿ��BuX^�@�zA�4@?jw���!?�U�(��@�ҫcp�ٿ��BuX^�@�zA�4@?jw���!?�U�(��@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@G.����ٿ�p^����@�J�k�4@&N��!?��7^ӈ�@���ӛٿ��3+���@jF`�w4@�).�z�!?�
��{�@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@�Ɖ�ٿ���T�@�n#�r4@�ݤ��!?� ����@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@5)2qޞٿM��p@��@�[.� 4@j�6��!?rg+(��@N��ٿE���#�@�F�� 4@2{�l�!?��2c���@N��ٿE���#�@�F�� 4@2{�l�!?��2c���@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@��M�ٿ���&i,�@�R��� 4@��ױ�!?�^�:�-�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�ǘ䈫ٿw%�Y�@ H,�Q 4@��fo��!?�~�4v�@�}.J��ٿZVި��@3\�޳�3@�D����!?֋�yu'�@�}.J��ٿZVި��@3\�޳�3@�D����!?֋�yu'�@�}.J��ٿZVި��@3\�޳�3@�D����!?֋�yu'�@