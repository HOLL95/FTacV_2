�NUMPY v {'descr': '<f8', 'fortran_order': False, 'shape': (3, 10000, 5), }                                                   
������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@b�Ԇƙٿ7������@a�u 4@� ?�Ր!?�k��(��@e����ٿY�����@��4{ 4@X���C�!?����(��@e����ٿY�����@��4{ 4@X���C�!?����(��@e����ٿY�����@��4{ 4@X���C�!?����(��@e����ٿY�����@��4{ 4@X���C�!?����(��@e����ٿY�����@��4{ 4@X���C�!?����(��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@�Xߨ��ٿ���b���@���� 4@"�%3�!?.�Xm)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@1	���ٿ�׏e���@Ё�� 4@��ȣ�!?��6S)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@%n�]�ٿj����@蕉� 4@���!?E@W)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@k����ٿ�р���@���� 4@��Ő!?[�.V)��@�$vAڙٿ}܁���@=<�� 4@I��%�!?�RhL)��@9�ʙٿ�&����@�� 4@��o���!?��j4)��@9�ʙٿ�&����@�� 4@��o���!?��j4)��@9�ʙٿ�&����@�� 4@��o���!?��j4)��@ȟq;ʙٿ����@���� 4@�@�8�!?�{()��@ȟq;ʙٿ����@���� 4@�@�8�!?�{()��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@ag��ϙٿ�/T���@�x- 4@��R��!?���*)��@���əٿ��kx���@毜N 4@eo����!?7�I.)��@���əٿ��kx���@毜N 4@eo����!?7�I.)��@���əٿ��kx���@毜N 4@eo����!?7�I.)��@���əٿ��kx���@毜N 4@eo����!?7�I.)��@���əٿ��kx���@毜N 4@eo����!?7�I.)��@F}�>Ιٿ��x���@x+�� 4@6�I��!?��x)��@F}�>Ιٿ��x���@x+�� 4@6�I��!?��x)��@F}�>Ιٿ��x���@x+�� 4@6�I��!?��x)��@F}�>Ιٿ��x���@x+�� 4@6�I��!?��x)��@F}�>Ιٿ��x���@x+�� 4@6�I��!?��x)��@�U�ϙٿ�K v���@��' 4@�T�ϐ!?"�{')��@�U�ϙٿ�K v���@��' 4@�T�ϐ!?"�{')��@�U�ϙٿ�K v���@��' 4@�T�ϐ!?"�{')��@�\�͙ٿh�7x���@7/�n 4@D�5���!?��()��@�\�͙ٿh�7x���@7/�n 4@D�5���!?��()��@�\�͙ٿh�7x���@7/�n 4@D�5���!?��()��@�\�͙ٿh�7x���@7/�n 4@D�5���!?��()��@�\�͙ٿh�7x���@7/�n 4@D�5���!?��()��@���<Ιٿ�o|{���@�T�� 4@��O�!?S�y&)��@���<Ιٿ�o|{���@�T�� 4@��O�!?S�y&)��@�%Gҙٿ�o���@WU"� 4@. ���!?��3)��@�?��ҙٿ�x�h���@n��b 4@(h��d�!?�e9)��@�?��ҙٿ�x�h���@n��b 4@(h��d�!?�e9)��@ �hRٙٿ�F�g���@���n 4@�ӭ��!? [%>)��@_/�ߙٿB�>g���@��� 4@|+�p��!?YF;)��@_/�ߙٿB�>g���@��� 4@|+�p��!?YF;)��@_/�ߙٿB�>g���@��� 4@|+�p��!?YF;)��@_/�ߙٿB�>g���@��� 4@|+�p��!?YF;)��@_/�ߙٿB�>g���@��� 4@|+�p��!?YF;)��@"R2J��ٿ�#g���@ލz 4@YI�`>�!?��"4)��@UD�ڙٿ� l���@�o�� 4@^٨M�!?r�9)��@��4#�ٿ�V�h���@�G�9 4@߼��q�!?~�=)��@��R��ٿ�fmg���@;��3 4@�`hu�!?A�:;)��@��R��ٿ�fmg���@;��3 4@�`hu�!?A�:;)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@�*е�ٿ��m���@Đjs 4@�W�uܐ!?;�@?)��@��)�ٿ,-l���@iߗ 4@Kpa�ߐ!?�^N5)��@,���ٿ��m���@��� 4@�,dN��!? 5G:)��@E+�g�ٿb�*r���@�֑ 4@�ĩ�!?q��:)��@�Κ	�ٿ��py���@���� 4@��ժ�!?v��:)��@�Κ	�ٿ��py���@���� 4@��ժ�!?v��:)��@�Κ	�ٿ��py���@���� 4@��ժ�!?v��:)��@�nd��ٿY2gx���@�'ߘ 4@����!?��=)��@�5GP�ٿN�����@��P� 4@de��Ґ!?<-�A)��@�5GP�ٿN�����@��P� 4@de��Ґ!?<-�A)��@�4�ٿЊ�z���@��U� 4@B'榲�!?$�CA)��@���ٿ�0�r���@�� 4@��U���!?sbWF)��@���ٿ�0�r���@�� 4@��U���!?sbWF)��@��V��ٿ��Gx���@�Կ 4@9�T̐!?��D)��@޵�h��ٿ�/�w���@\O� 4@ޡ���!?]�E)��@֫}��ٿ�Si{���@D$tM 4@��$���!?�?)��@֫}��ٿ�Si{���@D$tM 4@��$���!?�?)��@֫}��ٿ�Si{���@D$tM 4@��$���!?�?)��@֫}��ٿ�Si{���@D$tM 4@��$���!?�?)��@֫}��ٿ�Si{���@D$tM 4@��$���!?�?)��@xj��ٿW��}���@H7� 4@~l��!?��A)��@ڏl�ٿS������@$Lw� 4@-�#>��!?�j�B)��@��;8��ٿ�t����@ � 4@]�]~�!?�ޝ>)��@*5���ٿ�SF����@�5 _ 4@���mX�!?WK<)��@*5���ٿ�SF����@�5 _ 4@���mX�!?WK<)��@kB��ٿQ����@xц 4@��=�!?m>5)��@,	���ٿ�BO����@QP!� 4@���*�!?;��2)��@,	���ٿ�BO����@QP!� 4@���*�!?;��2)��@,	���ٿ�BO����@QP!� 4@���*�!?;��2)��@T����ٿ6=_����@��� 4@��P9�!?UM8)��@�;#�ٿp ����@��m� 4@�����!?��9)��@�UUv��ٿ��%z���@��� 4@6s�0�!?n�x9)��@�T<��ٿ°�w���@�$L% 4@ͬ�5_�!?�(�8)��@�~���ٿs1�v���@�^ 4@�Ck�!?��2)��@�~���ٿs1�v���@�^ 4@�Ck�!?��2)��@����ٿR�s���@f�� 4@�tIl�!?��5)��@����ٿR�s���@f�� 4@�tIl�!?��5)��@!�I�ٿ�+ts���@}�} 4@і�F��!?^Z!8)��@#9O	�ٿ@`�p���@���9 4@���*�!?���6)��@#9O	�ٿ@`�p���@���9 4@���*�!?���6)��@��
5	�ٿ���r���@y�X� 4@a�R/��!?p��3)��@xI_�ٿ�O�p���@B,l 4@ ڣ�!?�Ȫ4)��@xI_�ٿ�O�p���@B,l 4@ ڣ�!?�Ȫ4)��@��	�ٿ�#�r���@�b�� 4@J��8Ő!?Oa)5)��@�9�}�ٿj�t���@�Um� 4@�C�ΐ!?˝95)��@3�V��ٿҘ�p���@(�F 4@��֔�!?@o^8)��@�襦�ٿo��m���@���� 4@�I��!?� "9)��@�襦�ٿo��m���@���� 4@�I��!?� "9)��@����ٿS��q���@��ͮ 4@����!?�&+:)��@�J���ٿ7��t���@:H7 4@����!?�$�5)��@Ix��ٿ���x���@m�x� 4@�+�2��!?��$6)��@Ix��ٿ���x���@m�x� 4@�+�2��!?��$6)��@Ix��ٿ���x���@m�x� 4@�+�2��!?��$6)��@C��<�ٿ}�t���@c{�� 4@�J:£�!?�O�3)��@ɑ�+�ٿ�J"v���@A�� 4@�>4�Ր!?Q�M9)��@�tC�ٿ���v���@V�� 4@����!??0�A)��@��k�ٿ!
}y���@7��Y 4@y�̾א!?̲�<)��@��k�ٿ!
}y���@7��Y 4@y�̾א!?̲�<)��@h���ٿ*�zw���@Cu� 4@�,Z�D�!?`S�:)��@s@m��ٿJ��v���@�� 4@��a0�!?�:)��@<�D�ٿ�y"s���@]�8� 4@̫_�.�!?��8<)��@�ۦ�ٿ w%s���@.�� 4@
�y��!?��=?)��@�HJ��ٿ��am���@��,� 4@��uS�!?��H?)��@�����ٿ�Ij���@��}' 4@
�O,�!?�m�B)��@:���ٿp_Dj���@���� 4@̜א�!?��B)��@���]�ٿ�r6g���@�i�q 4@q�}�!?��=C)��@ {[��ٿ���d���@�A� 4@�K��!?��:A)��@ɱ4t�ٿ�l���@J�G' 4@�j~�!?�IA)��@M
���ٿܔ�m���@�_�D 4@>O�ϐ!?�l>)��@M
���ٿܔ�m���@�_�D 4@>O�ϐ!?�l>)��@M
���ٿܔ�m���@�_�D 4@>O�ϐ!?�l>)��@����ٿ�}ue���@��N 4@o���!? |@)��@�4@��ٿ/;Va���@F`�� 4@G����!?�S�A)��@$��+�ٿ��_���@ݹyb 4@����!?���B)��@$��+�ٿ��_���@ݹyb 4@����!?���B)��@e��+�ٿ�c���@v*F 4@�.6��!?v��@)��@e��+�ٿ�c���@v*F 4@�.6��!?v��@)��@6�L�.�ٿ�s�Z���@"Y 4@y��^ː!?�>)��@6�L�.�ٿ�s�Z���@"Y 4@y��^ː!?�>)��@�E�=@�ٿ�2�U���@��� 4@\m�)֐!?9�@)��@�bDA�ٿ{�tV���@�QS� 4@�yM�Ɛ!?(�=)��@,/x�?�ٿN�Q���@_' 4@�2.iސ!?˯/>)��@�&lNM�ٿ�YQI���@!S[� 4@*�/��!?�7iA)��@�� ;�ٿ�}�O���@�d� 4@&�����!?�SFA)��@�� ;�ٿ�}�O���@�d� 4@&�����!?�SFA)��@AI�N�ٿ�C1N���@Pk�= 4@��ܚ��!?�3�E)��@U�ۦ\�ٿ���F���@&	�2 4@.Q�ǐ!?�QI)��@���L�ٿ���P���@i�B� 4@�f�!?Y�C)��@���L�ٿ���P���@i�B� 4@�f�!?Y�C)��@gL�9�ٿ	�JW���@���C 4@~�kYg�!?�T�A)��@���-�ٿ2��_���@��N 4@	�Ev�!?O@)��@����ٿ��n���@�b�� 4@Oٜ�[�!?�$d@)��@K[�Y�ٿ�C�p���@C��s 4@��v��!?@�:)��@Ro8'�ٿ��a���@��ʷ 4@&��Ӑ!?�I]?)��@����>�ٿ�H�V���@�i� 4@�$��E�!?�-�B)��@����>�ٿ�H�V���@�i� 4@�$��E�!?�-�B)��@f
v3�ٿ���^���@'��* 4@����!?���B)��@��;�ٿ���\���@P��& 4@|~P蘐!?��tF)��@5��;�ٿ�[���@f(c 4@W��<Ð!?���F)��@ ��C�ٿ."fV���@Y�`w 4@oj��Ґ!?�Q�G)��@�^K�ٿa��M���@���3 4@���	�!?h˷G)��@��rk6�ٿL��Y���@�[�n 4@�Xې!?�H)��@
d��=�ٿ5��[���@�#E� 4@�|���!?>w"I)��@�a�cA�ٿ�|�X���@��g 4@4̝�!?�UC)��@�a�cA�ٿ�|�X���@��g 4@4̝�!?�UC)��@3�אA�ٿX�Y���@
b)� 4@�]�b+�!?�=�E)��@�0ok-�ٿ�7
^���@En�� 4@)R�'�!?�E)��@6�1�ٿ�f_���@b�f" 4@	ۼ�!?�Q�A)��@����D�ٿ���V���@L�8B 4@�����!?cR�E)��@����D�ٿ���V���@L�8B 4@�����!?cR�E)��@<���F�ٿVc}U���@,��E 4@��3e�!?1�D)��@đ|zQ�ٿ�$ P���@EP�� 4@y���̐!?�?G)��@đ|zQ�ٿ�$ P���@EP�� 4@y���̐!?�?G)��@Ɠx�J�ٿ���S���@;�bv 4@8�!?��H)��@Ɠx�J�ٿ���S���@;�bv 4@8�!?��H)��@�$mP�ٿ�s�P���@��*� 4@�==/��!?�AH)��@�$`�ٿfêK���@W�k 4@��>翐!?;1bJ)��@�⾲p�ٿ��<���@B��v 4@R�֐!?��)N)��@rZ��u�ٿq��;���@H�Zn 4@��5���!?���S)��@�D�~�ٿ<�4���@�5�� 4@�x3��!?;=�V)��@�D�~�ٿ<�4���@�5�� 4@�x3��!?;=�V)��@�G�"��ٿ�0R8���@�Y�� 4@��*�!?�Z)��@�{Mg��ٿb��-���@�.~	 4@B_�� �!?���^)��@�{Mg��ٿb��-���@�.~	 4@B_�� �!?���^)��@�{Mg��ٿb��-���@�.~	 4@B_�� �!?���^)��@%�K���ٿ�6P.���@��X 4@���c��!?��^\)��@��{D��ٿE	$ ���@�W�@ 4@Hh9��!?Sc)��@R��B��ٿ3��(���@!�x9 4@VJ��3�!?��L[)��@ C�V��ٿ������@�@�
 4@uÈ�-�!?�e)��@��馃�ٿ�m{3���@!U�Q 4@/=��(�!?�&v[)��@�T�Z��ٿƧq6���@!�Ư 4@K�ĺ/�!?�nY)��@���e��ٿX_)���@g�]� 4@��:*�!?��a)��@���߈�ٿ�7l2���@7��` 4@��f0ɐ!?�CQX)��@A�7��ٿe#�0���@
wD 4@���ޤ�!?Jt])��@2x���ٿ��5���@%Z 4@TxZ��!?z\X])��@2x���ٿ��5���@%Z 4@TxZ��!?z\X])��@�y��h�ٿ!�UB���@��4� 4@��zΪ�!?�#�P)��@n��n��ٿ���1���@g�?` 4@�S��!?��W)��@��K/��ٿ�L/!���@ν�q 4@��)���!?��])��@��K/��ٿ�L/!���@ν�q 4@��)���!?��])��@=74?��ٿ wO���@��K 4@f3��!?+3=^)��@-�b�c�ٿ�cGK���@zF 4@>����!?u?;I)��@-�b�c�ٿ�cGK���@zF 4@>����!?u?;I)��@�g�d��ٿ�1;���@5N*) 4@o ��|�!?W'�W)��@�dmȮ�ٿ&�,���@�rG8 4@*��ɭ�!?�_ZZ)��@�dmȮ�ٿ&�,���@�rG8 4@*��ɭ�!?�_ZZ)��@�z����ٿ��9���@:>�� 4@kwhݐ!?�X�T)��@�츣�ٿt��5���@�w�� 4@�t蕐!?�W)��@�츣�ٿt��5���@�w�� 4@�t蕐!?�W)��@*��˚ٿ�M!���@�� 4@�F�⍐!?�?�`)��@*��˚ٿ�M!���@�� 4@�F�⍐!?�?�`)��@�f:��ٿ��.(���@T9� 4@�
���!?߳O\)��@Pi����ٿ�1�6���@�4�� 4@}���!?]R�Y)��@$D���ٿ�C?2���@�8�� 4@�o�Q�!?]�^)��@$D���ٿ�C?2���@�8�� 4@�o�Q�!?]�^)��@���ɢ�ٿ�C�1���@���v 4@;N�I�!?R#�])��@���ɢ�ٿ�C�1���@���v 4@;N�I�!?R#�])��@���ɢ�ٿ�C�1���@���v 4@;N�I�!?R#�])��@�y�Uy�ٿ9�G���@vg= 4@�N���!?��T)��@�����ٿ3��7���@��K� 4@=�U��!?��n`)��@��(*�ٿ�ZU����@��s� 4@��-א!?�2�y)��@*�0�ٿk'W����@�9E� 4@�n�{�!?Q$��)��@*�0�ٿk'W����@�9E� 4@�n�{�!?Q$��)��@*�0�ٿk'W����@�9E� 4@�n�{�!?Q$��)��@Е�ߚٿ�����@�f � 4@2�M��!?㖉p)��@����ٿ T<���@a�� 4@!�bd��!?u��o)��@�E�3�ٿ[������@�;� 4@�}�5r�!?����)��@�� D��ٿ������@Ce� 4@ι�H��!?�b~v)��@��օ��ٿX������@B� 4@F�U!?���v)��@��օ��ٿX������@B� 4@F�U!?���v)��@��օ��ٿX������@B� 4@F�U!?���v)��@��օ��ٿX������@B� 4@F�U!?���v)��@��օ��ٿX������@B� 4@F�U!?���v)��@br����ٿM-e2���@SU	 4@��c�u�!?f�])��@'���ٿ?_���@p\Q' 4@�Vo�ǐ!?��Dv)��@'���ٿ?_���@p\Q' 4@�Vo�ǐ!?��Dv)��@��0��ٿ�=2���@=T� 4@6��R��!?���[)��@QF��ٿR�����@|��� 4@@�^9��!?��<{)��@����ٿ������@�6�� 4@W����!?����)��@����ٿ������@�6�� 4@W����!?����)��@����ٿ������@�6�� 4@W����!?����)��@����ٿ������@�6�� 4@W����!?����)��@�-�9��ٿ�(���@�7# 4@�Bil��!?��b)��@�T��a�ٿ
a4E���@yb 4@��5P��!?⫰S)��@i<ſ��ٿN�h.���@9�T 4@C��:{�!?�*h\)��@i<ſ��ٿN�h.���@9�T 4@C��:{�!?�*h\)��@i<ſ��ٿN�h.���@9�T 4@C��:{�!?�*h\)��@i<ſ��ٿN�h.���@9�T 4@C��:{�!?�*h\)��@�L�Ěٿ��,���@�f� 4@J�XY�!?�mq)��@z<-���ٿ9c����@m��g 4@R�_a�!?�HUp)��@������ٿ��f)���@��� 4@�,Y-ې!?�<�Z)��@����W�ٿ��G���@�U# 4@����!?T٦R)��@�:�Ds�ٿHΐ8���@H� 4@8K?��!?��])��@�>��ٿ�+���@���� 4@�]}��!?W�)a)��@P��q��ٿ�'���@�Kxa 4@ �%�!?o��q)��@P��q��ٿ�'���@�Kxa 4@ �%�!?o��q)��@�^t���ٿ�S�&���@�f� 4@C�g"�!?{l�d)��@^���N�ٿ��L���@�5�� 4@�ر�֐!?!i�N)��@�+D���ٿeq�-���@L�n 4@�����!?Oc)��@�,�|Z�ٿ��@���@���<	 4@��p�y�!?��s])��@�S/)�ٿe/q���@O�@� 4@��~敖!?" E)��@��4O�ٿ��O���@�\2� 4@\���!?R�R)��@�>̐�ٿ؎�+���@��" 4@��݁�!?�h)��@C�O���ٿ�6�8���@�7 4@�Mg�J�!?z�]k)��@l	��]�ٿw	N���@5��4 4@�t5t�!?��Z)��@�m�S�ٿ��z	���@ ��� 4@���!�!?��؇)��@�m�S�ٿ��z	���@ ��� 4@���!�!?��؇)��@�m�S�ٿ��z	���@ ��� 4@���!�!?��؇)��@ 9N�ٿ������@�8!� 4@4[�;7�!?��l�)��@�EMQ�ٿ�4����@�{�� 4@"�j�ΐ!?N�)��@�EMQ�ٿ�4����@�{�� 4@"�j�ΐ!?N�)��@�EMQ�ٿ�4����@�{�� 4@"�j�ΐ!?N�)��@����ٿ%������@�<Rg 4@�����!?��>�)��@o ����ٿX_���@�N�  4@�Y�#�!?��[�)��@o ����ٿX_���@�N�  4@�Y�#�!?��[�)��@o ����ٿX_���@�N�  4@�Y�#�!?��[�)��@o ����ٿX_���@�N�  4@�Y�#�!?��[�)��@z}�d�ٿ��)A���@?�n 4@���6�!?y��p)��@�:c�`�ٿ�p8���@���u��3@���֐!?]�v)��@�:c�`�ٿ�p8���@���u��3@���֐!?]�v)��@��D7ԙٿ��~���@Ȳ�: 4@�6����!?qD�()��@��D7ԙٿ��~���@Ȳ�: 4@�6����!?qD�()��@{0j-��ٿ��ߑ���@r�� 4@	��h�!?9��)��@{0j-��ٿ��ߑ���@r�� 4@	��h�!?9��)��@����ۙٿ<Jz���@��
 4@e�$~�!?�ɏ<)��@��d8�ٿ�^Q���@r�	 4@�Bjɐ!?8�T)��@�j����ٿ�[����@��� 4@v �n��!?Z9m)��@�j����ٿ�[����@��� 4@v �n��!?Z9m)��@�j����ٿ�[����@��� 4@v �n��!?Z9m)��@:����ٿ�G����@�" 4@�/�I̐!?6�o�)��@:����ٿ�G����@�" 4@�/�I̐!?6�o�)��@�r#��ٿ��pV���@�����3@��]�֐!?�Q*��@�r#��ٿ��pV���@�����3@��]�֐!?�Q*��@��h��ٿ�������@k)�  4@����Y�!? ��)��@5cq�-�ٿ������@��v 4@=K�}�!?5��)��@g����ٿш�����@��W 4@����y�!?9~A�)��@�AS\a�ٿ|�����@���. 4@	��酐!?�� )��@�AS\a�ٿ|�����@���. 4@	��酐!?�� )��@�AS\a�ٿ|�����@���. 4@	��酐!?�� )��@Q�_�]�ٿ�����@�]�� 4@ �I���!?�ǯ)��@���'�ٿע. ��@|��X 4@�%���!?�2�(��@E�ؘٿS�����@��X 4@����x�!?����(��@X���ٿ��҈���@�c*Z 4@q2N賐!?�$)��@ {��ٿf����@�B� 4@�O]���!?�N��)��@�^��ٿ�3�#���@GT. 4@JH/*��!?Z�ze)��@�lҫ�ٿ�!���@ "R	 4@�Q|��!?K8j})��@�lҫ�ٿ�!���@ "R	 4@�Q|��!?K8j})��@�Xq�_�ٿ��s����@��� 4@�"���!?�έ)��@�Xq�_�ٿ��s����@��� 4@�"���!?�έ)��@�2GT�ٿ��y���@VQ�B
 4@՟��!?
�R�)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@(��ٿ��C{���@p �^ 4@����!?�K��)��@�\\	�ٿ�
���@���\ 4@��B`�!?��R�)��@����ٿ4�71���@��� 4@�>�_h�!?%�?n)��@����ٿ4�71���@��� 4@�>�_h�!?%�?n)��@s�}�ٿN�	����@�� 4@�Y����!?�i�)��@s�}�ٿN�	����@�� 4@�Y����!?�i�)��@s�}�ٿN�	����@�� 4@�Y����!?�i�)��@���P0�ٿ�����@so'��3@yy3���!?��G�)��@���P0�ٿ�����@so'��3@yy3���!?��G�)��@���P0�ٿ�����@so'��3@yy3���!?��G�)��@�����ٿF��0���@0�z 4@���Ð!?t��})��@�X:F�ٿ۸#x���@ߩ·��3@e>;M��!?��*c)��@}Q]ԯ�ٿ������@�����3@3�,��!?4�@�)��@}Q]ԯ�ٿ������@�����3@3�,��!?4�@�)��@F����ٿN{�R���@���Y��3@�)�hא!?apf&*��@F����ٿN{�R���@���Y��3@�)�hא!?apf&*��@^�����ٿO����@;�B{��3@՝dխ�!?�b��*��@�H㠃�ٿ�G�����@<t��3@����!?`\^�+��@I>s�
�ٿs��y���@�����3@}L����!?��m,��@I>s�
�ٿs��y���@�����3@}L����!?��m,��@���ݥٿ���'���@ʿf��3@F��S��!?C���,��@1�>#��ٿ�����@�����3@�����!?��	,��@1�>#��ٿ�����@�����3@�����!?��	,��@����ٿ�kn���@�h3-��3@c�(��!?�=ņ*��@��+��ٿLԸ���@�'Z��3@�x�N�!?&�(;,��@��+��ٿLԸ���@�'Z��3@�x�N�!?&�(;,��@��PS��ٿ� ����@0Al�{�3@MR��!?)���,��@���9��ٿ�
����@oI�^��3@��q��!?��{,��@�����ٿ�v���@�>u���3@/�R���!?O��,��@�����ٿ�v���@�>u���3@/�R���!?O��,��@�����ٿ�v���@�>u���3@/�R���!?O��,��@�����ٿ�v���@�>u���3@/�R���!?O��,��@��k��ٿ�-Λ���@ɮ����3@�bȰq�!?򺜓+��@��k��ٿ�-Λ���@ɮ����3@�bȰq�!?򺜓+��@4*�*�ٿg��
���@��oS��3@-?�_��!?��/i*��@ć~:m�ٿӊ�"���@���O��3@ %ѐ!?�i�+��@ć~:m�ٿӊ�"���@���O��3@ %ѐ!?�i�+��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@�#�5��ٿ\������@�%P�m�3@~jM��!?7K{-��@J�i��ٿK�����@�H�} 4@a2䦫�!?,�<�(��@,Ԟ��ٿ��4���@�^?E��3@�b�as�!?oFvB+��@,Ԟ��ٿ��4���@�^?E��3@�b�as�!?oFvB+��@,Ԟ��ٿ��4���@�^?E��3@�b�as�!?oFvB+��@�#����ٿG}�����@3=��3@L����!?��-��@r��p�ٿ�i�����@��  4@Ϥ�}�!?�a/4*��@r��p�ٿ�i�����@��  4@Ϥ�}�!?�a/4*��@r��p�ٿ�i�����@��  4@Ϥ�}�!?�a/4*��@r��p�ٿ�i�����@��  4@Ϥ�}�!?�a/4*��@�n���ٿɷx����@HenA��3@Y����!?6�p�,��@�n���ٿɷx����@HenA��3@Y����!?6�p�,��@�n���ٿɷx����@HenA��3@Y����!?6�p�,��@���= �ٿ�%���@�`E?��3@� 5U��!?�eyu,��@»�ԢٿK������@=�h%w�3@���0ڐ!?��^,��@:��x�ٿE�`���@�8(#��3@��8h�!?���+��@�6�-�ٿq;�����@�Q;��3@�6�x�!?{��+��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@�x ��ٿ�w�����@:"���3@����4�!?��p�*��@��Y�D�ٿ�P����@�V���3@�螟,�!?@$�+��@��Y�D�ٿ�P����@�V���3@�螟,�!?@$�+��@!�{\�ٿ�������@v�ǫ�3@:���m�!?�E�i+��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@'��e�ٿq��m���@v�e�3@ʜ?��!?օ��,��@����ٿ�������@�0X�k�3@�Cv�!?�4#0+��@�/�ߟ�ٿ
�t���@R���3@�KU�ʐ!?�Ց.��@ZC)�ͨٿ���(���@�@m���3@��O�!?�3��-��@ZC)�ͨٿ���(���@�@m���3@��O�!?�3��-��@ZC)�ͨٿ���(���@�@m���3@��O�!?�3��-��@ZC)�ͨٿ���(���@�@m���3@��O�!?�3��-��@v��#�ٿXBi ��@�����3@���";�!?k��2)��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@�xX��ٿ��v���@��3K#�3@-@�v�!?}j[.��@ Q��ٿs/o���@����3@�Er�/�!?Q6�x-��@�
jM�ٿ�Jv��@O�4 4@3�U�!?$WX�'��@��ZМٿC[rr���@F�ڂ��3@���3V�!?R|��)��@'�E�Ϥٿu�T���@t�y�=�3@�C�$�!?�pz,��@'�E�Ϥٿu�T���@t�y�=�3@�C�$�!?�pz,��@'�E�Ϥٿu�T���@t�y�=�3@�C�$�!?�pz,��@�����ٿ���7 ��@HdNs 4@ъ�U��!?/4ѽ(��@�pr'ߜٿ�59����@��g�y�3@X���ː!?tZ��*��@�pr'ߜٿ�59����@��g�y�3@X���ː!?tZ��*��@���ٿ�)���@h�B�(�3@�])�Ր!?����,��@��B�^�ٿ(K�Z���@��GNe�3@lP��q�!?h�L�+��@��B�^�ٿ(K�Z���@��GNe�3@lP��q�!?h�L�+��@o��0�ٿ�Vm.���@+<K��3@|�rw�!?�m��*��@o��0�ٿ�Vm.���@+<K��3@|�rw�!?�m��*��@>�I7��ٿ���U���@:c�lB�3@{SV�!?.~�+��@>�I7��ٿ���U���@:c�lB�3@{SV�!?.~�+��@>�I7��ٿ���U���@:c�lB�3@{SV�!?.~�+��@���`�ٿ,jۮ���@.@V;�3@2���!?����+��@���`�ٿ,jۮ���@.@V;�3@2���!?����+��@���`�ٿ,jۮ���@.@V;�3@2���!?����+��@���`�ٿ,jۮ���@.@V;�3@2���!?����+��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@s8'9ġٿ��
���@�n���3@?WU��!?\�2�,��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@)B�p�ٿ�����@�V/�3@g�א!?+�4.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@_����ٿ*a�*���@l4a��3@�i�ݗ�!?/�|T.��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@)PѴ^�ٿ��`����@cQ�d�3@p�����!?}�"�+��@�@���ٿ%Q�����@� $A4@{�Ȑ!?N��(��@�@���ٿ%Q�����@� $A4@{�Ȑ!?N��(��@�@���ٿ%Q�����@� $A4@{�Ȑ!?N��(��@�ou��ٿ��&���@�m�2"4@�O����!? Ly�(��@|D�2��ٿ��4D���@#���3@}%� А!?M�]�-��@t�H�ٿHh|���@M�g��3@�*��!?~�v;1��@t�H�ٿHh|���@M�g��3@�*��!?~�v;1��@t�H�ٿHh|���@M�g��3@�*��!?~�v;1��@t�H�ٿHh|���@M�g��3@�*��!?~�v;1��@t�H�ٿHh|���@M�g��3@�*��!?~�v;1��@a50,�ٿgb�����@ف�[�3@RpJ��!?����0��@a50,�ٿgb�����@ف�[�3@RpJ��!?����0��@ ��&(�ٿ��\���@^�;�L�3@x)D,ː!?����3��@����ٿ�2̮���@v,�q��3@������!?�NR�9��@����ٿ�2̮���@v,�q��3@������!?�NR�9��@Z�YA��ٿ�t�����@ �����3@m�D��!?'S��1��@�%B�~�ٿ��q���@���O��3@�U�xܐ!?|B1��@�%B�~�ٿ��q���@���O��3@�U�xܐ!?|B1��@�>�h�ٿJwa����@�KLB�3@lOA�ِ!?����:��@�>�h�ٿJwa����@�KLB�3@lOA�ِ!?����:��@�>�h�ٿJwa����@�KLB�3@lOA�ِ!?����:��@�>�h�ٿJwa����@�KLB�3@lOA�ِ!?����:��@D�~�z�ٿk�����@��֎��3@��Vɐ!?A�GR0��@�x+|�ٿu(����@�WTw��3@g�:���!?�ӗA��@���@�ٿًQ)���@m��Ӭ�3@�����!?�:'N��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�aF-��ٿǔ����@v�����3@�e����!?��@U��@�����ٿP�s����@]�j"�3@�ۑNʐ!?��QeQ��@�����ٿP�s����@]�j"�3@�ۑNʐ!?��QeQ��@�����ٿP�s����@]�j"�3@�ۑNʐ!?��QeQ��@�����ٿP�s����@]�j"�3@�ۑNʐ!?��QeQ��@�����ٿP�s����@]�j"�3@�ۑNʐ!?��QeQ��@�=1l�ٿD͔v���@V`a�c�3@�)�߸�!?�w�=��@��-�ٿ�#O����@�Vo�3@��瘐!?�[ŀ:��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@-K�b+�ٿ:�����@��c�3@�/�!?j���<��@'��y�ٿ�y���@�_-�3@��%ű�!?[w�?��@'��y�ٿ�y���@�_-�3@��%ű�!?[w�?��@'��y�ٿ�y���@�_-�3@��%ű�!?[w�?��@'��y�ٿ�y���@�_-�3@��%ű�!?[w�?��@'��y�ٿ�y���@�_-�3@��%ű�!?[w�?��@8� :��ٿ�������@jf_�3@z�E�א!?T�VL��@8� :��ٿ�������@jf_�3@z�E�א!?T�VL��@8� :��ٿ�������@jf_�3@z�E�א!?T�VL��@�q+���ٿ���� ��@.��>E�3@�mh�!?Eً`@��@�q+���ٿ���� ��@.��>E�3@�mh�!?Eً`@��@�q+���ٿ���� ��@.��>E�3@�mh�!?Eً`@��@eR*�T�ٿ��� ��@�l����3@u��L�!?!��Q��@eR*�T�ٿ��� ��@�l����3@u��L�!?!��Q��@eR*�T�ٿ��� ��@�l����3@u��L�!?!��Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@��aJ�ٿ��%$ ��@� t�K�3@�zWd�!?��c?Q��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@P�+-�ٿ��Qw��@$3N[�3@�JԐ!?|�4!E��@���T�ٿ��1� ��@��~�W�3@ނn��!?n8�E��@���T�ٿ��1� ��@��~�W�3@ނn��!?n8�E��@tvU.U�ٿ�<A� ��@�V���3@z�A!Ӑ!?.���B��@tvU.U�ٿ�<A� ��@�V���3@z�A!Ӑ!?.���B��@tvU.U�ٿ�<A� ��@�V���3@z�A!Ӑ!?.���B��@tvU.U�ٿ�<A� ��@�V���3@z�A!Ӑ!?.���B��@tvU.U�ٿ�<A� ��@�V���3@z�A!Ӑ!?.���B��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@o��ơٿ��9$��@�;�P�3@AvƊ�!?�{�E��@ �]{�ٿ���
��@�u���3@�3+���!?��U|H��@ �]{�ٿ���
��@�u���3@�3+���!?��U|H��@ �]{�ٿ���
��@�u���3@�3+���!?��U|H��@ �]{�ٿ���
��@�u���3@�3+���!?��U|H��@ �]{�ٿ���
��@�u���3@�3+���!?��U|H��@���<�ٿ�Ք�
��@�@(���3@�n��!?�֩�3��@���<�ٿ�Ք�
��@�@(���3@�n��!?�֩�3��@��yܠٿ�H���@���3@��z!?���<��@t^$o	�ٿ Yl/!��@�]���3@�\��!?N��8��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@_7�`�ٿ+�T<.��@�-��=�3@H{���!?�6wH+��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@[@8ֺ�ٿ���H��@�=��3@��3ن�!?���"��@�����ٿ�����@��~�3@������!?��@l���@�����ٿ�����@��~�3@������!?��@l���@/f\lr�ٿ_�.{��@�Ͽj��3@��<��!?0�V���@/f\lr�ٿ_�.{��@�Ͽj��3@��<��!?0�V���@�f���ٿ���u��@UW��3@�z(hi�!?"�P���@��T�0�ٿ�����@���	h�3@Tԣ}�!?�넡Z��@��T�0�ٿ�����@���	h�3@Tԣ}�!?�넡Z��@��T�0�ٿ�����@���	h�3@Tԣ}�!?�넡Z��@�ş�ٿ�6�]r��@|�=*��3@2��̇�!?�w#��@ݤוٿ��Eb��@eZ�� �3@'�r���!?�,��@�Y?4�ٿL�R��@�Y)'w�3@=�`ʐ!?Wp[9��@�Y?4�ٿL�R��@�Y)'w�3@=�`ʐ!?Wp[9��@�Y?4�ٿL�R��@�Y)'w�3@=�`ʐ!?Wp[9��@����ٿm�2��@'�����3@�Ϟcx�!?������@��ǣٿ��\�-��@��F��3@�7��!?\�	.��@*����ٿ:�!���@����3@�X���!?3P!��@*����ٿ:�!���@����3@�X���!?3P!��@*����ٿ:�!���@����3@�X���!?3P!��@*����ٿ:�!���@����3@�X���!?3P!��@*����ٿ:�!���@����3@�X���!?3P!��@*����ٿ:�!���@����3@�X���!?3P!��@U�O�&�ٿ��Z���@ƈ4m��3@f���!?�r�t��@U�O�&�ٿ��Z���@ƈ4m��3@f���!?�r�t��@U�O�&�ٿ��Z���@ƈ4m��3@f���!?�r�t��@�;����ٿl�C$���@k����3@7*if�!?�O�Ղ��@�;����ٿl�C$���@k����3@7*if�!?�O�Ղ��@�;����ٿl�C$���@k����3@7*if�!?�O�Ղ��@��찾�ٿ)�����@��}���3@�A�x̐!?e��D��@��찾�ٿ)�����@��}���3@�A�x̐!?e��D��@��찾�ٿ)�����@��}���3@�A�x̐!?e��D��@��찾�ٿ)�����@��}���3@�A�x̐!?e��D��@S�����ٿ.?�����@�8Tt�3@2����!?�q��d��@�u$�F�ٿ�� �T��@�Z�M�3@mɐ!?I��!��@�u$�F�ٿ�� �T��@�Z�M�3@mɐ!?I��!��@�u$�F�ٿ�� �T��@�Z�M�3@mɐ!?I��!��@�u$�F�ٿ�� �T��@�Z�M�3@mɐ!?I��!��@�u$�F�ٿ�� �T��@�Z�M�3@mɐ!?I��!��@N�m��ٿd����@�4��3@��:$�!?��"����@�����ٿ+Bݹ<��@�����3@�+C���!?p�fk4��@�����ٿ+Bݹ<��@�����3@�+C���!?p�fk4��@	�rm�ٿ��)X��@�����3@߭� �!?��ju��@	!����ٿ�`堉�@��a��3@\X�͐!?[E�C��@	!����ٿ�`堉�@��a��3@\X�͐!?[E�C��@	!����ٿ�`堉�@��a��3@\X�͐!?[E�C��@	!����ٿ�`堉�@��a��3@\X�͐!?[E�C��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@J+�ٿ��ɑ��@s\7�3@�xP5h�!?��V��@S#1|�ٿl?�%��@�"a��3@���W
�!?  h���@-�Wf��ٿ�����@ڐS���3@�D�`�!?� F��@߇>�ٿ�ܫg��@���$��3@'B=:͐!?�¤���@߇>�ٿ�ܫg��@���$��3@'B=:͐!?�¤���@F�bΗٿ;�=�3��@[��N�3@�{P	q�!?V�=���@�#��ٿ<��b���@g�GA~�3@�i��!?�4jb��@�APؘٿo�X��@~��
/�3@;G.%А!?:�4ݫ��@�APؘٿo�X��@~��
/�3@;G.%А!?:�4ݫ��@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@	<��ΝٿThM��@�[�m�3@ݽ��!?�����@u��K�ٿC��|��@e�I���3@��ۿ�!?�w�!���@6��}�ٿ���H���@H����3@(���x�!?�ͯp��@6��}�ٿ���H���@H����3@(���x�!?�ͯp��@6��}�ٿ���H���@H����3@(���x�!?�ͯp��@6��}�ٿ���H���@H����3@(���x�!?�ͯp��@6��}�ٿ���H���@H����3@(���x�!?�ͯp��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@q(X%��ٿ������@���A�3@5sl�!?O�<2��@���LC�ٿ&Q3���@�Dw�3@.Q���!?�̮���@���LC�ٿ&Q3���@�Dw�3@.Q���!?�̮���@���LC�ٿ&Q3���@�Dw�3@.Q���!?�̮���@怓n�ٿoS#�%��@9I�[�3@�Z#��!?Vl����@怓n�ٿoS#�%��@9I�[�3@�Z#��!?Vl����@怓n�ٿoS#�%��@9I�[�3@�Z#��!?Vl����@#�C!�ٿ"��@)��R��3@?L���!? �I_x��@���$�ٿ�iل��@
�g`�3@�y�!?�C���@���$�ٿ�iل��@
�g`�3@�y�!?�C���@z'��ٿ@�H��@`D��
�3@O����!?�LW����@=2a{N�ٿ����w��@�u�3@�8�G��!?����R��@���ٿޒ#ƻ��@RH�a@�3@GjB���!?�!ĉ��@���ٿޒ#ƻ��@RH�a@�3@GjB���!?�!ĉ��@���ٿޒ#ƻ��@RH�a@�3@GjB���!?�!ĉ��@�ٿ.�����@D�L���3@�0sn�!?��N?��@�ٿ.�����@D�L���3@�0sn�!?��N?��@��L��ٿd?����@�����3@��<�?�!?�2�]��@��L��ٿd?����@�����3@��<�?�!?�2�]��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@c��	i�ٿn{9��@�)�<��3@�����!?Y�y�)��@}����ٿ"]�9��@nKô�3@��[�l�!?�g�t��@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@n�st��ٿ
H��Ċ�@���	�3@!�H*�!?nKP���@��U���ٿ�A5��@r��ُ�3@�h9��!?�{k���@��U���ٿ�A5��@r��ُ�3@�h9��!?�{k���@��U���ٿ�A5��@r��ُ�3@�h9��!?�{k���@��U���ٿ�A5��@r��ُ�3@�h9��!?�{k���@��U���ٿ�A5��@r��ُ�3@�h9��!?�{k���@Z�G��ٿd�gdK��@"X���3@��(���!?��3�(��@Z�G��ٿd�gdK��@"X���3@��(���!?��3�(��@Z�G��ٿd�gdK��@"X���3@��(���!?��3�(��@U�ۜٿH�f3���@OP�� �3@��K�5�!?��9����@U�ۜٿH�f3���@OP�� �3@��K�5�!?��9����@U�ۜٿH�f3���@OP�� �3@��K�5�!?��9����@�Fj��ٿ��U���@���c�3@�z��֐!?+��#}��@�Fj��ٿ��U���@���c�3@�z��֐!?+��#}��@�Fj��ٿ��U���@���c�3@�z��֐!?+��#}��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@���6�ٿ	W����@^Yˮ-�3@���%��!?�݈� ��@v �9�ٿ�o�>"��@���s��3@]�B�!?�֏͙��@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@i:�/��ٿ	c%�@��@),?���3@X��Ԑ!?e��%���@*�j[�ٿ�?�Q��@�o�w��3@��^���!?E��4w��@*�j[�ٿ�?�Q��@�o�w��3@��^���!?E��4w��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@Y���ٿ������@p8HC��3@�ģ�!?���V��@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@�T�ݠٿhiMw���@���ϰ�3@y{cސ!?�kM����@U"ON�ٿ#���@ ŀ�^�3@$
8ϐ!?�9b���@U"ON�ٿ#���@ ŀ�^�3@$
8ϐ!?�9b���@U"ON�ٿ#���@ ŀ�^�3@$
8ϐ!?�9b���@U"ON�ٿ#���@ ŀ�^�3@$
8ϐ!?�9b���@U"ON�ٿ#���@ ŀ�^�3@$
8ϐ!?�9b���@�1�<�ٿ����u��@� ���3@�<�}�!?(�C���@b�S�ٿ�i򰊉�@�S���3@q�=`��!?�o?�`��@b�S�ٿ�i򰊉�@�S���3@q�=`��!?�o?�`��@b�S�ٿ�i򰊉�@�S���3@q�=`��!?�o?�`��@7��u�ٿ;F��;��@�dJ�3@̖m�Ґ!?�:��i��@7��u�ٿ;F��;��@�dJ�3@̖m�Ґ!?�:��i��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@Z��
g�ٿ,���)��@2l2�G�3@.m׼�!?���X��@��4�ٿD�M|t��@�[S��3@�~'wƐ!?V���@��4�ٿD�M|t��@�[S��3@�~'wƐ!?V���@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@!�PVi�ٿ�g!��@k��1�3@�A��!?�7��	��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@j��ly�ٿ"x�
U��@}7�o��3@�f�i�!?��y*��@NFV��ٿ�R�HJ��@�#����3@�kM��!?��,_��@!�vNǥٿ���>��@׬����3@��H��!?�6����@!�vNǥٿ���>��@׬����3@��H��!?�6����@!�vNǥٿ���>��@׬����3@��H��!?�6����@Hqo�-�ٿ��i�W��@T�V��3@x����!?i��~$��@Hqo�-�ٿ��i�W��@T�V��3@x����!?i��~$��@Hqo�-�ٿ��i�W��@T�V��3@x����!?i��~$��@Hqo�-�ٿ��i�W��@T�V��3@x����!?i��~$��@Hqo�-�ٿ��i�W��@T�V��3@x����!?i��~$��@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@ws�z��ٿ��ˈ��@֌��Y�3@��7��!?������@|��眝ٿ>
�\��@�jd�3@A�&��!?�&��:��@�^�hR�ٿ�uNl�@%7�4"�3@�,�Ɛ!?[�Y�G��@��` �ٿm ��o�@x|c��3@T�Or�!?6��I�@�,ٿ��x�@_�T"?�3@����!?�K�.1��@��qtɞٿ�x��f��@"�9�Z�3@�G0}��!?��8���@��qtɞٿ�x��f��@"�9�Z�3@�G0}��!?��8���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�20�d�ٿQ>GW���@k�B !�3@f��K��!?�&L���@�;�i�ٿW�+�F��@$uPd��3@�'�i�!?p.�����@�;�i�ٿW�+�F��@$uPd��3@�'�i�!?p.�����@�;�i�ٿW�+�F��@$uPd��3@�'�i�!?p.�����@�;�i�ٿW�+�F��@$uPd��3@�'�i�!?p.�����@�;�i�ٿW�+�F��@$uPd��3@�'�i�!?p.�����@w̜DԜٿ�~�&:��@�o���3@YX�ѣ�!?m��F��@��3�ٿ�n�	c��@Dv��(�3@�Ȟ%��!?��]���@��3�ٿ�n�	c��@Dv��(�3@�Ȟ%��!?��]���@��3�ٿ�n�	c��@Dv��(�3@�Ȟ%��!?��]���@C�祬�ٿ�,}q��@\�ǽ�3@ǐ���!?�c���@-h�%x�ٿ�$3��t�@}u��~�3@ʞmː!?<oI�� �@-h�%x�ٿ�$3��t�@}u��~�3@ʞmː!?<oI�� �@k�&KW�ٿN���d�@x��3@������!?�V%�	�@k�&KW�ٿN���d�@x��3@������!?�V%�	�@k�&KW�ٿN���d�@x��3@������!?�V%�	�@k�&KW�ٿN���d�@x��3@������!?�V%�	�@k�&KW�ٿN���d�@x��3@������!?�V%�	�@k�&KW�ٿN���d�@x��3@������!?�V%�	�@���R9�ٿ)�ʮ�n�@lIb_��3@m�wr�!?<q,0�@���R9�ٿ)�ʮ�n�@lIb_��3@m�wr�!?<q,0�@���R9�ٿ)�ʮ�n�@lIb_��3@m�wr�!?<q,0�@���R9�ٿ)�ʮ�n�@lIb_��3@m�wr�!?<q,0�@���R9�ٿ)�ʮ�n�@lIb_��3@m�wr�!?<q,0�@AԼ+r�ٿ��[���@����/�3@vV�V�!?�t�۝��@AԼ+r�ٿ��[���@����/�3@vV�V�!?�t�۝��@AԼ+r�ٿ��[���@����/�3@vV�V�!?�t�۝��@�i5�/�ٿ/9��l��@�7^�L�3@F¨���!?�ɞr��@�i5�/�ٿ/9��l��@�7^�L�3@F¨���!?�ɞr��@�m�ʟٿe�`��@���g�3@��B>ʐ!?j����@����ٿ�DX����@Ā�8�3@]�"�!?3�+���@����ٿ�DX����@Ā�8�3@]�"�!?3�+���@(b�ۙٿ.�Xʭ#�@��$��3@n{��!?���T��@���[��ٿ�Q��w��@�����3@��K�!?�� ����@D�aU0�ٿ�8�"���@x�C�
�3@�R�}ʐ!?�^��xb�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@˙�R�ٿpG����@�{�u�3@Iw�!?��<�-�@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�x��ٿ��E�E�@��.���3@�"�QL�!?��h���@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@�P%�Оٿ�(_�"�@y(Þ�3@����`�!?���':�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����A�ٿM��4.��@��>��3@c����!?��ã�@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@����v�ٿ@����@�P��.�3@8����!?VT����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@#��8�ٿuV�%���@���P��3@)Y$��!?̲����@�2R�ܜٿ`[�;t��@��2���3@5�h̐�!?؛�4~	�@�2R�ܜٿ`[�;t��@��2���3@5�h̐�!?؛�4~	�@�,p�~�ٿ �̫�W�@�����3@X��!?;b�=���@�,p�~�ٿ �̫�W�@�����3@X��!?;b�=���@�,p�~�ٿ �̫�W�@�����3@X��!?;b�=���@�,p�~�ٿ �̫�W�@�����3@X��!?;b�=���@H��!�ٿ@�;���@c<b���3@3�����!?�jw��@H��!�ٿ@�;���@c<b���3@3�����!?�jw��@H��!�ٿ@�;���@c<b���3@3�����!?�jw��@H��!�ٿ@�;���@c<b���3@3�����!?�jw��@H��!�ٿ@�;���@c<b���3@3�����!?�jw��@|X�L�ٿZ+�fv��@{�8��3@I�B���!?�2{
��@|X�L�ٿZ+�fv��@{�8��3@I�B���!?�2{
��@|X�L�ٿZ+�fv��@{�8��3@I�B���!?�2{
��@|X�L�ٿZ+�fv��@{�8��3@I�B���!?�2{
��@'#Og7�ٿ`��x��@���n�3@�Ȉ�ؐ!?�����@'#Og7�ٿ`��x��@���n�3@�Ȉ�ؐ!?�����@'#Og7�ٿ`��x��@���n�3@�Ȉ�ؐ!?�����@'#Og7�ٿ`��x��@���n�3@�Ȉ�ؐ!?�����@'#Og7�ٿ`��x��@���n�3@�Ȉ�ؐ!?�����@_��v�ٿ���X��@\��YN�3@�)񑛐!?��:"c��@_��v�ٿ���X��@\��YN�3@�)񑛐!?��:"c��@�=l���ٿf�=�1a�@TȦg�3@Z�t�!?2cM7�K�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�,w0@�ٿ���&�U�@����l�3@�dې!?$0n�LR�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@�"oV��ٿ1tlp��@�&,��3@ߛX�Ȑ!?.�hj�&�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@޳�[�ٿ����T�@"/����3@w�欐!?L�9S�@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@C�3X�ٿjQ��G��@���:�3@̖�dΐ!?��D ��@t��
i�ٿ"�w�s��@��ƥ�3@��en�!?��~Z��@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��R<�ٿ�.����@�6l��3@(�.ː!?,U���@��0�ܜٿsu��I�@d؆���3@8['Uː!?i(���@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@@�^��ٿ��Q��!�@��%�3@���4�!?�?$�p�@ތ ^)�ٿ~k�O,��@4�n���3@��A��!?��U���@ތ ^)�ٿ~k�O,��@4�n���3@��A��!?��U���@ތ ^)�ٿ~k�O,��@4�n���3@��A��!?��U���@ތ ^)�ٿ~k�O,��@4�n���3@��A��!?��U���@ތ ^)�ٿ~k�O,��@4�n���3@��A��!?��U���@������ٿ@|5Q��@�x���3@�Z�>�!?�{�'��@������ٿ@|5Q��@�x���3@�Z�>�!?�{�'��@����ٿY��'c��@�c�V2�3@�(�͐!?c���]+�@����ٿY��'c��@�c�V2�3@�(�͐!?c���]+�@�F�բٿ�l���@<ZXu��3@�F1ϐ!?���׬z�@�F�բٿ�l���@<ZXu��3@�F1ϐ!?���׬z�@��ٿxV�(-�@�<����3@�|�W��!?y�=L��@��ٿxV�(-�@�<����3@�|�W��!?y�=L��@��ٿxV�(-�@�<����3@�|�W��!?y�=L��@��ٿxV�(-�@�<����3@�|�W��!?y�=L��@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@yɔ�~�ٿ�i���@��"��3@�(H���!?�t9���@���kQ�ٿ�v��S��@5�i��3@�1>7�!?|fҜ��@���kQ�ٿ�v��S��@5�i��3@�1>7�!?|fҜ��@���kQ�ٿ�v��S��@5�i��3@�1>7�!?|fҜ��@���kQ�ٿ�v��S��@5�i��3@�1>7�!?|fҜ��@���kQ�ٿ�v��S��@5�i��3@�1>7�!?|fҜ��@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@�=$��ٿ�&=�!}�@@�P�3@n^�Ő!?>��&C;�@~�*ܰ�ٿ8}�N���@�WCm�3@�����!?�֤t���@~�*ܰ�ٿ8}�N���@�WCm�3@�����!?�֤t���@~�*ܰ�ٿ8}�N���@�WCm�3@�����!?�֤t���@~�*ܰ�ٿ8}�N���@�WCm�3@�����!?�֤t���@~�*ܰ�ٿ8}�N���@�WCm�3@�����!?�֤t���@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�r���ٿ��'~u��@��oؒ�3@߷n��!?y�/����@�B��ٿ!z�%�@ ?L���3@_��+�!?l��-��@o��9o�ٿ��{���@HI{�3@�W�ڐ!?n�\��@o��9o�ٿ��{���@HI{�3@�W�ڐ!?n�\��@o��9o�ٿ��{���@HI{�3@�W�ڐ!?n�\��@�B��)�ٿ`E&�Pk�@��^w�3@�M/�ݐ!?e���2��@�B��)�ٿ`E&�Pk�@��^w�3@�M/�ݐ!?e���2��@�B��)�ٿ`E&�Pk�@��^w�3@�M/�ݐ!?e���2��@�B��)�ٿ`E&�Pk�@��^w�3@�M/�ݐ!?e���2��@�B��)�ٿ`E&�Pk�@��^w�3@�M/�ݐ!?e���2��@-&hӤ�ٿ�J�Yv�@R����3@%?08�!?��*���@Ȍ���ٿ��reR�@�;Nd�3@�0��!?��)2FT�@Ȍ���ٿ��reR�@�;Nd�3@�0��!?��)2FT�@Ȍ���ٿ��reR�@�;Nd�3@�0��!?��)2FT�@Ȍ���ٿ��reR�@�;Nd�3@�0��!?��)2FT�@Ȍ���ٿ��reR�@�;Nd�3@�0��!?��)2FT�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@"���ٿ�K��e�@~$D�!�3@l�ly!�!?')ސ]I�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@�4 �@�ٿf���u�@�����3@-�&h̐!?�&
@�@k��?�ٿ��&��@�y��A�3@yavt�!?�Ñ 7��@k��?�ٿ��&��@�y��A�3@yavt�!?�Ñ 7��@G�*y��ٿ3c��	h�@; �e�3@t��!?\2)���@G�*y��ٿ3c��	h�@; �e�3@t��!?\2)���@)vǘ�ٿf=a ��@ڙ:R�3@1`I$�!?�k�O���@)vǘ�ٿf=a ��@ڙ:R�3@1`I$�!?�k�O���@��!П�ٿ��7�=��@�ln��3@��Z.�!?ſ�ev��@ղv�ٿ�
�����@�В�8�3@L� �!?�u�%;��@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@q�N�'�ٿ71�D�C�@���� �3@z7��!?_����\�@�	_�âٿ�ER��	�@e��C��3@�Hr�!?���~�@�	_�âٿ�ER��	�@e��C��3@�Hr�!?���~�@[��,��ٿk�D����@1���=�3@I��6��!?�c1���@[��,��ٿk�D����@1���=�3@I��6��!?�c1���@[��,��ٿk�D����@1���=�3@I��6��!?�c1���@#�m&�ٿf�^�1�@sW�.�3@�Uce��!?��wg�@#�m&�ٿf�^�1�@sW�.�3@�Uce��!?��wg�@#�m&�ٿf�^�1�@sW�.�3@�Uce��!?��wg�@� `$�ٿ��d�|�@B[(j�3@4����!?��k��;�@� `$�ٿ��d�|�@B[(j�3@4����!?��k��;�@� `$�ٿ��d�|�@B[(j�3@4����!?��k��;�@� `$�ٿ��d�|�@B[(j�3@4����!?��k��;�@Rd�~�ٿ4 z��h�@��><��3@����!?2o��G�@�����ٿM[>�߇�@�4��3@�����!?H�Pl��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@i%� �ٿJ��{S`�@�Op�3@���R��!? Y�+o��@�LR���ٿB���3a�@W�BG[�3@�th⬐!? ������@�LR���ٿB���3a�@W�BG[�3@�th⬐!? ������@�LR���ٿB���3a�@W�BG[�3@�th⬐!? ������@�LR���ٿB���3a�@W�BG[�3@�th⬐!? ������@���E1�ٿ��\&��@a�TN�3@!���!?- 1����@��(�s�ٿr�x"�@���%�3@�6
�!?��o2p�@��(�s�ٿr�x"�@���%�3@�6
�!?��o2p�@��(�s�ٿr�x"�@���%�3@�6
�!?��o2p�@�a��Z�ٿ����Č�@H	���3@�y@��!?*5�{��@�a��Z�ٿ����Č�@H	���3@�y@��!?*5�{��@�a��Z�ٿ����Č�@H	���3@�y@��!?*5�{��@�6o���ٿ�9+�-�@���D@�3@2vo�@�!?0��I~��@�6o���ٿ�9+�-�@���D@�3@2vo�@�!?0��I~��@�6o���ٿ�9+�-�@���D@�3@2vo�@�!?0��I~��@�6o���ٿ�9+�-�@���D@�3@2vo�@�!?0��I~��@�6o���ٿ�9+�-�@���D@�3@2vo�@�!?0��I~��@Z��H�ٿ��1R��@�9�9�3@
f(v�!?��~��7�@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@�0�E�ٿ'h��b�@V3�F��3@�R?"�!?/�����@� �:b�ٿv�O�R�@>�u>y�3@C`ߐ!?��0	�@]#��ʤٿ�3�=�d�@B�T�3@�x���!?���s���@]#��ʤٿ�3�=�d�@B�T�3@�x���!?���s���@]#��ʤٿ�3�=�d�@B�T�3@�x���!?���s���@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@Qɨנٿ ��;�G�@�̞��3@M�r��!?	�a����@���#�ٿ�֭��i�@x����3@�|����!?>u����@���#�ٿ�֭��i�@x����3@�|����!?>u����@���#�ٿ�֭��i�@x����3@�|����!?>u����@뷝��ٿ7��f�@4�'L�3@�bVj��!?��O��@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@������ٿ:3�m��@Hw�2G�3@R@r(��!?���-�0�@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@�yI^�ٿˌZ����@�P�3@��m��!?hN����@	D�@+�ٿ�i�Q8��@6�	�+�3@,v%��!?��k��@	D�@+�ٿ�i�Q8��@6�	�+�3@,v%��!?��k��@	D�@+�ٿ�i�Q8��@6�	�+�3@,v%��!?��k��@	D�@+�ٿ�i�Q8��@6�	�+�3@,v%��!?��k��@	D�@+�ٿ�i�Q8��@6�	�+�3@,v%��!?��k��@��d���ٿ�U����@��Р�3@��yׄ�!?	 �R��@��d���ٿ�U����@��Р�3@��yׄ�!?	 �R��@}}?[�ٿ#��h�@G=����3@߮昼�!?|��-�G�@�q�wr�ٿ��M:��@US��3@���e͐!?�i"/D��@�q�wr�ٿ��M:��@US��3@���e͐!?�i"/D��@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@d�2><�ٿ�E��@oŚ]��3@��CѮ�!?���+���@�u��ٿ�*��N��@��n��3@90�̐!?g\���@�� _��ٿ�(�FY�@ms9��3@����!?��F��@�� _��ٿ�(�FY�@ms9��3@����!?��F��@�� _��ٿ�(�FY�@ms9��3@����!?��F��@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@7nEj��ٿ|�!�(5�@YW�#��3@AGǍ��!?������@f'���ٿЙ}��@M4 C��3@J��s|�!?�ߥ-}�@f'���ٿЙ}��@M4 C��3@J��s|�!?�ߥ-}�@��H�ٿ�'�$��@�sq� 4@���_Ґ!?$�K�_��@��H�ٿ�'�$��@�sq� 4@���_Ґ!?$�K�_��@��H�ٿ�'�$��@�sq� 4@���_Ґ!?$�K�_��@��H�ٿ�'�$��@�sq� 4@���_Ґ!?$�K�_��@�^6�ٿ���87�@Dຖ�3@�M��!?#|��u��@�^6�ٿ���87�@Dຖ�3@�M��!?#|��u��@�^6�ٿ���87�@Dຖ�3@�M��!?#|��u��@?��8��ٿԵ����@L���3@ڗ蓐!?�2"���@�����ٿ���F�@2�kq�3@���l�!?c��f(\�@�����ٿ���F�@2�kq�3@���l�!?c��f(\�@�����ٿ���F�@2�kq�3@���l�!?c��f(\�@�����ٿ���F�@2�kq�3@���l�!?c��f(\�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@f��t�ٿ<��� �@ T��N�3@������!?���>zp�@U�1i��ٿzL�ſ��@�eIڱ�3@(�`���!?�g&U��@U�1i��ٿzL�ſ��@�eIڱ�3@(�`���!?�g&U��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�����ٿ�~"=z�@�uR��3@Q(�ɐ!?�Y�g��@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@�GA�ٿ]j�9j�@�����3@����s�!?T��kz�@����ʞٿ:ל}9K�@�@��3�3@�`����!?�v{yX�@����ʞٿ:ל}9K�@�@��3�3@�`����!?�v{yX�@�<���ٿ�]�P��@�ܼh��3@t
�0Ӑ!?�+HT�{�@�<���ٿ�]�P��@�ܼh��3@t
�0Ӑ!?�+HT�{�@�<���ٿ�]�P��@�ܼh��3@t
�0Ӑ!?�+HT�{�@�<���ٿ�]�P��@�ܼh��3@t
�0Ӑ!?�+HT�{�@�<���ٿ�]�P��@�ܼh��3@t
�0Ӑ!?�+HT�{�@��v��ٿꖐ��&�@P����3@��j��!?��W� �@��v��ٿꖐ��&�@P����3@��j��!?��W� �@��v��ٿꖐ��&�@P����3@��j��!?��W� �@��v��ٿꖐ��&�@P����3@��j��!?��W� �@��v��ٿꖐ��&�@P����3@��j��!?��W� �@��v��ٿꖐ��&�@P����3@��j��!?��W� �@�rr��ٿk����@��� 6�3@�6���!?b����	�@�rr��ٿk����@��� 6�3@�6���!?b����	�@�rr��ٿk����@��� 6�3@�6���!?b����	�@�rr��ٿk����@��� 6�3@�6���!?b����	�@Dmϐ�ٿ���m>�@&E�5&�3@�}�[�!?�5�����@Dmϐ�ٿ���m>�@&E�5&�3@�}�[�!?�5�����@�J^�j�ٿ%����@��uɸ�3@}�+���!?�O����@�J^�j�ٿ%����@��uɸ�3@}�+���!?�O����@�J^�j�ٿ%����@��uɸ�3@}�+���!?�O����@��v���ٿ�p7�x�@~��	�3@1�Z}��!?g��g�@��v���ٿ�p7�x�@~��	�3@1�Z}��!?g��g�@��v���ٿ�p7�x�@~��	�3@1�Z}��!?g��g�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@,!g�g�ٿ:di���@�y�3@�lJ[�!?/(c	".�@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@~�7F�ٿ^qSjSg�@ރ�̈́�3@�����!?�����@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@U
�Q��ٿ\M�~��@"�����3@0K���!?lG3d��@�~��ٿԇ�rE�@�NU	��3@<���!?�r����@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@.�^�ٿ�F�y���@@Q�3c�3@�s]�#�!?q�?A��@xܦ�Ρٿ��J� ��@�����3@��VK�!?�u�£��@xܦ�Ρٿ��J� ��@�����3@��VK�!?�u�£��@xܦ�Ρٿ��J� ��@�����3@��VK�!?�u�£��@x�7���ٿ��ø���@���R��3@f!��ʐ!?e|��@̽[�_�ٿ�)pM�@���'��3@{����!?�ǂ��s�@̽[�_�ٿ�)pM�@���'��3@{����!?�ǂ��s�@̽[�_�ٿ�)pM�@���'��3@{����!?�ǂ��s�@̽[�_�ٿ�)pM�@���'��3@{����!?�ǂ��s�@�Y�n�ٿ����@�c<Y��3@0q.�l�!?�Ċu?��@E.��ٿ8/�0z-�@V���3@Cﴘ�!?�S����@E.��ٿ8/�0z-�@V���3@Cﴘ�!?�S����@E.��ٿ8/�0z-�@V���3@Cﴘ�!?�S����@E.��ٿ8/�0z-�@V���3@Cﴘ�!?�S����@\��Wڝٿ9����@�59���3@��o�!?4��G(�@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@���ٿ�����@�EԝY�3@�F秐!?�J���@Bsnu�ٿ<��)H��@?���u�3@%�d���!?IA�}��@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@:��G�ٿ��B���@3��p��3@*V���!?`�ʚ���@��Y�ٿ�UHP��@�.7�4�3@ ١;��!?��!Mt�@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@&�t�֠ٿ�@w��@wm2>�3@���#��!?���o���@��fw��ٿ�GMj(�@�NJ^��3@F��T2�!?���sr�@��fw��ٿ�GMj(�@�NJ^��3@F��T2�!?���sr�@��fw��ٿ�GMj(�@�NJ^��3@F��T2�!?���sr�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@9�nߠٿ�c8aG��@��3���3@B����!?���s�.�@�Z�uC�ٿ[S�(BU�@�oh�)�3@��i�̐!?v$�0P�@�Z�uC�ٿ[S�(BU�@�oh�)�3@��i�̐!?v$�0P�@�Z�uC�ٿ[S�(BU�@�oh�)�3@��i�̐!?v$�0P�@�Z�uC�ٿ[S�(BU�@�oh�)�3@��i�̐!?v$�0P�@���wۜٿ+T�Df�@'�G] �3@�s��!?1"tF�@���wۜٿ+T�Df�@'�G] �3@�s��!?1"tF�@���wۜٿ+T�Df�@'�G] �3@�s��!?1"tF�@���wۜٿ+T�Df�@'�G] �3@�s��!?1"tF�@M0bI�ٿ�[�5b��@<>�Xu�3@�$�7��!?�7��5'�@�����ٿD���=�@F*
���3@r���!?Pv2�_�@������ٿL0g���@�ں�3@�OE�ِ!?��J���@������ٿL0g���@�ں�3@�OE�ِ!?��J���@������ٿL0g���@�ں�3@�OE�ِ!?��J���@������ٿL0g���@�ں�3@�OE�ِ!?��J���@������ٿL0g���@�ں�3@�OE�ِ!?��J���@���g�ٿK~��c�@�#u�-�3@���.�!?���t�P�@���g�ٿK~��c�@�#u�-�3@���.�!?���t�P�@�J���ٿxp��)�@�G���3@)�J���!?8�8(�t�@�J���ٿxp��)�@�G���3@)�J���!?8�8(�t�@�J���ٿxp��)�@�G���3@)�J���!?8�8(�t�@�J���ٿxp��)�@�G���3@)�J���!?8�8(�t�@\�R7]�ٿ���̥��@HmDQ�3@J��O��!?�
	ֿ�@\�R7]�ٿ���̥��@HmDQ�3@J��O��!?�
	ֿ�@\�R7]�ٿ���̥��@HmDQ�3@J��O��!?�
	ֿ�@�}ݵ]�ٿ�-�©{�@`#�G�3@.�����!?I^$S���@�}ݵ]�ٿ�-�©{�@`#�G�3@.�����!?I^$S���@�}ݵ]�ٿ�-�©{�@`#�G�3@.�����!?I^$S���@ȥP���ٿ�G�d%r�@n��d�3@ě�A�!?��>D�@��6Ð�ٿ2/j܄�@�����3@J=�@�!?�f����@�Ų���ٿ͐� �@����3@���!?�g?}�@�Ų���ٿ͐� �@����3@���!?�g?}�@�Ų���ٿ͐� �@����3@���!?�g?}�@�Ų���ٿ͐� �@����3@���!?�g?}�@ʅ?c��ٿ��Ȭw�@I&��3@YR�}��!?�Ns7�@�8�h�ٿ��7i��@8b�9��3@�Q�,Ԑ!?m(�6>��@�8�h�ٿ��7i��@8b�9��3@�Q�,Ԑ!?m(�6>��@�8�h�ٿ��7i��@8b�9��3@�Q�,Ԑ!?m(�6>��@�8�h�ٿ��7i��@8b�9��3@�Q�,Ԑ!?m(�6>��@�8�h�ٿ��7i��@8b�9��3@�Q�,Ԑ!?m(�6>��@��Sr��ٿ��I`]�@�}y��3@�IZ�!?sT*7�O�@�w>��ٿf�;V��@6u5q��3@�ݖ���!?x���@%#鏤ٿ�_� ��@m=�o|�3@sW���!?�.Z|� �@�mLUX�ٿ�-�ⱊ�@�����3@Waz!?G�C���@�mLUX�ٿ�-�ⱊ�@�����3@Waz!?G�C���@�mLUX�ٿ�-�ⱊ�@�����3@Waz!?G�C���@���=��ٿ�������@���<��3@�ȹ��!?�;����@�8��ٿ7�4յ��@�.8��3@�:��!?�d�y��@�8��ٿ7�4յ��@�.8��3@�:��!?�d�y��@��AJ�ٿ8���~��@��X���3@�7��֐!?�����@��AJ�ٿ8���~��@��X���3@�7��֐!?�����@��AJ�ٿ8���~��@��X���3@�7��֐!?�����@��AJ�ٿ8���~��@��X���3@�7��֐!?�����@L�U�o�ٿAG�A�y�@P0�r��3@֔��!?�����@L�U�o�ٿAG�A�y�@P0�r��3@֔��!?�����@L�U�o�ٿAG�A�y�@P0�r��3@֔��!?�����@L�U�o�ٿAG�A�y�@P0�r��3@֔��!?�����@L�U�o�ٿAG�A�y�@P0�r��3@֔��!?�����@;��ٿ����N�@��l���3@�>����!?��H\�@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@��#x�ٿ�
iz��@������3@�&���!?�L���@.v�P��ٿ/FsS��@�e���3@)>�ߌ�!?����5��@.v�P��ٿ/FsS��@�e���3@)>�ߌ�!?����5��@Qf�Ėٿӓ�����@���3@z�6��!?��%��@Qf�Ėٿӓ�����@���3@z�6��!?��%��@Qf�Ėٿӓ�����@���3@z�6��!?��%��@Qf�Ėٿӓ�����@���3@z�6��!?��%��@�-����ٿB����@��꼨�3@��rU�!?�:ᛋ�@�-����ٿB����@��꼨�3@��rU�!?�:ᛋ�@�-����ٿB����@��꼨�3@��rU�!?�:ᛋ�@�-����ٿB����@��꼨�3@��rU�!?�:ᛋ�@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@tヾڟٿ��	��@{oM8�3@���!?�F���@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@�� m�ٿEd���.�@|_3���3@������!?tQ<�n�@��̾�ٿ�>P��8�@`�R�3@�)��!?Z�~��]�@��̾�ٿ�>P��8�@`�R�3@�)��!?Z�~��]�@��̾�ٿ�>P��8�@`�R�3@�)��!?Z�~��]�@��̾�ٿ�>P��8�@`�R�3@�)��!?Z�~��]�@Wc�y�ٿS�Fa���@��D2�3@E�����!?���ņ��@Wc�y�ٿS�Fa���@��D2�3@E�����!?���ņ��@Wc�y�ٿS�Fa���@��D2�3@E�����!?���ņ��@Wc�y�ٿS�Fa���@��D2�3@E�����!?���ņ��@e�珞ٿ��[t���@L�A���3@��^gϐ!?޴���@�0�d�ٿ��k��@ߨH�_�3@�=Y�Ԑ!?�����@d|n��ٿ�H�C���@塨���3@��oZ��!?����,�@d|n��ٿ�H�C���@塨���3@��oZ��!?����,�@d|n��ٿ�H�C���@塨���3@��oZ��!?����,�@d|n��ٿ�H�C���@塨���3@��oZ��!?����,�@XC���ٿ���=n��@������3@����!?�^�;���@;�;�V�ٿ)9�����@g ��&�3@m�	�ݐ!?;��ƾ�@;�;�V�ٿ)9�����@g ��&�3@m�	�ݐ!?;��ƾ�@;�;�V�ٿ)9�����@g ��&�3@m�	�ݐ!?;��ƾ�@丅e�ٿ�:3_�]�@;)�3@����!?V,�2�M�@�I�/}�ٿO�����@��/��3@�'i��!?�n^���@�I�/}�ٿO�����@��/��3@�'i��!?�n^���@X����ٿqz�G�;�@jT���3@ŀ^#�!?+���Q�@X����ٿqz�G�;�@jT���3@ŀ^#�!?+���Q�@X����ٿqz�G�;�@jT���3@ŀ^#�!?+���Q�@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@EB�;�ٿw�Ob��@�$�B��3@��xސ!?%]'����@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@�a:�d�ٿ�#mm��@�kJ�3@k0����!?��O���@TpH2��ٿ�o;N��@��8�3@3��ˠ�!?Zٯ��@TpH2��ٿ�o;N��@��8�3@3��ˠ�!?Zٯ��@TpH2��ٿ�o;N��@��8�3@3��ˠ�!?Zٯ��@�����ٿ�X�ك��@�5��3@�.G쮐!?�^��Y��@gg)�ٿ��r���@��"�3@R8[���!?�Kg��@�%1�ٿ��:t b�@�c{R�3@D�����!?i[StAn�@�%1�ٿ��:t b�@�c{R�3@D�����!?i[StAn�@���ٿP���>�@�K0w4@�[M�ې!?�k����@���ٿP���>�@�K0w4@�[M�ې!?�k����@WO���ٿ�C�����@ل�3@%@�/ϐ!?�8;��@WO���ٿ�C�����@ل�3@%@�/ϐ!?�8;��@9�ڭ��ٿc�c`���@�
d�3@/�2��!?�?%����@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@��W�ٿ%�,6 �@���#�3@Ҁ�!?w��Ĕ��@#��E^�ٿ��*�]�@T/dQ�3@����!?�l]�9Y�@#��E^�ٿ��*�]�@T/dQ�3@����!?�l]�9Y�@�{US�ٿE;�1�'�@*�	
r�3@" ��!?9r"7�@�{US�ٿE;�1�'�@*�	
r�3@" ��!?9r"7�@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@܍ ٿ	�B5
��@Y\D��3@�1�ΐ!?'-�/��@z?��ٿ�{��P��@dѶ�4@��&�!?����n��@�B�N�ٿ�Gi�6+�@�~��F�3@Uܗò�!?q�?ŝ��@�B�N�ٿ�Gi�6+�@�~��F�3@Uܗò�!?q�?ŝ��@�B�N�ٿ�Gi�6+�@�~��F�3@Uܗò�!?q�?ŝ��@�B�N�ٿ�Gi�6+�@�~��F�3@Uܗò�!?q�?ŝ��@cؽ�d�ٿd�U�r�@�����3@ä	!ɐ!?�r�r7�@�3�E�ٿ��^���@n�h�3@ \u��!?�����@�3�E�ٿ��^���@n�h�3@ \u��!?�����@m�}sv�ٿ֕���@���3@8�U͚�!?f>���r�@m�}sv�ٿ֕���@���3@8�U͚�!?f>���r�@m�}sv�ٿ֕���@���3@8�U͚�!?f>���r�@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@�#1I�ٿ1,��1�@H����3@�~l3��!?�@YCf��@��P�ٿz��f�@��Bѹ�3@�饂�!?R<����@��P�ٿz��f�@��Bѹ�3@�饂�!?R<����@��P�ٿz��f�@��Bѹ�3@�饂�!?R<����@���0�ٿ��Ù4��@)�j}+ 4@Z�{�!?g暔`�@U8��ٿtY��&��@�X1Y�3@߈��ɐ!?�?���1�@U8��ٿtY��&��@�X1Y�3@߈��ɐ!?�?���1�@U8��ٿtY��&��@�X1Y�3@߈��ɐ!?�?���1�@U8��ٿtY��&��@�X1Y�3@߈��ɐ!?�?���1�@U8��ٿtY��&��@�X1Y�3@߈��ɐ!?�?���1�@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@��ԑ�ٿ��r&��@�c�� �3@�H��ΐ!?�,2�j��@?f��ٿ���5��@>�1<�3@�&D��!?�������@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@�Ï-�ٿ���ϭ��@��	~<�3@�oq�Ԑ!?����@���L�ٿR�����@}����3@��ߪ��!?�O�p
��@���L�ٿR�����@}����3@��ߪ��!?�O�p
��@O�@�ٿ�ܹ;v�@M�����3@?Ѡ�ܐ!?$\N����@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@mG��Ҩٿ��QG�@�- ќ�3@<�Y\�!?|�H��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@�0�
�ٿ��%����@4;;ӏ�3@u��!?c�<0&��@N�팢ٿ#��)��@+,�6�3@��0�Đ!?爫Ŭ��@}MJ���ٿC�>�(��@�I���3@p�A�ؐ!?')R#9�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@2n�=��ٿ��p�T��@S�t>t�3@!�~Ԑ!?ϊ �(8�@�I]ޘٿ4���}�@��p�3@�é���!?b��",+�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@`d�^��ٿ��O��@�L��3@v�M��!?��_Lwi�@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@���?W�ٿ�+2'��@�G�X��3@U;FB��!?MxY���@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@<G�Xj�ٿ�wJ�@e�o���3@*=eL��!?�?��+W�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�$��ٿ�="��@��.?!�3@���@ɐ!?)��r*�@�*\�1�ٿ/�](*��@
U�k��3@��d�ڐ!?5�K:��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@SY���ٿ�Ւ����@5/d{��3@��p��!?����{��@u�H+�ٿ�V����@�+��3@�|F67�!?S�P��@:?��ٿ ���Q�@��>�3@$��!?����0�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@E�n�v�ٿj,r�@T�����3@(��'�!?�Eg��>�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@�6ϊ��ٿ`����@/-����3@"��ͷ�!?(���|�@<v�Gèٿ�����@;����3@�2d���!?�--�
3�@�����ٿע�4A�@�'Zf��3@=��:ѐ!?ENU
���@L��U�ٿ��7d.��@�h�>�3@TR��!?�ln���@L��U�ٿ��7d.��@�h�>�3@TR��!?�ln���@L��U�ٿ��7d.��@�h�>�3@TR��!?�ln���@L��U�ٿ��7d.��@�h�>�3@TR��!?�ln���@�,�́�ٿ�}t����@B=�N��3@,����!?x�3���@�,�́�ٿ�}t����@B=�N��3@,����!?x�3���@�,�́�ٿ�}t����@B=�N��3@,����!?x�3���@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��� �ٿ��G]��@���t�3@߄�oȐ!?�J{y_�@��v���ٿ�V�t-��@�E]��3@6��b�!?�l
���@��v���ٿ�V�t-��@�E]��3@6��b�!?�l
���@��v���ٿ�V�t-��@�E]��3@6��b�!?�l
���@I�1�(�ٿ|��Ƭ�@���jH�3@C�(�!?�-�9r��@I�1�(�ٿ|��Ƭ�@���jH�3@C�(�!?�-�9r��@j���b�ٿdQ�Q0��@(�v+��3@�_U뜐!?}mC	��@j���b�ٿdQ�Q0��@(�v+��3@�_U뜐!?}mC	��@j���b�ٿdQ�Q0��@(�v+��3@�_U뜐!?}mC	��@��*$�ٿ8T��,�@/)�3@d��B�!?0�&W��@Fc�S�ٿ�1���@ ��1�3@���ڐ!?Z�Jx�h�@Fc�S�ٿ�1���@ ��1�3@���ڐ!?Z�Jx�h�@j��+�ٿ�x͋x�@�NQ��3@�m�ؐ!?�(+��@j��+�ٿ�x͋x�@�NQ��3@�m�ؐ!?�(+��@\����ٿ�n�����@b	+�x�3@vh���!?`v��u�@\����ٿ�n�����@b	+�x�3@vh���!?`v��u�@\����ٿ�n�����@b	+�x�3@vh���!?`v��u�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@��
4�ٿ���H��@¶�C��3@�����!?x�`��#�@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@�p�ٿ�G��͒�@����3@"t����!?������@��?>�ٿ�}���4�@�F�(�3@��<1��!?b�i+=s�@��?>�ٿ�}���4�@�F�(�3@��<1��!?b�i+=s�@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@�C�5�ٿ��l���@�l�W��3@ȁ�^��!?����@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@A����ٿ�����@�t���3@���8��!?�Ei!f�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@ ��uk�ٿ52�يm�@Oq
:��3@�y�wƐ!?���E�@���]�ٿ\��O�@p��jU�3@�#����!?<Dѹ68�@�qX,�ٿ"R�|���@~��R�3@f0]ˊ�!?*���9�@�qX,�ٿ"R�|���@~��R�3@f0]ˊ�!?*���9�@�qX,�ٿ"R�|���@~��R�3@f0]ˊ�!?*���9�@�qX,�ٿ"R�|���@~��R�3@f0]ˊ�!?*���9�@�qX,�ٿ"R�|���@~��R�3@f0]ˊ�!?*���9�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��O+�ٿ�~	����@��N���3@��9̐!?�B�w�2�@��dN��ٿ�� ���@Q��Pz�3@u�`ۼ�!?L�����@��dN��ٿ�� ���@Q��Pz�3@u�`ۼ�!?L�����@��dN��ٿ�� ���@Q��Pz�3@u�`ۼ�!?L�����@7�]��ٿI%�YB�@�)+D�3@����!?AVPz��@7�]��ٿI%�YB�@�)+D�3@����!?AVPz��@7�]��ٿI%�YB�@�)+D�3@����!?AVPz��@����ٿ�He+���@�� y��3@n���!?�bW*�O�@����ٿ�He+���@�� y��3@n���!?�bW*�O�@����ٿ�He+���@�� y��3@n���!?�bW*�O�@����ٿ�He+���@�� y��3@n���!?�bW*�O�@��B%�ٿ�Or�<�@;5q8��3@��j�Ӑ!?:v�iq�@��B%�ٿ�Or�<�@;5q8��3@��j�Ӑ!?:v�iq�@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@uŽ=�ٿ��Cc<�@���v��3@�%p켐!?�_����@Iڼ�ԥٿ�Dww6�@"SDO�3@.Eʷ�!?�j�	���@��	)��ٿ�f�O��@٨�{_�3@��P�S�!?f����@��	)��ٿ�f�O��@٨�{_�3@��P�S�!?f����@��	)��ٿ�f�O��@٨�{_�3@��P�S�!?f����@��	)��ٿ�f�O��@٨�{_�3@��P�S�!?f����@��	)��ٿ�f�O��@٨�{_�3@��P�S�!?f����@����ٿ��P�˖�@�v�t�3@�e�~��!?3�����@����ٿ��P�˖�@�v�t�3@�e�~��!?3�����@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�fv+��ٿ&M����@1����3@Ă�<Ő!?�k`�!�@�X�s��ٿQ�Ռ��@ӕ��3@P�Rʐ!?���s1�@�X�s��ٿQ�Ռ��@ӕ��3@P�Rʐ!?���s1�@�X�s��ٿQ�Ռ��@ӕ��3@P�Rʐ!?���s1�@�X�s��ٿQ�Ռ��@ӕ��3@P�Rʐ!?���s1�@����d�ٿ��g1���@yg1��3@�¡��!?��ѩ ��@����d�ٿ��g1���@yg1��3@�¡��!?��ѩ ��@����d�ٿ��g1���@yg1��3@�¡��!?��ѩ ��@����d�ٿ��g1���@yg1��3@�¡��!?��ѩ ��@0�!�Q�ٿ7~��z�@�,Qv �3@I ��!?�sV����@0�!�Q�ٿ7~��z�@�,Qv �3@I ��!?�sV����@0�!�Q�ٿ7~��z�@�,Qv �3@I ��!?�sV����@0�!�Q�ٿ7~��z�@�,Qv �3@I ��!?�sV����@0�!�Q�ٿ7~��z�@�,Qv �3@I ��!?�sV����@�;_�$�ٿ��銅��@�����3@(���!?�/@�;.�@�;_�$�ٿ��銅��@�����3@(���!?�/@�;.�@�;_�$�ٿ��銅��@�����3@(���!?�/@�;.�@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@Sps�L�ٿ����8��@�M	l��3@��B��!?s�I7��@��Kʠٿ���n=�@��zeC�3@@�|�!?�E娪g�@��Kʠٿ���n=�@��zeC�3@@�|�!?�E娪g�@��Kʠٿ���n=�@��zeC�3@@�|�!?�E娪g�@��Kʠٿ���n=�@��zeC�3@@�|�!?�E娪g�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@3"Im��ٿ�lP�@K���3@�>f��!?��a]�K�@��ڟ��ٿ,L+�[�@���|X�3@똯���!?��>s	��@�i��t�ٿ�8�ǋ��@�Sp���3@I�����!?b��dN�@�i��t�ٿ�8�ǋ��@�Sp���3@I�����!?b��dN�@O�U�.�ٿZ�O[�"�@o ����3@A�D���!?��]�}��@O�U�.�ٿZ�O[�"�@o ����3@A�D���!?��]�}��@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@&�x��ٿ�COG��@�|d�X�3@K�E���!?SkC �@��o9�ٿ{�7��@v�%��3@T��t͐!?�U_����@j$���ٿ:�Z��@ʹ��3@�n{�!?��NO��@j$���ٿ:�Z��@ʹ��3@�n{�!?��NO��@j$���ٿ:�Z��@ʹ��3@�n{�!?��NO��@j$���ٿ:�Z��@ʹ��3@�n{�!?��NO��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@S��Q�ٿiPy�a��@᭻��3@\�3j��!?S��o��@�����ٿ���I�F�@�XV�d�3@�����!?�'�齌�@�����ٿ���I�F�@�XV�d�3@�����!?�'�齌�@�����ٿ���I�F�@�XV�d�3@�����!?�'�齌�@�����ٿ���I�F�@�XV�d�3@�����!?�'�齌�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@��W��ٿ��"��<�@E~�ǵ�3@���娐!?m���t�@|6a`�ٿb9ǝ��@�ʵ��3@e��kː!?8Q�b��@|6a`�ٿb9ǝ��@�ʵ��3@e��kː!?8Q�b��@|6a`�ٿb9ǝ��@�ʵ��3@e��kː!?8Q�b��@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@XS7�B�ٿ�~�?��@mo�+�3@>�z>��!?["���B�@	�]�ٿ1����@Z�bU��3@t����!?H���\�@	�]�ٿ1����@Z�bU��3@t����!?H���\�@	�]�ٿ1����@Z�bU��3@t����!?H���\�@�榣ޡٿ���!E��@��̉�3@|��y��!?v�L�@�榣ޡٿ���!E��@��̉�3@|��y��!?v�L�@�i_��ٿ��nf�@=U�J&�3@}���I�!?6�5�@�i_��ٿ��nf�@=U�J&�3@}���I�!?6�5�@�i_��ٿ��nf�@=U�J&�3@}���I�!?6�5�@�A�ǜٿ��$Xy�@�L���3@;��~�!?�ce'�h�@�A�ǜٿ��$Xy�@�L���3@;��~�!?�ce'�h�@�A�ǜٿ��$Xy�@�L���3@;��~�!?�ce'�h�@�A�ǜٿ��$Xy�@�L���3@;��~�!?�ce'�h�@�A�ǜٿ��$Xy�@�L���3@;��~�!?�ce'�h�@b�����ٿT�f���@��,�F�3@� <��!?���q�@��De�ٿA%L�! �@�s����3@?%Y�t�!?LS^�!��@��De�ٿA%L�! �@�s����3@?%Y�t�!?LS^�!��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@@�P���ٿ��g���@d�G��3@j��/i�!?��4��@��ӕ�ٿ�TV�M��@��A,��3@�lZꈐ!?;�n�`��@��ӕ�ٿ�TV�M��@��A,��3@�lZꈐ!?;�n�`��@=��b5�ٿ������@���
�3@�	)퍐!?5#�D2�@���ٿ��ڪ��@�x��C�3@do9�ː!?5���@���ٿ��ڪ��@�x��C�3@do9�ː!?5���@���ٿ��ڪ��@�x��C�3@do9�ː!?5���@�լ.j�ٿ蟎��@��\�3@�>����!?5wO&�@�լ.j�ٿ蟎��@��\�3@�>����!?5wO&�@�լ.j�ٿ蟎��@��\�3@�>����!?5wO&�@�լ.j�ٿ蟎��@��\�3@�>����!?5wO&�@/�;L�ٿ�,��m��@�'Hb3�3@��9��!?��P�_�@/�;L�ٿ�,��m��@�'Hb3�3@��9��!?��P�_�@�n�6&�ٿyh�r�i�@M��3@��+Ő!?e2��$��@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@���X2�ٿ4�;�]�@�K�Հ�3@��(0��!?�wa���@n��v�ٿH�	O��@�^���3@jlQ�V�!?�1R~1�@n��v�ٿH�	O��@�^���3@jlQ�V�!?�1R~1�@ػ�\U�ٿQ9��@]�@����>�3@7u��y�!?�܀���@�H�/�ٿ�'�-���@+��L�3@�Il�!?"������@�H�/�ٿ�'�-���@+��L�3@�Il�!?"������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�&���ٿ���@"n��^�3@��[��!?������@�����ٿ���ai��@H��3@��d��!?������@�����ٿ���ai��@H��3@��d��!?������@�����ٿ���ai��@H��3@��d��!?������@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@4��ٿ�7Y�7s�@R�X�3@�q�!?�߽��@��=�ٿ��O�<��@��or�3@�1p���!?��u���@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�ʷ1�ٿ���ܩ��@�AX�3@����!?���+}�@�7��נٿ��pr��@��[�3@�ǋ�Ԑ!?r.d%�-�@wX�Wx�ٿ�t�:�@U�E�A�3@!�C��!?��z���@wX�Wx�ٿ�t�:�@U�E�A�3@!�C��!?��z���@wX�Wx�ٿ�t�:�@U�E�A�3@!�C��!?��z���@wX�Wx�ٿ�t�:�@U�E�A�3@!�C��!?��z���@wX�Wx�ٿ�t�:�@U�E�A�3@!�C��!?��z���@�C
6�ٿ*{Ï1�@y}���3@���pՐ!?@5�jB�@�C
6�ٿ*{Ï1�@y}���3@���pՐ!?@5�jB�@�C
6�ٿ*{Ï1�@y}���3@���pՐ!?@5�jB�@�C
6�ٿ*{Ï1�@y}���3@���pՐ!?@5�jB�@��̠ٿ"��
��@�g�M��3@��}ѐ!?��݇�@��̠ٿ"��
��@�g�M��3@��}ѐ!?��݇�@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@��כٿp��6�@q.��3@^�!?Np����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@*�$�њٿ��ҭ��@N�����3@Ŷ�z��!?'����@���1�ٿ�Q�/
�@P�I�3@��Cv��!?ǘ�=�n�@���1�ٿ�Q�/
�@P�I�3@��Cv��!?ǘ�=�n�@���1�ٿ�Q�/
�@P�I�3@��Cv��!?ǘ�=�n�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@�D�m�ٿ�M�@�@虮�j�3@�AԈ�!?���$�@��gk��ٿ��$��@��c�1�3@���_א!?��'4:��@��gk��ٿ��$��@��c�1�3@���_א!?��'4:��@��gk��ٿ��$��@��c�1�3@���_א!?��'4:��@��gk��ٿ��$��@��c�1�3@���_א!?��'4:��@����'�ٿ~��q��@馪h��3@9��3��!?��T��@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@N$��D�ٿ������@\S�1�3@��]Y��!?!���I�@��6��ٿ�/�����@(����3@C57ِ!?� ~��l�@��6��ٿ�/�����@(����3@C57ِ!?� ~��l�@��6��ٿ�/�����@(����3@C57ِ!?� ~��l�@��6��ٿ�/�����@(����3@C57ِ!?� ~��l�@��6��ٿ�/�����@(����3@C57ِ!?� ~��l�@���E�ٿt�/1��@u��I0�3@W u�!?�fk��@���E�ٿt�/1��@u��I0�3@W u�!?�fk��@Ax�M��ٿ�U/�@_��~n�3@�G���!?�V|*�@Ax�M��ٿ�U/�@_��~n�3@�G���!?�V|*�@Ax�M��ٿ�U/�@_��~n�3@�G���!?�V|*�@��j�_�ٿ$���d�@*�4�3@!!iG��!?`yn�w��@��j�_�ٿ$���d�@*�4�3@!!iG��!?`yn�w��@��j�_�ٿ$���d�@*�4�3@!!iG��!?`yn�w��@�l�YОٿ)�W
�V�@�~���3@�;���!?������@0� ��ٿE�u���@�����3@n'*��!?��uJ��@0� ��ٿE�u���@�����3@n'*��!?��uJ��@0� ��ٿE�u���@�����3@n'*��!?��uJ��@0� ��ٿE�u���@�����3@n'*��!?��uJ��@0� ��ٿE�u���@�����3@n'*��!?��uJ��@0� ��ٿE�u���@�����3@n'*��!?��uJ��@�];�a�ٿ)� N�{�@,J�m��3@�[��)�!?Q?��p��@�];�a�ٿ)� N�{�@,J�m��3@�[��)�!?Q?��p��@k񯕟�ٿ�OaRCM�@q����3@v6�Ր!?�j���@k񯕟�ٿ�OaRCM�@q����3@v6�Ր!?�j���@k񯕟�ٿ�OaRCM�@q����3@v6�Ր!?�j���@k񯕟�ٿ�OaRCM�@q����3@v6�Ր!?�j���@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@����ٿmN=�@�q�w�3@�����!?)���W��@�T㳭�ٿ�\N�I�@:Y
1��3@�S�U��!?x�k,�]�@/�`���ٿk�̚��@�Ha
��3@ ��)��!?�=��;�@�.]ޥٿ�~��.=�@�/�8(�3@,)H�$�!?����@�.]ޥٿ�~��.=�@�/�8(�3@,)H�$�!?����@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@}�P4�ٿMo2@�(�@����3@��R���!?���.7#�@���h��ٿ�*��0��@+�w���3@ ��co�!?�����@jf��,�ٿ�U�	o��@����3@�����!?"(� �@��Xڭ�ٿ�vx̓�@���#�3@���״�!?b>����@]Bc�Y�ٿ�;��|��@�8K> �3@�_,Ԑ!?�����~�@]Bc�Y�ٿ�;��|��@�8K> �3@�_,Ԑ!?�����~�@<2px��ٿ&�͟�@ϕ(���3@[]�S�!?zy�0��@<2px��ٿ&�͟�@ϕ(���3@[]�S�!?zy�0��@�����ٿ#�[����@F�pL�3@��l5Ɛ!?*<z�Z�@�����ٿ#�[����@F�pL�3@��l5Ɛ!?*<z�Z�@�b��ٿ�~���@=a>�W�3@��K��!?��L�>K�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@������ٿ:^"��*�@7Mn�3@e�5	�!?2 ��8�@��NƝٿ>�a�@�C�,�3@�8��!?J�a�P�@��NƝٿ>�a�@�C�,�3@�8��!?J�a�P�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@�^j�ٿ\�h���@�8Q@�3@U-l��!?���;�@���H�ٿ��r�"�@��5�>�3@�r{Xː!?��&��F�@���H�ٿ��r�"�@��5�>�3@�r{Xː!?��&��F�@���H�ٿ��r�"�@��5�>�3@�r{Xː!?��&��F�@Q�X��ٿ@��X�_�@<�h��3@���4ΐ!?T_�0���@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@���`E�ٿ�=��m��@Q�^x��3@ ��?Ð!?�5&�a�@��m,��ٿ������@ڌJ��3@!��켐!?z��΋�@��m,��ٿ������@ڌJ��3@!��켐!?z��΋�@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�&�E�ٿ�-���B�@���~�3@@a�'$�!?b��h���@�;�ۃ�ٿ*S���@C�'M��3@^�:"��!?Ć��@�;�ۃ�ٿ*S���@C�'M��3@^�:"��!?Ć��@�;�ۃ�ٿ*S���@C�'M��3@^�:"��!?Ć��@�;�ۃ�ٿ*S���@C�'M��3@^�:"��!?Ć��@nA���ٿ�R�C�Z�@��N$��3@K�s��!?�T1�ݒ�@nA���ٿ�R�C�Z�@��N$��3@K�s��!?�T1�ݒ�@nA���ٿ�R�C�Z�@��N$��3@K�s��!?�T1�ݒ�@�<�$��ٿژAvҾ�@�9��3@q�L��!?]��[�l�@B���Лٿ1����@����X�3@���w��!?O��V`�@B���Лٿ1����@����X�3@���w��!?O��V`�@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@ڳ�c�ٿΈɛ��@����3@�/�l��!?�l����@(��夡ٿ��5a�@���?�3@2�I��!?v���@(��夡ٿ��5a�@���?�3@2�I��!?v���@(��夡ٿ��5a�@���?�3@2�I��!?v���@(��夡ٿ��5a�@���?�3@2�I��!?v���@(��夡ٿ��5a�@���?�3@2�I��!?v���@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@���3?�ٿ��b�5$�@ZG!�Z�3@���!?�P�'�@�'��M�ٿ*p�V���@�LJ�e�3@�iw���!?
v\��@�'��M�ٿ*p�V���@�LJ�e�3@�iw���!?
v\��@�'��M�ٿ*p�V���@�LJ�e�3@�iw���!?
v\��@�'��M�ٿ*p�V���@�LJ�e�3@�iw���!?
v\��@�'��M�ٿ*p�V���@�LJ�e�3@�iw���!?
v\��@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@��8[�ٿ�!B�@�;0�3@Sn�d��!? N�V�@�k݀�ٿ�,Y)y�@J��w�3@��|��!?�?3�9�@�k݀�ٿ�,Y)y�@J��w�3@��|��!?�?3�9�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@|��z�ٿ�K�U��@0D�\�3@�R9���!?d�w�3y�@���t�ٿ��e�e�@�&�t�3@������!?�N�*���@���t�ٿ��e�e�@�&�t�3@������!?�N�*���@���t�ٿ��e�e�@�&�t�3@������!?�N�*���@�T.�}�ٿ�5!�R�@xoUC�3@:?��ː!?Ŷ�Q�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@ cݼI�ٿ�m���@bd_J�3@x5�y|�!?�.&�=^�@9CY0��ٿR����@­'U�3@�@�^��!?�RF�i�@9CY0��ٿR����@­'U�3@�@�^��!?�RF�i�@9CY0��ٿR����@­'U�3@�@�^��!?�RF�i�@kV
(�ٿ�_ڜd.�@U�yA�3@�;���!?�i?("��@kV
(�ٿ�_ڜd.�@U�yA�3@�;���!?�i?("��@kV
(�ٿ�_ڜd.�@U�yA�3@�;���!?�i?("��@kV
(�ٿ�_ڜd.�@U�yA�3@�;���!?�i?("��@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@�H�,�ٿ�h����@������3@EE@��!?/E-:ܻ�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@���ٿ��A��@�^K�3@K̄h!?�s< �O�@.�2>�ٿ�IxYK��@q��5��3@p��ː!?���5��@.�2>�ٿ�IxYK��@q��5��3@p��ː!?���5��@.�2>�ٿ�IxYK��@q��5��3@p��ː!?���5��@.�2>�ٿ�IxYK��@q��5��3@p��ː!?���5��@�2��ٿmJ�g��@���/7�3@Zg(���!?(�\�k�@�2��ٿmJ�g��@���/7�3@Zg(���!?(�\�k�@ ��xG�ٿؐ���@?���3@����D�!?XΑp8��@ ��xG�ٿؐ���@?���3@����D�!?XΑp8��@ ��xG�ٿؐ���@?���3@����D�!?XΑp8��@ ��xG�ٿؐ���@?���3@����D�!?XΑp8��@����ٿ�8W��@L[ :��3@�0�k�!?I-e�@����ٿ�8W��@L[ :��3@�0�k�!?I-e�@����ٿ�8W��@L[ :��3@�0�k�!?I-e�@����ٿ�8W��@L[ :��3@�0�k�!?I-e�@�y��	�ٿ#�q��Y�@�}`��3@|\,�z�!?!.��}��@���q�ٿ�.`��@�s�m��3@@&��!?V,�����@���q�ٿ�.`��@�s�m��3@@&��!?V,�����@���q�ٿ�.`��@�s�m��3@@&��!?V,�����@���q�ٿ�.`��@�s�m��3@@&��!?V,�����@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@�1ؘݞٿ��1�{�@=�۸��3@��T��!?g~��h��@?~y.r�ٿ�ZE4���@������3@��@Ր!?o�����@?~y.r�ٿ�ZE4���@������3@��@Ր!?o�����@?~y.r�ٿ�ZE4���@������3@��@Ր!?o�����@?~y.r�ٿ�ZE4���@������3@��@Ր!?o�����@?~y.r�ٿ�ZE4���@������3@��@Ր!?o�����@���F��ٿ'�����@���8�3@��`��!?��LV��@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@^5�燛ٿA�!��_�@���c�3@rW��!?	J����@1�46Ңٿm�i���@Q�=;�3@G����!?�� ��@1�46Ңٿm�i���@Q�=;�3@G����!?�� ��@�⌫��ٿ��H���@{\�5�3@�cx���!?GVW|�M�@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@DWh���ٿ�'&+`�@�Ϸ��3@������!?G0� �@r��h@�ٿ�v�37�@�ͻ��3@����!?O6�DGb�@r��h@�ٿ�v�37�@�ͻ��3@����!?O6�DGb�@���r�ٿ�� û`�@�$��3@�7'���!?pH��zr�@���r�ٿ�� û`�@�$��3@�7'���!?pH��zr�@�T���ٿ������@�E%h�3@�7���!?��3'�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@�Z��ٿ쇖�-��@� hq-�3@*�E��!?���q�!�@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@ߔ�"��ٿ�q���@�T\�~�3@&rub��!?�<�(��@\F�gۡٿa�����@��]d��3@�\�X^�!?��ҩ��@\F�gۡٿa�����@��]d��3@�\�X^�!?��ҩ��@����o�ٿ�yl�B��@��_S��3@qψp��!?f�_��@����o�ٿ�yl�B��@��_S��3@qψp��!?f�_��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@� =Q�ٿFO��@�%KB�3@�bU���!?RA�W��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�߸N;�ٿ�Px���@�\����3@|�'E�!?1I�u��@�C���ٿʫ����@����3@�Se���!?ƾ�$p�@i�J�ٿ��� �@v�p6��3@A��͐!?n �����@i�J�ٿ��� �@v�p6��3@A��͐!?n �����@i�J�ٿ��� �@v�p6��3@A��͐!?n �����@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@+�?�ٿH,��`@�@Gt?F�3@%�{��!?Df�O��@6B,n��ٿ~K���@5�L�q�3@k�X{��!?��[W���@6B,n��ٿ~K���@5�L�q�3@k�X{��!?��[W���@6B,n��ٿ~K���@5�L�q�3@k�X{��!?��[W���@6B,n��ٿ~K���@5�L�q�3@k�X{��!?��[W���@6B,n��ٿ~K���@5�L�q�3@k�X{��!?��[W���@B��ٿ�g�j�@d�C��3@��ߕ�!?:��8;�@B��ٿ�g�j�@d�C��3@��ߕ�!?:��8;�@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@U��ٿa	���W�@5wp��3@�Y��!?�����@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@--�+z�ٿ��P��@�[<��3@�E3�z�!?��9�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@=>P��ٿ��3s�"�@�og��3@I���!?$�{�"�@�����ٿ3�:���@�^u�C�3@�ҵ��!?�¶0V�@�����ٿ3�:���@�^u�C�3@�ҵ��!?�¶0V�@/ͯN�ٿ�෺d��@&���e�3@2�R��!?r���\�@��ϲ,�ٿT�G}���@-,�3@��_��!?B;{-,��@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@w1�?��ٿ��'D��@�B
�1�3@sU���!?������@g�]�ٿPV�^@B�@A����3@�<� �!?�'���@�c�Ȅ�ٿ����@����E�3@Ɋ��!?|tX��@�c�Ȅ�ٿ����@����E�3@Ɋ��!?|tX��@�c�Ȅ�ٿ����@����E�3@Ɋ��!?|tX��@�c�Ȅ�ٿ����@����E�3@Ɋ��!?|tX��@�c�Ȅ�ٿ����@����E�3@Ɋ��!?|tX��@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@Y��)y�ٿ¬�js�@�����3@��x���!?h+<�$�@��+e�ٿ�Su��@�5����3@��d�t�!?_����@��+e�ٿ�Su��@�5����3@��d�t�!?_����@��+e�ٿ�Su��@�5����3@��d�t�!?_����@��+e�ٿ�Su��@�5����3@��d�t�!?_����@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@]Y���ٿ6dёLo�@�]GkY�3@�?�S��!?������@Q8�W�ٿ���>u"�@Y�C�3@��f!v�!?������@Q8�W�ٿ���>u"�@Y�C�3@��f!v�!?������@Q8�W�ٿ���>u"�@Y�C�3@��f!v�!?������@Q8�W�ٿ���>u"�@Y�C�3@��f!v�!?������@by�^p�ٿs� ҁ�@���k�3@M�9���!?����a�@����F�ٿ!b�]�@�N��3@l��9̐!?L�8X��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@�7��ٿ'v�_��@���	��3@�S�� �!?��
�~��@��鬞ٿ�;��&�@�!���3@e����!?Y3KƳ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@���狢ٿ{�����@GYF���3@̓�{�!?�Nʘ�@ ��(-�ٿᯮ���@֙*�3@AxA˿�!?�C�V��@ ��(-�ٿᯮ���@֙*�3@AxA˿�!?�C�V��@ ��(-�ٿᯮ���@֙*�3@AxA˿�!?�C�V��@ ��(-�ٿᯮ���@֙*�3@AxA˿�!?�C�V��@ ��(-�ٿᯮ���@֙*�3@AxA˿�!?�C�V��@�X�ٿ�����k�@�y�Q�3@l�e�ِ!?U����@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@J���؜ٿ�8 ���@T*=Sj�3@���ِ!?�C�%�@�]aեٿԙo�x��@�����3@��z�!?1��M���@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@�Bf���ٿI�)�5x�@i/N���3@t���Ő!?Rؠ�[!�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@���7z�ٿ��6r��@/�`:��3@�v�<�!?��1^\q�@y���j�ٿ��l%��@p��3*�3@�6�N	�!?hɔޙ	�@y���j�ٿ��l%��@p��3*�3@�6�N	�!?hɔޙ	�@y���j�ٿ��l%��@p��3*�3@�6�N	�!?hɔޙ	�@y���j�ٿ��l%��@p��3*�3@�6�N	�!?hɔޙ	�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@,-�?�ٿ͡oH���@,��4�3@ b�� �!?L�5�J#�@:���ٿؔ?j)�@��,J�3@��� �!?�����O�@:���ٿؔ?j)�@��,J�3@��� �!?�����O�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@��('�ٿ0`���@H��q{�3@�[�h��!?P9c�j@�@�
�1��ٿ:̅�v�@#���3@�er��!?�gNrb�@�
�1��ٿ:̅�v�@#���3@�er��!?�gNrb�@�
�1��ٿ:̅�v�@#���3@�er��!?�gNrb�@a:�.�ٿ���d�@��D��3@l4���!?7�5���@a:�.�ٿ���d�@��D��3@l4���!?7�5���@a:�.�ٿ���d�@��D��3@l4���!?7�5���@a:�.�ٿ���d�@��D��3@l4���!?7�5���@a:�.�ٿ���d�@��D��3@l4���!?7�5���@a:�.�ٿ���d�@��D��3@l4���!?7�5���@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@Ϲ�Cp�ٿ���`X�@���\�3@�L����!?:1�7�@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@:�4���ٿ
2|����@��TH��3@�S���!?�iR8��@g���ٿ�3Cal��@�����3@��9ܐ!?�h!m���@g���ٿ�3Cal��@�����3@��9ܐ!?�h!m���@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@P{�gߞٿg4�0���@���D�3@�A�ʐ!?���B�@!Z�ٿ�����@%���3@f>Ԑ!?B;�x!�@!Z�ٿ�����@%���3@f>Ԑ!?B;�x!�@O��ܹ�ٿ����F�@y�)��3@�9�֐!?�_�Y�*�@O��ܹ�ٿ����F�@y�)��3@�9�֐!?�_�Y�*�@�_

	�ٿ��W4��@�0k�E�3@��5��!?�B�+�@�_

	�ٿ��W4��@�0k�E�3@��5��!?�B�+�@�_

	�ٿ��W4��@�0k�E�3@��5��!?�B�+�@�_

	�ٿ��W4��@�0k�E�3@��5��!?�B�+�@�_

	�ٿ��W4��@�0k�E�3@��5��!?�B�+�@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�]l^�ٿ���^��@�vK�X�3@�11,�!? C�׺��@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@�a"��ٿ���K�@Y��R�3@��f��!?�[��w�@r� �T�ٿ�wb�9y�@d�4=�3@�k���!?�c:Vq�@r� �T�ٿ�wb�9y�@d�4=�3@�k���!?�c:Vq�@r� �T�ٿ�wb�9y�@d�4=�3@�k���!?�c:Vq�@�:����ٿ`ʮ��@�*����3@�6+�!?��4���@�:����ٿ`ʮ��@�*����3@�6+�!?��4���@vx�_ٟٿq��6|��@�Ӏ���3@&����!?N��6��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@R�g�ٿ�����@�67�V�3@�j:���!?Ԯ�x��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@�;t�*�ٿf�	x;��@�INq��3@𘏴��!?�ͫ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@|�eC�ٿ�-Y�>�@�X�@�3@:�J��!?���aZ��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@�L}O�ٿz��,�h�@�}=�8�3@�A���!?,e�r��@���|��ٿ�-6���@���i�3@G_����!?�rt_��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@��U�ٿH�߭X��@>��N�3@�	?А!?�r�4��@?ꉇd�ٿ�6�7�@�����3@������!?\M/TC�@?ꉇd�ٿ�6�7�@�����3@������!?\M/TC�@�w�ܨٿXO>���@���u��3@֑���!?�a7�"�@ �r�Z�ٿ��h>�!�@,-�&�3@���ݐ!?�����M�@ �r�Z�ٿ��h>�!�@,-�&�3@���ݐ!?�����M�@ �r�Z�ٿ��h>�!�@,-�&�3@���ݐ!?�����M�@ �r�Z�ٿ��h>�!�@,-�&�3@���ݐ!?�����M�@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@����ٿb���p�@CL��3@U>1���!?������@[��3I�ٿ˳k���@֚�)0�3@Ry��	�!?=s���@[��3I�ٿ˳k���@֚�)0�3@Ry��	�!?=s���@[��3I�ٿ˳k���@֚�)0�3@Ry��	�!?=s���@[��3I�ٿ˳k���@֚�)0�3@Ry��	�!?=s���@�*�ٿ���I^��@J���3@�A$��!?�o���.�@�*�ٿ���I^��@J���3@�A$��!?�o���.�@�*�ٿ���I^��@J���3@�A$��!?�o���.�@�*�ٿ���I^��@J���3@�A$��!?�o���.�@�*�ٿ���I^��@J���3@�A$��!?�o���.�@�L��%�ٿ(>�?�@8;��c�3@"����!?S���.��@�a�(�ٿ1����@��-���3@�.���!?�G��$��@�a�(�ٿ1����@��-���3@�.���!?�G��$��@�a�(�ٿ1����@��-���3@�.���!?�G��$��@�}SZ�ٿ�L�3��@�%�G�3@��L��!?����@v��ٿ���c�4�@	�f�6�3@��-6��!?�����|�@v��ٿ���c�4�@	�f�6�3@��-6��!?�����|�@v��ٿ���c�4�@	�f�6�3@��-6��!?�����|�@v��ٿ���c�4�@	�f�6�3@��-6��!?�����|�@a��8֟ٿW2�d��@U�f��3@D�Ǹ�!?�M�~�@a��8֟ٿW2�d��@U�f��3@D�Ǹ�!?�M�~�@a��8֟ٿW2�d��@U�f��3@D�Ǹ�!?�M�~�@a��8֟ٿW2�d��@U�f��3@D�Ǹ�!?�M�~�@a��8֟ٿW2�d��@U�f��3@D�Ǹ�!?�M�~�@!��i�ٿ>�m�Z�@�����3@l.\���!?��>װ�@!��i�ٿ>�m�Z�@�����3@l.\���!?��>װ�@!��i�ٿ>�m�Z�@�����3@l.\���!?��>װ�@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@N�A��ٿ���)�@I~ϷI�3@��]o�!?6������@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@^���8�ٿ�^����@_��U�3@OE�9��!?E�mY�@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�x"/ʙٿ�`i�'�@���)h�3@orm��!?/��g��@�p���ٿ,r޷̠�@b�Y5��3@������!?`�0mG�@�p���ٿ,r޷̠�@b�Y5��3@������!?`�0mG�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@�ׂ��ٿ�0���@���Q<�3@\ξ�!?�,�qs�@��25R�ٿ����@��� ��3@����!?t�8��@��25R�ٿ����@��� ��3@����!?t�8��@��25R�ٿ����@��� ��3@����!?t�8��@���r_�ٿ����W?�@���My�3@e��f��!?�z����@���r_�ٿ����W?�@���My�3@e��f��!?�z����@���r_�ٿ����W?�@���My�3@e��f��!?�z����@���r_�ٿ����W?�@���My�3@e��f��!?�z����@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@tb8��ٿ�Q���"�@��J�e�3@,=�ǐ!?O��i���@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�ъ (�ٿ����5�@�޳���3@D~�x��!?0t6����@�J<�E�ٿ���@���@۝��n�3@�����!?��l�h��@�J<�E�ٿ���@���@۝��n�3@�����!?��l�h��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@�ƹ�ٿ�X8Bx�@f� ��3@�I_А!?�IC(>��@eU^��ٿhQ���@m�����3@U*���!?���xk��@��e;Ӡٿ�����@��3S��3@�H��Ő!?V�A��@��e;Ӡٿ�����@��3S��3@�H��Ő!?V�A��@��e;Ӡٿ�����@��3S��3@�H��Ő!?V�A��@��e;Ӡٿ�����@��3S��3@�H��Ő!?V�A��@��e;Ӡٿ�����@��3S��3@�H��Ő!?V�A��@����ٿ�M�b��@�Q���3@:�c�!?�J����@����ٿ�M�b��@�Q���3@:�c�!?�J����@�r��ٿ�Tj�@$�'��3@T0���!?�ah]V*�@�\��ٿ) (&�@V���3@7y���!?�[�XM�@�\��ٿ) (&�@V���3@7y���!?�[�XM�@�\��ٿ) (&�@V���3@7y���!?�[�XM�@J{��Z�ٿt�%G��@+	Ձ��3@9�zѐ!?	���+�@�a�%G�ٿ�M-H��@{����3@v��d�!?��]�V�@�a�%G�ٿ�M-H��@{����3@v��d�!?��]�V�@���)=�ٿ�K�	�@�Aߎ��3@�لDÐ!?R�W���@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@��-P�ٿl�@T��@��3@T�Ú�!?�'߲R��@@��ߜٿFV����@�i'��3@�5��!?<I����@@��ߜٿFV����@�i'��3@�5��!?<I����@@��ߜٿFV����@�i'��3@�5��!?<I����@K�rɟٿ*����@L�rς�3@� �!?[����@K�rɟٿ*����@L�rς�3@� �!?[����@ag��'�ٿ�1]}���@�7ƾ`�3@��l=Ґ!?�e�I���@ag��'�ٿ�1]}���@�7ƾ`�3@��l=Ґ!?�e�I���@�Mn�)�ٿ�v��v��@��
���3@������!?� ����@�Mn�)�ٿ�v��v��@��
���3@������!?� ����@�Mn�)�ٿ�v��v��@��
���3@������!?� ����@�Mn�)�ٿ�v��v��@��
���3@������!?� ����@�Mn�)�ٿ�v��v��@��
���3@������!?� ����@���_ �ٿ6��*���@4����3@�I��!?8ƈ���@�YB
O�ٿ?j�U�%�@�P#9��3@
�h��!?�ً��a�@���>�ٿ%$X�U��@§����3@�Y�E��!?��8-��@���>�ٿ%$X�U��@§����3@�Y�E��!?��8-��@���>�ٿ%$X�U��@§����3@�Y�E��!?��8-��@���>�ٿ%$X�U��@§����3@�Y�E��!?��8-��@m�!^�ٿ��a~A��@�����3@I��S��!?��=���@m�!^�ٿ��a~A��@�����3@I��S��!?��=���@i��7�ٿ����i�@�A�3@����!?�ڛ�*�@i��7�ٿ����i�@�A�3@����!?�ڛ�*�@�<�ou�ٿ�FJD`��@���t�3@�R��ː!?���$+�@�<�ou�ٿ�FJD`��@���t�3@�R��ː!?���$+�@�<�ou�ٿ�FJD`��@���t�3@�R��ː!?���$+�@��?�X�ٿev��o.�@M�W��3@5<<�!?G- �7`�@�]�_�ٿR#-$���@�����3@Sb��!?��#A���@�]�_�ٿR#-$���@�����3@Sb��!?��#A���@�]�_�ٿR#-$���@�����3@Sb��!?��#A���@�1_���ٿʻִ�%�@�Z?ޔ�3@�#����!?�ln���@�1_���ٿʻִ�%�@�Z?ޔ�3@�#����!?�ln���@���i�ٿ2�3蠵�@m'J���3@�H:���!?�^�랥�@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@�E|:<�ٿ�R	�7�@h�x@k�3@���Ő!?���H��@:eZu7�ٿ]`bD�@�h����3@ �kxݐ!?^ ��b��@:eZu7�ٿ]`bD�@�h����3@ �kxݐ!?^ ��b��@:eZu7�ٿ]`bD�@�h����3@ �kxݐ!?^ ��b��@:eZu7�ٿ]`bD�@�h����3@ �kxݐ!?^ ��b��@:eZu7�ٿ]`bD�@�h����3@ �kxݐ!?^ ��b��@��[�ٿ��}M��@�l) �3@���xА!?�Uf� �@��[�ٿ��}M��@�l) �3@���xА!?�Uf� �@��[�ٿ��}M��@�l) �3@���xА!?�Uf� �@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@Gx� �ٿ��m=�@��cL�3@�$��!?�&�cq�@8��l`�ٿ�dETje�@4BUb�3@ �����!?$��.�r�@8��l`�ٿ�dETje�@4BUb�3@ �����!?$��.�r�@�dW�,�ٿdǆm1|�@���Ǔ�3@YBM�ސ!?.�Y���@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@�z�R0�ٿ��\�:��@��95�3@9�|�ѐ!?r(��		�@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@3�K�M�ٿ�T4�@���R�3@�X����!?v���@]�xƳ�ٿG���s�@�F���3@{��q��!? p�]��@]�xƳ�ٿG���s�@�F���3@{��q��!? p�]��@]�xƳ�ٿG���s�@�F���3@{��q��!? p�]��@�a��ٿ��T�`��@�F�d3�3@V����!?��X���@�a��ٿ��T�`��@�F�d3�3@V����!?��X���@�a��ٿ��T�`��@�F�d3�3@V����!?��X���@�a��ٿ��T�`��@�F�d3�3@V����!?��X���@�a��ٿ��T�`��@�F�d3�3@V����!?��X���@`R\��ٿץ���l�@p����3@&Z#�ߐ!?"��P�@�zj��ٿ-CG��@ԥ��3@͒_��!?n<!K��@�zj��ٿ-CG��@ԥ��3@͒_��!?n<!K��@�zj��ٿ-CG��@ԥ��3@͒_��!?n<!K��@�zj��ٿ-CG��@ԥ��3@͒_��!?n<!K��@�zj��ٿ-CG��@ԥ��3@͒_��!?n<!K��@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@���ٿXc4i��@Ә'�%�3@;�1֣�!?��a����@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@n��%E�ٿ1-et�@���ʑ�3@D�TŐ!?�d�u�c�@��_E[�ٿ�����@���3@�(�Mِ!?��i~h��@տ_)��ٿ�Ir�t��@b��3@��G�!?&$�궺�@տ_)��ٿ�Ir�t��@b��3@��G�!?&$�궺�@տ_)��ٿ�Ir�t��@b��3@��G�!?&$�궺�@��͉�ٿ�>���J�@�`�|J�3@ ���!?W�K����@��͉�ٿ�>���J�@�`�|J�3@ ���!?W�K����@��͉�ٿ�>���J�@�`�|J�3@ ���!?W�K����@ D�B�ٿ�V%����@򸷕��3@��䀟�!?X��*��@4��y�ٿ�+����@L�S�>�3@ᲞG��!?)������@4��y�ٿ�+����@L�S�>�3@ᲞG��!?)������@4��y�ٿ�+����@L�S�>�3@ᲞG��!?)������@ɼ8���ٿa��#�O�@�����3@$�|��!?�g5���@ɼ8���ٿa��#�O�@�����3@$�|��!?�g5���@��[;�ٿ�=�k��@Z��$b�3@��d���!?�57�f��@��[;�ٿ�=�k��@Z��$b�3@��d���!?�57�f��@��[;�ٿ�=�k��@Z��$b�3@��d���!?�57�f��@��[;�ٿ�=�k��@Z��$b�3@��d���!?�57�f��@��[;�ٿ�=�k��@Z��$b�3@��d���!?�57�f��@�����ٿ	O/���@a�	��3@qby��!?���Ƒ�@�X���ٿ	��&���@�|�û�3@��k���!?t�і���@�X���ٿ	��&���@�|�û�3@��k���!?t�і���@�X���ٿ	��&���@�|�û�3@��k���!?t�і���@�X���ٿ	��&���@�|�û�3@��k���!?t�і���@�X���ٿ	��&���@�|�û�3@��k���!?t�і���@̬��ܟٿ�1C7��@}��^�3@�9����!?Q���w��@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@*�gC�ٿ5�Iq#��@�&�/�3@K����!?�����@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@3����ٿPI{.f�@����3@b8���!?�P?I��@��O�ٿ4j��@*6�	�3@?,����!?
��U�@��O�ٿ4j��@*6�	�3@?,����!?
��U�@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@��H�n�ٿҙ���@�;_�;�3@ﻚӍ�!?��&ݲ��@(�	�P�ٿ ���^�@��&���3@���Ȑ!? R�x��@(�	�P�ٿ ���^�@��&���3@���Ȑ!? R�x��@(�'�ٿs+7d�@��!���3@Ek�ѐ!?�hV�lz�@(�'�ٿs+7d�@��!���3@Ek�ѐ!?�hV�lz�@(�'�ٿs+7d�@��!���3@Ek�ѐ!?�hV�lz�@�m��ٿvƚ��-�@���3��3@�E���!?�U5���@�m��ٿvƚ��-�@���3��3@�E���!?�U5���@�`0Ƞٿҥ4�@&�@��s��3@���֐!?��i2w��@�`0Ƞٿҥ4�@&�@��s��3@���֐!?��i2w��@�`0Ƞٿҥ4�@&�@��s��3@���֐!?��i2w��@�`0Ƞٿҥ4�@&�@��s��3@���֐!?��i2w��@�Q^�Z�ٿ���[�w�@#D��3@�P���!?�ڢ���@�Q^�Z�ٿ���[�w�@#D��3@�P���!?�ڢ���@�Q^�Z�ٿ���[�w�@#D��3@�P���!?�ڢ���@�Q^�Z�ٿ���[�w�@#D��3@�P���!?�ڢ���@@R�&�ٿL��/A�@��d��3@=����!?�A$���@(�1���ٿ��$�@0�5���3@]�u�!?�Na_)�@(�1���ٿ��$�@0�5���3@]�u�!?�Na_)�@(�1���ٿ��$�@0�5���3@]�u�!?�Na_)�@(�1���ٿ��$�@0�5���3@]�u�!?�Na_)�@{a�ٿc�Ϙ�@v�D���3@�_.��!?��+X��@��>�,�ٿ8+����@@��pR�3@bP�y�!?�v)�@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�z(b�ٿ�{i�@�C�"R�3@���ΐ!?f��ɚ��@�|�{\�ٿXx)	��@�wf'�3@������!?@�4��,�@�|�{\�ٿXx)	��@�wf'�3@������!?@�4��,�@�|�{\�ٿXx)	��@�wf'�3@������!?@�4��,�@�5�f��ٿ�ꮛ��@��*2H�3@���|��!?�V��x!�@�Pf���ٿRL���@=�J��3@޴
���!?(�_K��@�Pf���ٿRL���@=�J��3@޴
���!?(�_K��@�Pf���ٿRL���@=�J��3@޴
���!?(�_K��@P�Lm�ٿ���Oe��@�kf���3@�7�N��!?�HQ�o�@P�Lm�ٿ���Oe��@�kf���3@�7�N��!?�HQ�o�@>C�W�ٿ}�tZU��@S/���3@M��ki�!?7�U<`��@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�|�q�ٿ�����@#�j��3@{d���!?]i�zׁ�@�?�9��ٿ�|I=2��@D�%G�3@���!?� Ա���@�?�9��ٿ�|I=2��@D�%G�3@���!?� Ա���@�?�9��ٿ�|I=2��@D�%G�3@���!?� Ա���@�l�NРٿ��r��J�@%Z����3@E��	�!?С��U��@ ����ٿ��}���@S�^�c�3@���r��!?g_X9X��@ ����ٿ��}���@S�^�c�3@���r��!?g_X9X��@(Գq��ٿ�u��QC�@�S���3@P�!?���/�@(Գq��ٿ�u��QC�@�S���3@P�!?���/�@C����ٿ<c�%��@��n��3@�X~�!?����E�@C����ٿ<c�%��@��n��3@�X~�!?����E�@C����ٿ<c�%��@��n��3@�X~�!?����E�@���ٿ�����@sh{��3@�tb2��!?�����1�@���ٿ�����@sh{��3@�tb2��!?�����1�@���ٿ�����@sh{��3@�tb2��!?�����1�@���ٿ�����@sh{��3@�tb2��!?�����1�@���ٿ�����@sh{��3@�tb2��!?�����1�@���ٿ�����@sh{��3@�tb2��!?�����1�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@y����ٿ��j FK�@C����3@e�Q=�!?8�
2OV�@	�ۇ��ٿ[�
F��@ާX�B�3@3�|��!?� ��(�@	�ۇ��ٿ[�
F��@ާX�B�3@3�|��!?� ��(�@	�ۇ��ٿ[�
F��@ާX�B�3@3�|��!?� ��(�@�ś�åٿ�z�#-�@]��4�3@~4��Ɛ!?L=�~�@�Ss(�ٿ9��4�@�q����3@{���!?y1��>�@g�J�=�ٿ���Y��@��u��3@�N�А!?��:���@�i���ٿ�8�W��@�X����3@Q�)��!?��zG���@�i���ٿ�8�W��@�X����3@Q�)��!?��zG���@�i���ٿ�8�W��@�X����3@Q�)��!?��zG���@��D��ٿS����@|b�EB�3@���⢐!?Jg�	���@��V�r�ٿ�#A9�@�&����3@2cM�!?�T�Ad��@��rѶ�ٿ�}؆,�@�Lv�z�3@��Nِ!?�7</*�@��rѶ�ٿ�}؆,�@�Lv�z�3@��Nِ!?�7</*�@��rѶ�ٿ�}؆,�@�Lv�z�3@��Nِ!?�7</*�@��rѶ�ٿ�}؆,�@�Lv�z�3@��Nِ!?�7</*�@��rѶ�ٿ�}؆,�@�Lv�z�3@��Nِ!?�7</*�@�b��x�ٿ�@(N��@�yV�3@�
{�!?�L���_�@�b��x�ٿ�@(N��@�yV�3@�
{�!?�L���_�@�5�g�ٿ�5,�z�@�hU���3@0CȎ��!?f����W�@�5�g�ٿ�5,�z�@�hU���3@0CȎ��!?f����W�@�5�g�ٿ�5,�z�@�hU���3@0CȎ��!?f����W�@�5�g�ٿ�5,�z�@�hU���3@0CȎ��!?f����W�@�5�g�ٿ�5,�z�@�hU���3@0CȎ��!?f����W�@	��ٿR�Ad
�@���]��3@��ސ!?36q�@��Y5�ٿ�ʸV���@���Kv�3@�1dF֐!?����u��@��Y5�ٿ�ʸV���@���Kv�3@�1dF֐!?����u��@��Y5�ٿ�ʸV���@���Kv�3@�1dF֐!?����u��@��Y5�ٿ�ʸV���@���Kv�3@�1dF֐!?����u��@9Vi~��ٿ8���w�@�|����3@�]>ʐ!?�*����@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@䛗�t�ٿ�V����@`�t0!�3@�����!?�[���@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@���c]�ٿO�;���@2��IA�3@�Q듻�!?���{&�@�����ٿ���
-q�@��0G~�3@|M�'��!?w�o�.T�@�����ٿ���
-q�@��0G~�3@|M�'��!?w�o�.T�@�����ٿ���
-q�@��0G~�3@|M�'��!?w�o�.T�@�����ٿ���
-q�@��0G~�3@|M�'��!?w�o�.T�@�����ٿ���
-q�@��0G~�3@|M�'��!?w�o�.T�@gn�`�ٿUh�|�6�@A$4�"�3@��	ѐ!?	�]�.�@gn�`�ٿUh�|�6�@A$4�"�3@��	ѐ!?	�]�.�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@Z��ٿcH5=�@�v�`X�3@l�2x�!?�8,N�]�@o��|9�ٿSI�2c�@��щ��3@<fh��!?���n��@o��|9�ٿSI�2c�@��щ��3@<fh��!?���n��@o��|9�ٿSI�2c�@��щ��3@<fh��!?���n��@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@׌6i�ٿ�j����@q	
�f�3@�	��!?����c�@���&�ٿ�A]{�@�!&>��3@ӱ6��!?��s����@��%�!�ٿ�;T�!��@�?��e�3@E	վ�!?�����@5��$>�ٿ������@,��'��3@7�#͌�!?~�����@5��$>�ٿ������@,��'��3@7�#͌�!?~�����@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@XBg���ٿ��⊬��@^����3@�r�,F�!?�8�ݯ��@��i�6�ٿ݀�/��@7�4���3@��c�[�!?��'9��@���n�ٿ�l���@�D�4T�3@wE�V�!?C=A"�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�q����ٿ�z�~e��@/��k�3@t܈���!?}AAZ�@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�b�8��ٿ֞����@Y����3@�	����!?������@�$���ٿ�*^:�1�@�N��3@�Ր!?��Q$'�@�$���ٿ�*^:�1�@�N��3@�Ր!?��Q$'�@�$���ٿ�*^:�1�@�N��3@�Ր!?��Q$'�@�$���ٿ�*^:�1�@�N��3@�Ր!?��Q$'�@�$���ٿ�*^:�1�@�N��3@�Ր!?��Q$'�@��y�ٿ-D����@�x/��3@}z�B�!?��P���@��y�ٿ-D����@�x/��3@}z�B�!?��P���@7�;���ٿ�z�����@&�����3@]���!?��y�e�@7�;���ٿ�z�����@&�����3@]���!?��y�e�@7�;���ٿ�z�����@&�����3@]���!?��y�e�@�0�ўٿ��K
[��@0\ ��3@��P,ؐ!?�=^���@�0�ўٿ��K
[��@0\ ��3@��P,ؐ!?�=^���@'vd��ٿ���1D�@�W>:��3@��k�ʐ!?��*q/��@'vd��ٿ���1D�@�W>:��3@��k�ʐ!?��*q/��@'vd��ٿ���1D�@�W>:��3@��k�ʐ!?��*q/��@<�\ϻ�ٿ�� �>�@m��W�3@�t�!?��F����@<�\ϻ�ٿ�� �>�@m��W�3@�t�!?��F����@<�\ϻ�ٿ�� �>�@m��W�3@�t�!?��F����@<�\ϻ�ٿ�� �>�@m��W�3@�t�!?��F����@<�\ϻ�ٿ�� �>�@m��W�3@�t�!?��F����@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@|���ٿf��?��@�s�N�3@�C�͐!?�������@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@U~mu]�ٿI��Wu�@�t��3@�u����!?>c���@q�nS��ٿ��P;��@|�2��3@`\�o�!?ȴ!����@r�d;�ٿ	J���X�@�*x���3@!�Ȑ!?u̽J�@r�d;�ٿ	J���X�@�*x���3@!�Ȑ!?u̽J�@r�d;�ٿ	J���X�@�*x���3@!�Ȑ!?u̽J�@r�d;�ٿ	J���X�@�*x���3@!�Ȑ!?u̽J�@r�d;�ٿ	J���X�@�*x���3@!�Ȑ!?u̽J�@�4��ٿV0���@�_2���3@����!?�{��q�@��B�ٿ�V��4��@��)s�3@�����!?�ﷵ��@��B�ٿ�V��4��@��)s�3@�����!?�ﷵ��@��B�ٿ�V��4��@��)s�3@�����!?�ﷵ��@��B�ٿ�V��4��@��)s�3@�����!?�ﷵ��@҄&k��ٿ3���q�@б���3@ɶސ!?j�����@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@��\$[�ٿ��B'r�@?&����3@]pqߐ!?��z��@�.Q�Ρٿ �$z��@��X���3@�׫���!?tV��4�@�.Q�Ρٿ �$z��@��X���3@�׫���!?tV��4�@o�8��ٿT����@�;�!�3@��E�!?��F�v��@�3�N�ٿ����'��@�����3@��~cǐ!?�\�����@�3�N�ٿ����'��@�����3@��~cǐ!?�\�����@c�lH�ٿj0���h�@A�Y��3@_�Î��!?1��m�@��f�b�ٿ�l䭎��@���2��3@��ݛې!?�����@��f�b�ٿ�l䭎��@���2��3@��ݛې!?�����@��f�b�ٿ�l䭎��@���2��3@��ݛې!?�����@:U����ٿy,��%�@u̮�	�3@E��!?���W��@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@��ͻ3�ٿ��R�[B�@3]B�R�3@�}+��!?�2��'z�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@䬪Lw�ٿ7A��&��@;����3@���S��!?�Ԡ��P�@���p�ٿS�0�SP�@ٞ�L��3@��sE֐!?�	P�t3�@���p�ٿS�0�SP�@ٞ�L��3@��sE֐!?�	P�t3�@���0�ٿNd�gq�@7��~��3@�stC��!?.�e����@���0�ٿNd�gq�@7��~��3@�stC��!?.�e����@���0�ٿNd�gq�@7��~��3@�stC��!?.�e����@����ٿ��Y���@?���3@�*�$Ő!?�ԝS1�@����ٿ��Y���@?���3@�*�$Ő!?�ԝS1�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@crdc�ٿ��e�@�y
��3@�.[��!?�a4M=s�@���s�ٿ/���v��@/��!�3@Ѣx��!?ߊ���"�@���s�ٿ/���v��@/��!�3@Ѣx��!?ߊ���"�@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@��/i!�ٿR{��<8�@m>e�3@��6-��!?�k��Q��@����ٿ�m��� �@&C�*�3@w�a�f�!?���U0�@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��Jz˥ٿ:��<��@ѹ_��3@����Ð!?鷎P"��@��6�ҝٿ5���Y��@v����3@u"����!?�]�k�4�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@hn��Уٿ\%4��z�@9����3@�\[���!?��M�2�@�h#[A�ٿbZu����@/�Wg6�3@s'z(�!?�ݬ��X�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@�H懟ٿ�	D��@�����3@�nS�!?J8���n�@z�yCL�ٿ�K�E��@�AK�s�3@����!?+�y7�@��2U�ٿ��K_�@�����3@K2�8��!?�l��*��@�CȄʤٿ�;|�1��@�~ں�3@��g$ِ!?�cr���@�CȄʤٿ�;|�1��@�~ں�3@��g$ِ!?�cr���@�CȄʤٿ�;|�1��@�~ں�3@��g$ِ!?�cr���@�CȄʤٿ�;|�1��@�~ں�3@��g$ِ!?�cr���@�CȄʤٿ�;|�1��@�~ں�3@��g$ِ!?�cr���@��c֟ٿ�п��@����l�3@ʶv�p�!?!���@��c֟ٿ�п��@����l�3@ʶv�p�!?!���@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@R�	�ٿ�U���@.�<9��3@��>��!?��r�g��@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@b��ٿ��YY�U�@��zp��3@�kɐ!?�d���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@{54��ٿey�W��@T
̊��3@��P��!?��\���@)���Ȧٿ��D��@���	�3@{��!?�2�����@)���Ȧٿ��D��@���	�3@{��!?�2�����@0\��T�ٿ�$A�F4�@�B�av�3@4ﮘ��!?�_���_�@zUn6��ٿ+�z��@�#���3@��t���!?��2�-��@zUn6��ٿ+�z��@�#���3@��t���!?��2�-��@zUn6��ٿ+�z��@�#���3@��t���!?��2�-��@zUn6��ٿ+�z��@�#���3@��t���!?��2�-��@IS�3�ٿ��э�@�Y"��3@�FJ}ʐ!?��g��@IS�3�ٿ��э�@�Y"��3@�FJ}ʐ!?��g��@IS�3�ٿ��э�@�Y"��3@�FJ}ʐ!?��g��@��ٿ���S��@o{y3��3@�N�I��!?��$���@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@��wƢٿF%�}�Z�@l����3@3��f�!?��͆Q�@J��ћٿ�Sq����@Hķ��3@��K��!?�Q�0�@0NgԔٿ��!���@~�眴�3@Rm�q��!?�k�m�@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@���c�ٿE }�5��@l5�3@�BV�!?���U���@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@�K���ٿ���Ի�@a�!���3@�����!?�TJv��@���1��ٿj M�@���K�3@�G!$�!?fg$�p`�@���1��ٿj M�@���K�3@�G!$�!?fg$�p`�@���1��ٿj M�@���K�3@�G!$�!?fg$�p`�@���1��ٿj M�@���K�3@�G!$�!?fg$�p`�@���1��ٿj M�@���K�3@�G!$�!?fg$�p`�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@��t0�ٿ���mz��@1@-��3@5)��!?(i��H�@z��:$�ٿ�K�ޙ;�@��a*h�3@[-酐!?sv�l!��@z��:$�ٿ�K�ޙ;�@��a*h�3@[-酐!?sv�l!��@z��:$�ٿ�K�ޙ;�@��a*h�3@[-酐!?sv�l!��@z��:$�ٿ�K�ޙ;�@��a*h�3@[-酐!?sv�l!��@z��:$�ٿ�K�ޙ;�@��a*h�3@[-酐!?sv�l!��@i��n�ٿm�V�:�@6����3@:���!?*l�ťY�@i��n�ٿm�V�:�@6����3@:���!?*l�ťY�@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@/�ϴA�ٿ�}���|�@<�>-J�3@�;f�Ԑ!?������@#�2��ٿ�����@B5!
&�3@o�ҋ�!?'�y(�^�@#�2��ٿ�����@B5!
&�3@o�ҋ�!?'�y(�^�@Sp�D�ٿ�����@īfڪ�3@R!m>�!?"	ٲ�@Sp�D�ٿ�����@īfڪ�3@R!m>�!?"	ٲ�@s˕o�ٿY��ݥ�@��+��3@�T�`�!?����t�@s˕o�ٿY��ݥ�@��+��3@�T�`�!?����t�@s˕o�ٿY��ݥ�@��+��3@�T�`�!?����t�@s˕o�ٿY��ݥ�@��+��3@�T�`�!?����t�@�l��ٿ<��
SI�@��Ҝ��3@����!?�A�p��@�l��ٿ<��
SI�@��Ҝ��3@����!?�A�p��@�l��ٿ<��
SI�@��Ҝ��3@����!?�A�p��@�l��ٿ<��
SI�@��Ҝ��3@����!?�A�p��@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@�g�ǯ�ٿY8�z��@�C
n�3@�6ܐ!?��ii�@z�@f�ٿ(�R�@��� �3@e�YO��!?�E�?���@���,�ٿ�^��E�@�Q�I�3@f�ZW�!?sۓ����@���,�ٿ�^��E�@�Q�I�3@f�ZW�!?sۓ����@���,�ٿ�^��E�@�Q�I�3@f�ZW�!?sۓ����@���,�ٿ�^��E�@�Q�I�3@f�ZW�!?sۓ����@Ӌ<�8�ٿ���"���@,tw3��3@�1iS��!?Z3l���@K�L�ٿ�����@g<����3@��%��!?���R���@K�L�ٿ�����@g<����3@��%��!?���R���@K�L�ٿ�����@g<����3@��%��!?���R���@K�L�ٿ�����@g<����3@��%��!?���R���@K�L�ٿ�����@g<����3@��%��!?���R���@K�L�ٿ�����@g<����3@��%��!?���R���@;T���ٿ�цn2�@4Oc�V�3@}��X��!?,:$U���@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@씂��ٿ׳rդ�@�/}&��3@e�
��!?
B�(k>�@�l��F�ٿKR��@L���P�3@�H�G �!?��w�Ұ�@�l��F�ٿKR��@L���P�3@�H�G �!?��w�Ұ�@�l��F�ٿKR��@L���P�3@�H�G �!?��w�Ұ�@�?�ٿ$��mΊ�@���3@��L�!?���!��@�?�ٿ$��mΊ�@���3@��L�!?���!��@�?�ٿ$��mΊ�@���3@��L�!?���!��@�?�ٿ$��mΊ�@���3@��L�!?���!��@�?�ٿ$��mΊ�@���3@��L�!?���!��@�?�ٿ$��mΊ�@���3@��L�!?���!��@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@���A�ٿ���إ�@21�z��3@�Q3W��!?G�J�@B�u��ٿ��Y�h��@�ś�-�3@�֚��!?�Z���@B�u��ٿ��Y�h��@�ś�-�3@�֚��!?�Z���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�L����ٿ5r�K���@$ju)�3@�mD��!?|���@�l~Ԡٿ�k���s�@��y�W�3@��t���!?�����@�l~Ԡٿ�k���s�@��y�W�3@��t���!?�����@�l~Ԡٿ�k���s�@��y�W�3@��t���!?�����@�a b��ٿ��{�_��@Kܦi��3@!)��s�!?��w��@�a b��ٿ��{�_��@Kܦi��3@!)��s�!?��w��@�a b��ٿ��{�_��@Kܦi��3@!)��s�!?��w��@^�]�_�ٿ2�B ��@N*C*�3@a�ᗏ�!?�Bf�]��@+A�7��ٿr�&��@�B�^4�3@
1���!?MK-�Q�@+A�7��ٿr�&��@�B�^4�3@
1���!?MK-�Q�@3*���ٿ� �6��@�k!"�3@ܥ�Đ!?(/5����@�� ��ٿ�
4��@��?��3@9鉞�!?2U�%�S�@�� ��ٿ�
4��@��?��3@9鉞�!?2U�%�S�@�� ��ٿ�
4��@��?��3@9鉞�!?2U�%�S�@�� ��ٿ�
4��@��?��3@9鉞�!?2U�%�S�@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@���1��ٿMWv>ߤ�@
�����3@�/�l�!?g�v��@�����ٿ:d����@ɟ4���3@E~Оؐ!?�x�1��@�����ٿ:d����@ɟ4���3@E~Оؐ!?�x�1��@๧�٥ٿ���N| �@&���3@y�f�!?.�j7���@๧�٥ٿ���N| �@&���3@y�f�!?.�j7���@๧�٥ٿ���N| �@&���3@y�f�!?.�j7���@�о�s�ٿ�~�x{q�@S��(�3@�I����!?���(xB�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@x~�Gr�ٿ"��ՠ�@�|�&��3@9vK{��!?]�u�:T�@�{G'�ٿbRMp�@�g>ӊ�3@o.��А!?jAˡ#9�@�{G'�ٿbRMp�@�g>ӊ�3@o.��А!?jAˡ#9�@�{G'�ٿbRMp�@�g>ӊ�3@o.��А!?jAˡ#9�@�{G'�ٿbRMp�@�g>ӊ�3@o.��А!?jAˡ#9�@e1����ٿ�w3�D�@7Jq��3@19dN�!?�L5ID�@e1����ٿ�w3�D�@7Jq��3@19dN�!?�L5ID�@e1����ٿ�w3�D�@7Jq��3@19dN�!?�L5ID�@e1����ٿ�w3�D�@7Jq��3@19dN�!?�L5ID�@��w���ٿ������@��&8�3@2����!?|�Uk�V�@f�1�ҞٿK�/�qi�@�(����3@qipr�!?��O)j��@f�1�ҞٿK�/�qi�@�(����3@qipr�!?��O)j��@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@�m�x՛ٿvB�Wt�@Z�� �3@c��ċ�!?���{���@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@��˫^�ٿ$3���@�.u�?�3@�5��!?y�va��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@Os�.Z�ٿ5T����@�����3@mT��!?�)�"
��@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@CBj�ٿEK@�y"�@�v�_�3@�KƆ�!?�t���@�U!�ٿ�X��-�@������3@�b��!?���3j�@ְld?�ٿ��p���@��@��3@�����!?��<����@ְld?�ٿ��p���@��@��3@�����!?��<����@^ߎ�Q�ٿ���I�:�@�Vk�3@����͐!?���@V�~,�ٿ=7�j�@�D�cG�3@��_ΐ!?4��}o��@V�~,�ٿ=7�j�@�D�cG�3@��_ΐ!?4��}o��@V�~,�ٿ=7�j�@�D�cG�3@��_ΐ!?4��}o��@V�~,�ٿ=7�j�@�D�cG�3@��_ΐ!?4��}o��@V�~,�ٿ=7�j�@�D�cG�3@��_ΐ!?4��}o��@��W���ٿN,|�7g�@5�_���3@	jڛ��!?X�%8u��@��W���ٿN,|�7g�@5�_���3@	jڛ��!?X�%8u��@��W���ٿN,|�7g�@5�_���3@	jڛ��!?X�%8u��@��W���ٿN,|�7g�@5�_���3@	jڛ��!?X�%8u��@��W���ٿN,|�7g�@5�_���3@	jڛ��!?X�%8u��@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@d�!��ٿ˞�p�@h�EB�3@�\����!?l�U`�@��`w�ٿ�\���@���3@ޖ6I��!?h�~��@��`w�ٿ�\���@���3@ޖ6I��!?h�~��@��`w�ٿ�\���@���3@ޖ6I��!?h�~��@���뾧ٿ)��I�K�@HAht�3@�3 �!?Md���@���뾧ٿ)��I�K�@HAht�3@�3 �!?Md���@���뾧ٿ)��I�K�@HAht�3@�3 �!?Md���@���뾧ٿ)��I�K�@HAht�3@�3 �!?Md���@��y+�ٿm�I>��@��0lu�3@&���̐!?�̄+nB�@��y+�ٿm�I>��@��0lu�3@&���̐!?�̄+nB�@��y+�ٿm�I>��@��0lu�3@&���̐!?�̄+nB�@i�<���ٿ�!�{�@�pĽ�3@3���!?X�]uH��@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@V�*LB�ٿ��?6P�@m}a��3@�Q�~��!?hU�*�@�_්�ٿ�._ZU�@�B���3@z��!?,��&� �@�_්�ٿ�._ZU�@�B���3@z��!?,��&� �@�_්�ٿ�._ZU�@�B���3@z��!?,��&� �@F�,]�ٿW`*�@S/)�3@�����!?RA��B��@F�,]�ٿW`*�@S/)�3@�����!?RA��B��@F�,]�ٿW`*�@S/)�3@�����!?RA��B��@~ժ��ٿ�H#A��@QI�8��3@l2 �ː!?ܣ����@\BN"p�ٿR� �ǯ�@��|�3@"#V�!?��dU���@�/S�Ʀٿyb�K-�@�2���3@����Ɛ!?7��7��@�/S�Ʀٿyb�K-�@�2���3@����Ɛ!?7��7��@�2�\��ٿ�
���@J����3@:����!?�	�PZ�@�2�\��ٿ�
���@J����3@:����!?�	�PZ�@p|hl�ٿ��g n��@�
2x�3@B�ϐ!? �2O�@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�SQv�ٿ&nV2T��@�K�2��3@�e�Ȑ!?>!Dw��@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@�R���ٿ���U��@#-�q�3@|xS��!?� 6��|�@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@R(T�˟ٿr6�1H@�@�P����3@V����!?�'Y���@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�Ҋ��ٿ/�K8�@�[��3@l*e�Đ!?�����@�ܩG��ٿݢ�"�@9X*��3@j�ː!?���N�@�ܩG��ٿݢ�"�@9X*��3@j�ː!?���N�@�ܩG��ٿݢ�"�@9X*��3@j�ː!?���N�@�ܩG��ٿݢ�"�@9X*��3@j�ː!?���N�@�ܩG��ٿݢ�"�@9X*��3@j�ː!?���N�@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�Z�Cm�ٿ�ل��@%�/J��3@J��nِ!?�:C�]��@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�B;���ٿoԾ����@D�����3@���ڔ�!?�(yS�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@�MG��ٿ���!c�@�E���3@O��ړ�!?.�k�X�@+ϒ2�ٿ��j���@��~��3@]c�J��!?6R
އ��@+ϒ2�ٿ��j���@��~��3@]c�J��!?6R
އ��@+ϒ2�ٿ��j���@��~��3@]c�J��!?6R
އ��@b
�KV�ٿf_|&�t�@�k�m�3@�D�Ɛ!?|#�f��@b
�KV�ٿf_|&�t�@�k�m�3@�D�Ɛ!?|#�f��@���Y2�ٿ-:@P���@���3@O��0��!?���K��@:��h�ٿ֘W*���@�_��3@p/T��!?n*^=���@:��h�ٿ֘W*���@�_��3@p/T��!?n*^=���@8��V͟ٿ��K�;\�@��UN�3@�Ⱥ��!?��t�Q�@8��V͟ٿ��K�;\�@��UN�3@�Ⱥ��!?��t�Q�@8��V͟ٿ��K�;\�@��UN�3@�Ⱥ��!?��t�Q�@q����ٿ��>��@먰��3@p�YJߐ!?�g���@q����ٿ��>��@먰��3@p�YJߐ!?�g���@q����ٿ��>��@먰��3@p�YJߐ!?�g���@q����ٿ��>��@먰��3@p�YJߐ!?�g���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@����K�ٿ��8'��@��K;��3@����!?�!-���@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@5nW�/�ٿf����@�ɤ#��3@CW���!?����S��@'� ���ٿ*��nj�@dP���3@E3���!?nK}3@��@v"|�ٿDk��'�@s�+��3@��Ρ��!?���Ùc�@v"|�ٿDk��'�@s�+��3@��Ρ��!?���Ùc�@v"|�ٿDk��'�@s�+��3@��Ρ��!?���Ùc�@v"|�ٿDk��'�@s�+��3@��Ρ��!?���Ùc�@v"|�ٿDk��'�@s�+��3@��Ρ��!?���Ùc�@b��A��ٿ���}�@�W&���3@W
��!?	����@Q���ٿ|jDȎ�@T���3@��B!x�!?'��@���@Q���ٿ|jDȎ�@T���3@��B!x�!?'��@���@Q���ٿ|jDȎ�@T���3@��B!x�!?'��@���@Q���ٿ|jDȎ�@T���3@��B!x�!?'��@���@'�wx�ٿ�#a�h��@V�=y�3@�jM��!?�4P��@'�wx�ٿ�#a�h��@V�=y�3@�jM��!?�4P��@�9�ߟٿfcn���@kd�:(�3@E@e���!?[����P�@��2�,�ٿ��K���@eh���3@�?�Y�!?2������@��2�,�ٿ��K���@eh���3@�?�Y�!?2������@��2�,�ٿ��K���@eh���3@�?�Y�!?2������@��2�,�ٿ��K���@eh���3@�?�Y�!?2������@��2�,�ٿ��K���@eh���3@�?�Y�!?2������@ٺ>�F�ٿc!h�r�@�����3@����̐!?%z��F�@ٺ>�F�ٿc!h�r�@�����3@����̐!?%z��F�@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@톙S@�ٿ������@�՘���3@\0kĸ�!?n�����@Ԁ�6�ٿ��2���@��1���3@n�7��!?���Ė�@Ԁ�6�ٿ��2���@��1���3@n�7��!?���Ė�@Ԁ�6�ٿ��2���@��1���3@n�7��!?���Ė�@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@���ƞٿ���":��@��QT��3@�+��!?W�wo��@;����ٿͦ�(��@�>K�J�3@XN��!? hǳ;a�@;����ٿͦ�(��@�>K�J�3@XN��!? hǳ;a�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@W�?�МٿJ͘#&��@�3�� �3@�7���!?	��_x�@Zm�1ȡٿ3��f��@�ky|��3@� �S�!?�M}N���@K����ٿt�bM��@�l����3@���ː!?Y/Ƅ8��@K����ٿt�bM��@�l����3@���ː!?Y/Ƅ8��@����/�ٿ20�kɣ�@�>��3@`^"�!?�+���@�Ex�ٿE]E��@s)��3@�DD��!?�x�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@���}��ٿjՖ�)�@/B Z�3@��\�!?�3�����@K["���ٿ�:�/7�@4�-�3@c�h��!?��_)-�@K["���ٿ�:�/7�@4�-�3@c�h��!?��_)-�@K["���ٿ�:�/7�@4�-�3@c�h��!?��_)-�@K["���ٿ�:�/7�@4�-�3@c�h��!?��_)-�@�W����ٿ����@��p��3@�,ss��!?�1���@�W����ٿ����@��p��3@�,ss��!?�1���@�W����ٿ����@��p��3@�,ss��!?�1���@�W����ٿ����@��p��3@�,ss��!?�1���@����9�ٿh��W�@ꎏOk�3@WE�A��!?��` ���@����9�ٿh��W�@ꎏOk�3@WE�A��!?��` ���@����9�ٿh��W�@ꎏOk�3@WE�A��!?��` ���@����9�ٿh��W�@ꎏOk�3@WE�A��!?��` ���@��`4۝ٿ��q�P�@+��:��3@�6���!?g�iBO@�@��`4۝ٿ��q�P�@+��:��3@�6���!?g�iBO@�@��`4۝ٿ��q�P�@+��:��3@�6���!?g�iBO@�@��`4۝ٿ��q�P�@+��:��3@�6���!?g�iBO@�@��`4۝ٿ��q�P�@+��:��3@�6���!?g�iBO@�@��/��ٿ�"��:�@~o�"��3@�|M���!?2S�Z��@��/��ٿ�"��:�@~o�"��3@�|M���!?2S�Z��@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�ڬ���ٿq���i��@%JdU��3@[_4*ǐ!?!|��Q�@�U����ٿk�"���@lȡ8��3@�]�ῐ!?N!i�~�@��`V�ٿ:�Q���@���cJ 4@����!?1�f}��@��`V�ٿ:�Q���@���cJ 4@����!?1�f}��@��`V�ٿ:�Q���@���cJ 4@����!?1�f}��@��`V�ٿ:�Q���@���cJ 4@����!?1�f}��@��`V�ٿ:�Q���@���cJ 4@����!?1�f}��@�IlUC�ٿ���n�@QO(6��3@��q���!?^���E�@�IlUC�ٿ���n�@QO(6��3@��q���!?^���E�@�IlUC�ٿ���n�@QO(6��3@��q���!?^���E�@�IlUC�ٿ���n�@QO(6��3@��q���!?^���E�@G}HX��ٿH�&�܊�@"�׋��3@a�����!?�l�)�d�@G}HX��ٿH�&�܊�@"�׋��3@a�����!?�l�)�d�@G}HX��ٿH�&�܊�@"�׋��3@a�����!?�l�)�d�@W1��ٿ�;˚�@��do�3@�~�]��!?����^r�@W1��ٿ�;˚�@��do�3@�~�]��!?����^r�@W1��ٿ�;˚�@��do�3@�~�]��!?����^r�@W1��ٿ�;˚�@��do�3@�~�]��!?����^r�@W1��ٿ�;˚�@��do�3@�~�]��!?����^r�@=�l�àٿV�+C`�@��n��3@~;H$Ӑ!?����2��@=�l�àٿV�+C`�@��n��3@~;H$Ӑ!?����2��@.����ٿH"6)M�@td��3@z�:��!?l�!F�d�@S~�/�ٿݏA��@�Jr*��3@҇,�!?w}v�e��@S~�/�ٿݏA��@�Jr*��3@҇,�!?w}v�e��@S~�/�ٿݏA��@�Jr*��3@҇,�!?w}v�e��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@]����ٿI	G�\Q�@^4}��3@m5ǐ!?j��J"��@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@)�l'�ٿ��n��@x�'���3@]bu���!?���6;0�@|�XY�ٿ fc�r��@���3@7��W�!?�*	_��@�����ٿ��V@
P�@]�֚G�3@�b[Ȑ!?m�P�@s�#�̜ٿ���bc�@G	0n#�3@�G�5��!?��ʦ��@s�#�̜ٿ���bc�@G	0n#�3@�G�5��!?��ʦ��@s�#�̜ٿ���bc�@G	0n#�3@�G�5��!?��ʦ��@���2�ٿ��^��@�'*�3@�H3̐!?�Ʉq=)�@�����ٿ���_���@���3@��u��!?��P ��@xh�I�ٿ�=�xT��@�Yk�d�3@�=�`��!?}�v�$�@�#���ٿuM���@�T���3@�a�H��!?�q�U70�@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@���!��ٿ�	���@ܨ�C��3@:h{5v�!?��*0��@D2#�ٿ����{�@E8�t�3@����!?�.�רd�@D2#�ٿ����{�@E8�t�3@����!?�.�רd�@��.L�ٿ2L��M��@��yb�3@t��;�!?����'�@��.L�ٿ2L��M��@��yb�3@t��;�!?����'�@�����ٿ+���@�+���3@f�`��!?yt3[��@�����ٿ+���@�+���3@f�`��!?yt3[��@�����ٿ+���@�+���3@f�`��!?yt3[��@�����ٿ+���@�+���3@f�`��!?yt3[��@�����ٿ+���@�+���3@f�`��!?yt3[��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@�0n՗ٿ�pR �~�@�ݽ�x�3@��!��!?k*��@AO,Mg�ٿ��r��@L���3@W�Đ!?o49M���@AO,Mg�ٿ��r��@L���3@W�Đ!?o49M���@AO,Mg�ٿ��r��@L���3@W�Đ!?o49M���@sA�v�ٿ&LUYC��@�����3@�B�E��!?�����@�Ѐɪ�ٿR��	���@#ZO��3@Y�Id�!?c���6�@�Ѐɪ�ٿR��	���@#ZO��3@Y�Id�!?c���6�@C{�vP�ٿ=G��_�@�zZ}�3@����!?�E����@C{�vP�ٿ=G��_�@�zZ}�3@����!?�E����@C{�vP�ٿ=G��_�@�zZ}�3@����!?�E����@C{�vP�ٿ=G��_�@�zZ}�3@����!?�E����@���뜢ٿV��0��@&_�I��3@h{P��!?ݵ�z9^�@���뜢ٿV��0��@&_�I��3@h{P��!?ݵ�z9^�@���뜢ٿV��0��@&_�I��3@h{P��!?ݵ�z9^�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�$]h�ٿ^fGI1��@�sN�4@V3[ː!?��9��V�@�P	W�ٿA��'*�@�^Ÿ�3@��:)��!?�!�'��@�P	W�ٿA��'*�@�^Ÿ�3@��:)��!?�!�'��@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@�pp���ٿ"`��c�@B'!���3@*�Hx��!?�ѵ\�@��U(��ٿ5E���@)~��3@s�L��!?o��o��@��U(��ٿ5E���@)~��3@s�L��!?o��o��@�d.�h�ٿm7�����@��<j�3@�JT���!?��\OM�@�d.�h�ٿm7�����@��<j�3@�JT���!?��\OM�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@x*1�ٿ����+ �@#�Q��3@��x笐!?�sq�Sy�@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@���ٿ Y�����@�/H��3@Y�Z✐!?/���<��@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@y���ٿ��c?]��@�r���3@pH��Ɛ!?7\i���@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@h ZW�ٿʔ3�W�@�� ��3@� 0P�!?nC;#��@���Tǝٿ z6�C��@}�pt]�3@c�68��!?z��z�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@��wﮘٿ�8�5���@:�Mp(�3@�6 ʃ�!?��p�
�@���%�ٿ�G-G~�@�͍��3@��R|�!?��T���@���%�ٿ�G-G~�@�͍��3@��R|�!?��T���@���%�ٿ�G-G~�@�͍��3@��R|�!?��T���@�>Ϸ�ٿ�qR���@�$zO��3@�Á�>�!?��t�<N�@�>Ϸ�ٿ�qR���@�$zO��3@�Á�>�!?��t�<N�@�>Ϸ�ٿ�qR���@�$zO��3@�Á�>�!?��t�<N�@�:�Z؝ٿ�z���@:|^���3@�,@.ې!?9u�2���@"��v��ٿ�$|�>�@�����3@�jj��!?`��V��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@�� ��ٿ^�m����@E�ƥ��3@�ѱ<�!?�HW@��@��)�ٿ���?r�@[Z��3@N�S�!?)��^��@�)��ԡٿ;��z\�@;S���3@ɾ���!?�u W��@�)��ԡٿ;��z\�@;S���3@ɾ���!?�u W��@�)��ԡٿ;��z\�@;S���3@ɾ���!?�u W��@͜�ٿZ ��+b�@�y��3@�U�ސ!?�)�Jo��@͜�ٿZ ��+b�@�y��3@�U�ސ!?�)�Jo��@͜�ٿZ ��+b�@�y��3@�U�ސ!?�)�Jo��@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@���q�ٿL�)""�@C�����3@��t#А!?����w�@d%󼰥ٿ�o�Зb�@����2�3@ն�!?��z��@��$S�ٿ�����@DDVh�3@�B�!?&,�g-�@<��ٿd/t/�@������3@1}�X��!?	�6�9�@R���x�ٿ��
i��@,�Ɏ�3@?�kd�!?U� c���@R���x�ٿ��
i��@,�Ɏ�3@?�kd�!?U� c���@I�{��ٿ}��7�@�+��3@�*����!?�N3��Z�@������ٿ]�)v���@����3@ﶻ�!?"%-�6$�@if�ٿ�������@ ��_H�3@�Nnʐ!??¥	K��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@h1B�r�ٿO���|��@�5ʷo�3@���~�!?��{��@U�s�ٿU�?Ȃ�@�3-��3@ҍJ�ߐ!?�sh2��@Kt�]l�ٿ�K��%��@���.[�3@|ߘt�!?Z��ؽ-�@Kt�]l�ٿ�K��%��@���.[�3@|ߘt�!?Z��ؽ-�@�#�)�ٿ��y��@�E��u�3@9awh�!?PcD.!��@�#�)�ٿ��y��@�E��u�3@9awh�!?PcD.!��@�#�)�ٿ��y��@�E��u�3@9awh�!?PcD.!��@�	�KўٿP��C0��@Þ�3@1n���!? hU���@��C�ٿ?���@�{�e�3@%j#��!?���.�@��C�ٿ?���@�{�e�3@%j#��!?���.�@��C�ٿ?���@�{�e�3@%j#��!?���.�@��C�ٿ?���@�{�e�3@%j#��!?���.�@2!�%-�ٿ%?�����@%�<��3@�9gn�!?v�h����@2!�%-�ٿ%?�����@%�<��3@�9gn�!?v�h����@:�����ٿ�g�5��@ӞHE�3@ �0��!?��M��@�@:�����ٿ�g�5��@ӞHE�3@ �0��!?��M��@�@:�����ٿ�g�5��@ӞHE�3@ �0��!?��M��@�@:�����ٿ�g�5��@ӞHE�3@ �0��!?��M��@�@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@�,�i̥ٿ�Z?YU��@)e��3@ƨ'\��!?l�}A���@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@I�c�ٿdd�����@��2�3@�K�Ѐ�!?#؜{~��@X��ٿ*ʔZ�i�@'ô_��3@"��A��!?"��:���@X��ٿ*ʔZ�i�@'ô_��3@"��A��!?"��:���@X��ٿ*ʔZ�i�@'ô_��3@"��A��!?"��:���@X��ٿ*ʔZ�i�@'ô_��3@"��A��!?"��:���@`=�{�ٿ�P#ր��@��M/F�3@�+ᐐ!?_z�&��@`=�{�ٿ�P#ր��@��M/F�3@�+ᐐ!?_z�&��@0z:O~�ٿ���u8�@�	k��3@L�����!?竈h��@0z:O~�ٿ���u8�@�	k��3@L�����!?竈h��@����n�ٿ�?L�@��\M�3@ b$���!? 95�8�@����n�ٿ�?L�@��\M�3@ b$���!? 95�8�@A#�eM�ٿ8�|a��@��
\��3@��
�!?��#- �@A#�eM�ٿ8�|a��@��
\��3@��
�!?��#- �@A#�eM�ٿ8�|a��@��
\��3@��
�!?��#- �@�xϝQ�ٿ�θ��{�@H6R+�3@��o��!?4'c�Te�@�xϝQ�ٿ�θ��{�@H6R+�3@��o��!?4'c�Te�@�xϝQ�ٿ�θ��{�@H6R+�3@��o��!?4'c�Te�@�xϝQ�ٿ�θ��{�@H6R+�3@��o��!?4'c�Te�@z���ٿf�t"��@�ܤ���3@�y��%�!?� �5�3�@rX����ٿ�{���@��E���3@߆����!?�҂���@rX����ٿ�{���@��E���3@߆����!?�҂���@���0�ٿ�um�]��@:��U��3@J��h��!?�0Vs�l�@���0�ٿ�um�]��@:��U��3@J��h��!?�0Vs�l�@�y\w�ٿ�2�3���@sd�:��3@@C��!?�Q+l���@�y\w�ٿ�2�3���@sd�:��3@@C��!?�Q+l���@�y\w�ٿ�2�3���@sd�:��3@@C��!?�Q+l���@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@�y�5+�ٿ�ܘ�@�P#�3@侀�ؐ!?���w��@��q�p�ٿ��6G�@G*�!��3@5&���!?�Ec��@��q�p�ٿ��6G�@G*�!��3@5&���!?�Ec��@��q�p�ٿ��6G�@G*�!��3@5&���!?�Ec��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@v��� �ٿ�!�7��@��8�/�3@��ul�!?�>#=v��@��X��ٿ���� Y�@�*y��3@�)	�!?�꫐��@��X��ٿ���� Y�@�*y��3@�)	�!?�꫐��@?w&:�ٿ����E�@�n<b�3@.W��s�!?og\���@��z� �ٿ É�T�@�����3@����!?��L���@��z� �ٿ É�T�@�����3@����!?��L���@��z� �ٿ É�T�@�����3@����!?��L���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@&�ٯ��ٿV�RU���@����3@��l��!?[�E���@/�3��ٿ�9j��@�<L)��3@�����!?P|��d�@/�3��ٿ�9j��@�<L)��3@�����!?P|��d�@��G�ٿL(�^U	�@�.?���3@��!��!?�t7���@�����ٿ�MŸ��@}�<;��3@�ˇ6�!?��,�7�@��EK��ٿ=MP�
��@�����3@,���Đ!?E�t�
 �@��EK��ٿ=MP�
��@�����3@,���Đ!?E�t�
 �@��EK��ٿ=MP�
��@�����3@,���Đ!?E�t�
 �@��EK��ٿ=MP�
��@�����3@,���Đ!?E�t�
 �@��EK��ٿ=MP�
��@�����3@,���Đ!?E�t�
 �@�]��ٿ���>f��@�|^�D�3@��O/��!?:�q\��@�]��ٿ���>f��@�|^�D�3@��O/��!?:�q\��@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@}/#o�ٿ�#6��@�H�4(�3@䝜���!?ד�&�V�@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+'z�E�ٿ�_�����@�?�C7�3@�!�&o�!?�m�����@+��C�ٿt�Q��@{9�F��3@E����!?��%�Q�@+��C�ٿt�Q��@{9�F��3@E����!?��%�Q�@+��C�ٿt�Q��@{9�F��3@E����!?��%�Q�@^vZ��ٿ���.��@����3@��/ߐ!?�3�ghM�@��`�ٿ��5d�@��7M�3@�I҄�!?8lHeV��@��`�ٿ��5d�@��7M�3@�I҄�!?8lHeV��@'x�W��ٿ������@�ՠ��3@�	S�!?;�6 ^_�@'x�W��ٿ������@�ՠ��3@�	S�!?;�6 ^_�@O�D��ٿFT��t�@�+q�3@�5���!?~�^NaB�@O�D��ٿFT��t�@�+q�3@�5���!?~�^NaB�@O�D��ٿFT��t�@�+q�3@�5���!?~�^NaB�@c�dƢٿ���8N��@1K�Q��3@�٢��!?��F��@c�dƢٿ���8N��@1K�Q��3@�٢��!?��F��@c�dƢٿ���8N��@1K�Q��3@�٢��!?��F��@c�dƢٿ���8N��@1K�Q��3@�٢��!?��F��@���)�ٿf���:�@������3@�*�;��!?SC� ���@���)�ٿf���:�@������3@�*�;��!?SC� ���@���)�ٿf���:�@������3@�*�;��!?SC� ���@���)�ٿf���:�@������3@�*�;��!?SC� ���@�]�Y�ٿ�� �~�@�����3@j���ϐ!?��D���@�]�Y�ٿ�� �~�@�����3@j���ϐ!?��D���@������ٿ�j����@we}���3@��l��!?����@������ٿ�j����@we}���3@��l��!?����@������ٿ�j����@we}���3@��l��!?����@������ٿ�j����@we}���3@��l��!?����@�C	_G�ٿ������@�1��3@T}L��!?�|���@�C	_G�ٿ������@�1��3@T}L��!?�|���@�C	_G�ٿ������@�1��3@T}L��!?�|���@�C	_G�ٿ������@�1��3@T}L��!?�|���@�C	_G�ٿ������@�1��3@T}L��!?�|���@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@���|�ٿ�I���`�@̠ã�3@�� &ΐ!?q�cc��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�с[�ٿ����� �@�r�3@	��!?-�R��@�y��ٿJc	eO�@z�9�L�3@�/���!?�i�}w�@�H~�*�ٿ�Re^K\�@��U�h�3@��}���!?n���U��@�H~�*�ٿ�Re^K\�@��U�h�3@��}���!?n���U��@�H~�*�ٿ�Re^K\�@��U�h�3@��}���!?n���U��@�H~�*�ٿ�Re^K\�@��U�h�3@��}���!?n���U��@�H~�*�ٿ�Re^K\�@��U�h�3@��}���!?n���U��@���~�ٿv���;��@aӺ4��3@ڣ�H��!?"7-aM�@���~�ٿv���;��@aӺ4��3@ڣ�H��!?"7-aM�@���~�ٿv���;��@aӺ4��3@ڣ�H��!?"7-aM�@���~�ٿv���;��@aӺ4��3@ڣ�H��!?"7-aM�@4!��s�ٿJT����@����y�3@q~6���!?c�5r1��@4!��s�ٿJT����@����y�3@q~6���!?c�5r1��@4!��s�ٿJT����@����y�3@q~6���!?c�5r1��@4!��s�ٿJT����@����y�3@q~6���!?c�5r1��@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@��lL�ٿ5籹�r�@��L�1�3@C���!?��}�zU�@���z�ٿ±.���@:�v��3@[�����!?�މ
`��@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@�)s�ɟٿ1 �+L��@z�8F�3@��l���!?���� 5�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@����ٿJ��]�@V3����3@��!?MFQ�<�@? 5K�ٿ��=�*��@8�6�3@���ΐ!?i��=t�@? 5K�ٿ��=�*��@8�6�3@���ΐ!?i��=t�@#N��]�ٿ'��Po��@�A�4�3@Y��W��!?�^�\�^�@#N��]�ٿ'��Po��@�A�4�3@Y��W��!?�^�\�^�@#N��]�ٿ'��Po��@�A�4�3@Y��W��!?�^�\�^�@#N��]�ٿ'��Po��@�A�4�3@Y��W��!?�^�\�^�@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@�E�q�ٿ��Y���@޴E���3@s��t��!?BA����@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@���K�ٿG��C��@t�;�x�3@��5̆�!?������@�K�̦ٿd�7�}}�@t'Ϟ��3@�٤x�!?���� �@^;�j�ٿ�`u���@_�j�G�3@�Y#X�!?L{#�L��@�A�ĝٿ�&u	���@~�/��3@�<�3�!?�ԣZk�@�A�ĝٿ�&u	���@~�/��3@�<�3�!?�ԣZk�@�A�ĝٿ�&u	���@~�/��3@�<�3�!?�ԣZk�@�r@CR�ٿ���I��@]E����3@�ʉ���!?mc㧀��@�r@CR�ٿ���I��@]E����3@�ʉ���!?mc㧀��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@0eh�a�ٿ��+.+ �@�����3@�nIѐ!?�f��J��@@7���ٿP� L��@����3@��ڡ�!?bC 1TB�@@7���ٿP� L��@����3@��ڡ�!?bC 1TB�@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@4�;D�ٿ�Z�݅N�@9d�v��3@!Q�(��!?��r���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ٿ��wZ,�@������3@R�a���!?N2���@���ˆ�ٿD�b0�@�{���3@�u[�}�!?�L�Y&�@���ˆ�ٿD�b0�@�{���3@�u[�}�!?�L�Y&�@��L�j�ٿ�6��G��@�	����3@�́�!?AvkY�@�.Y��ٿ���c�@{�*�8�3@��A��!?�6*Rn��@�.Y��ٿ���c�@{�*�8�3@��A��!?�6*Rn��@�.Y��ٿ���c�@{�*�8�3@��A��!?�6*Rn��@�.Y��ٿ���c�@{�*�8�3@��A��!?�6*Rn��@�.Y��ٿ���c�@{�*�8�3@��A��!?�6*Rn��@�4S�ٿR��y�@Hj�t��3@:%�А!?{�*���@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@-�a��ٿ>ey��9�@v�kQr�3@�X���!?ڀ"�N�@Ne ���ٿ�^�����@�ɯ&��3@���AҐ!?�5����@Ne ���ٿ�^�����@�ɯ&��3@���AҐ!?�5����@Ne ���ٿ�^�����@�ɯ&��3@���AҐ!?�5����@Ne ���ٿ�^�����@�ɯ&��3@���AҐ!?�5����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@�&|��ٿ�\+��P�@7m�Y��3@���!?�h����@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@DU�f�ٿm���K@�@�;�3@�Ң[�!?|(> �%�@�S؜�ٿ���{g�@Eߓ��3@��&�x�!?H�a۪;�@�S؜�ٿ���{g�@Eߓ��3@��&�x�!?H�a۪;�@�S؜�ٿ���{g�@Eߓ��3@��&�x�!?H�a۪;�@�s�W��ٿ^!�����@��G��3@����U�!?<�$Bt�@�4W5��ٿ�f�mH�@4ژ6�3@߈E=d�!?!3$�Z%�@�4W5��ٿ�f�mH�@4ژ6�3@߈E=d�!?!3$�Z%�@�4W5��ٿ�f�mH�@4ژ6�3@߈E=d�!?!3$�Z%�@.�qũٿ�ݤ*$s�@��<���3@r���!?��}�N�@�$�	��ٿ4�K���@Y�����3@;z;֐!?�1nɺ{�@�$�	��ٿ4�K���@Y�����3@;z;֐!?�1nɺ{�@a��ٿ�lh�6�@1���R�3@� �%�!?�e}+Y�@o�X}�ٿ��:�� �@�*L^�3@��O��!?���yb�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@�H�eĠٿV�]�y��@fw����3@�J��!?����}�@i�2ʢٿ��eQ�@ow�Q�3@�	�X͐!?���0^�@���^�ٿ�@�O�@�k�Ϸ�3@ d��!?������@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@[����ٿ�)�Ob�@������3@� �!?��f�Y��@6^�P��ٿt���P�@o�u���3@������!?x��t��@6^�P��ٿt���P�@o�u���3@������!?x��t��@6^�P��ٿt���P�@o�u���3@������!?x��t��@6^�P��ٿt���P�@o�u���3@������!?x��t��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@j���ٿ�����@�����3@#�܌��!?V�c�&��@�:��5�ٿ�C�_a�@�a����3@s𘞹�!?�F����@�:��5�ٿ�C�_a�@�a����3@s𘞹�!?�F����@�:��5�ٿ�C�_a�@�a����3@s𘞹�!?�F����@|�D��ٿ{������@�2��3@��t�!?���q�$�@|�D��ٿ{������@�2��3@��t�!?���q�$�@|�D��ٿ{������@�2��3@��t�!?���q�$�@|�D��ٿ{������@�2��3@��t�!?���q�$�@|�D��ٿ{������@�2��3@��t�!?���q�$�@;�l�l�ٿ��"x�?�@W�QM�3@f�Q�!?u�n^x��@��q���ٿ������@�[����3@�9M���!?�%X�WA�@��q���ٿ������@�[����3@�9M���!?�%X�WA�@���OP�ٿ�4Ѳ�k�@4W���3@�+�,{�!?�'�N��@��[p�ٿ��C�+��@W��34�3@Kr��^�!?�����@�6$03�ٿ�o���@�;�K��3@�,��h�!?����>u�@�6$03�ٿ�o���@�;�K��3@�,��h�!?����>u�@uӶ$��ٿ��B&j�@��3��3@!❜��!?���:���@����*�ٿ�a�S1�@���+��3@��#Q��!?�+��@Q8�_�ٿ��H�|�@9*{K��3@g���!?�7�w&�@Q8�_�ٿ��H�|�@9*{K��3@g���!?�7�w&�@Q8�_�ٿ��H�|�@9*{K��3@g���!?�7�w&�@Q8�_�ٿ��H�|�@9*{K��3@g���!?�7�w&�@�>E��ٿ*�a�
��@��;�3@��;�ߐ!?N�J�h�@�>E��ٿ*�a�
��@��;�3@��;�ߐ!?N�J�h�@�����ٿ�qᕊ�@io�3@�m6��!?q�J�
�@�����ٿ�qᕊ�@io�3@�m6��!?q�J�
�@�����ٿ�qᕊ�@io�3@�m6��!?q�J�
�@e2�E��ٿ%�t���@(y*{��3@eiP<��!?�.73b��@e2�E��ٿ%�t���@(y*{��3@eiP<��!?�.73b��@e2�E��ٿ%�t���@(y*{��3@eiP<��!?�.73b��@Ǻ V�ٿ`bP�ox�@����3@�:	А!?dNz_���@Ǻ V�ٿ`bP�ox�@����3@�:	А!?dNz_���@Ǻ V�ٿ`bP�ox�@����3@�:	А!?dNz_���@eC��ݞٿq�`E��@�6CI��3@�I#!?����,��@eC��ݞٿq�`E��@�6CI��3@�I#!?����,��@5��ٿ���\��@PxGTt�3@l7��Ґ!?ѹ�̖��@5��ٿ���\��@PxGTt�3@l7��Ґ!?ѹ�̖��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@���d��ٿ��y�+7�@N�����3@b��`Ɛ!?���7��@�߄��ٿY��9���@�d�!�3@LU�l�!?�n(����@�߄��ٿY��9���@�d�!�3@LU�l�!?�n(����@�߄��ٿY��9���@�d�!�3@LU�l�!?�n(����@�߄��ٿY��9���@�d�!�3@LU�l�!?�n(����@��g�{�ٿĭl�;�@��~��3@�7�Kː!?���z���@��g�{�ٿĭl�;�@��~��3@�7�Kː!?���z���@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@�k*���ٿ%��	�#�@�.���3@}E�ꇐ!?�A�D��@����ٿ�ZSE4l�@���
�3@��Ϻ��!?"K5���@l3�z�ٿ-ӽ'!�@�2�0�3@`Dx���!?���Vj�@l3�z�ٿ-ӽ'!�@�2�0�3@`Dx���!?���Vj�@l3�z�ٿ-ӽ'!�@�2�0�3@`Dx���!?���Vj�@T���؜ٿ�_��C�@����3@я����!? )s³��@�,��ʞٿ�Zp0���@���T�3@�XQ���!?p���K�@�,��ʞٿ�Zp0���@���T�3@�XQ���!?p���K�@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@M�0��ٿ3����b�@y�Ť)�3@����!?��ڢ��@������ٿ����@�����3@���Pϐ!?rF��]*�@������ٿ����@�����3@���Pϐ!?rF��]*�@������ٿ����@�����3@���Pϐ!?rF��]*�@������ٿ����@�����3@���Pϐ!?rF��]*�@������ٿ����@�����3@���Pϐ!?rF��]*�@������ٿ����@�����3@���Pϐ!?rF��]*�@J�[L[�ٿ �@�-�@Lψe��3@m+��!?���.��@J�[L[�ٿ �@�-�@Lψe��3@m+��!?���.��@J�[L[�ٿ �@�-�@Lψe��3@m+��!?���.��@J�[L[�ٿ �@�-�@Lψe��3@m+��!?���.��@J�[L[�ٿ �@�-�@Lψe��3@m+��!?���.��@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@y)��ҥٿ�UD�+^�@K)Z��3@�o��ϐ!?}������@���*g�ٿ��6�}�@��2Q�3@ݿ����!?�D����@z�E�$�ٿ��Α,�@������3@U-�b��!?
9�I��@z�E�$�ٿ��Α,�@������3@U-�b��!?
9�I��@z�E�$�ٿ��Α,�@������3@U-�b��!?
9�I��@�J槧ٿ�3!�K�@b�4� �3@�͘:��!?Y2t��@�bQ���ٿ�����B�@���,<�3@�hk��!?K��aZ�@�bQ���ٿ�����B�@���,<�3@�hk��!?K��aZ�@�bQ���ٿ�����B�@���,<�3@�hk��!?K��aZ�@WF�ٿ�tP��@q��3�3@�[����!?���Wt��@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��E8�ٿpe�o���@���Q��3@=W��!?�JFWh
�@��u�Οٿ���$N�@j���[�3@#N3��!?�i��J��@��u�Οٿ���$N�@j���[�3@#N3��!?�i��J��@��u�Οٿ���$N�@j���[�3@#N3��!?�i��J��@4�v���ٿ;�����@�c3���3@Whb�!?���Er��@4�v���ٿ;�����@�c3���3@Whb�!?���Er��@4�v���ٿ;�����@�c3���3@Whb�!?���Er��@4�v���ٿ;�����@�c3���3@Whb�!?���Er��@4�v���ٿ;�����@�c3���3@Whb�!?���Er��@΅Z\��ٿ_�BlT'�@���A�3@�����!?�����@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@AB"�1�ٿ\��I]	�@r�G?��3@�x乐!? |��N�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@Z6���ٿ�27 ��@:S�g�3@���!?Wą6e�@�}�H�ٿk�){#�@Eʭ�3@הV��!?���J���@�}�H�ٿk�){#�@Eʭ�3@הV��!?���J���@��Ce�ٿ�/l� ��@ayL�J�3@���М�!?�������@��.?�ٿz<J}\�@fx^[�3@�8U��!?�`U�R�@��.?�ٿz<J}\�@fx^[�3@�8U��!?�`U�R�@��.?�ٿz<J}\�@fx^[�3@�8U��!?�`U�R�@lDU�W�ٿpS����@��Z���3@�q���!?�.�����@lDU�W�ٿpS����@��Z���3@�q���!?�.�����@lDU�W�ٿpS����@��Z���3@�q���!?�.�����@lDU�W�ٿpS����@��Z���3@�q���!?�.�����@lDU�W�ٿpS����@��Z���3@�q���!?�.�����@��E���ٿ��귀�@`^�G�3@fQ����!?�����@��E���ٿ��귀�@`^�G�3@fQ����!?�����@��E���ٿ��귀�@`^�G�3@fQ����!?�����@�w�?��ٿ"�n���@����3@߰ed�!?�ӟ�2�@Zû�u�ٿ|�9�W1�@4��3@���!?��"�|�@Zû�u�ٿ|�9�W1�@4��3@���!?��"�|�@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�8>��ٿ��#����@��(���3@״	!?��7���@�O����ٿ����@���N�3@+u���!?�5�W��@�O����ٿ����@���N�3@+u���!?�5�W��@�O����ٿ����@���N�3@+u���!?�5�W��@�O����ٿ����@���N�3@+u���!?�5�W��@�O����ٿ����@���N�3@+u���!?�5�W��@o<hU�ٿ���{�@wpk��3@gH|�]�!?��T$��@o<hU�ٿ���{�@wpk��3@gH|�]�!?��T$��@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@ԒP�}�ٿlǬ��a�@���o�3@���{Ր!??S����@�����ٿ�6J���@ϵ!
��3@��}ճ�!?F��Y(&�@�����ٿ�6J���@ϵ!
��3@��}ճ�!?F��Y(&�@�����ٿ�6J���@ϵ!
��3@��}ճ�!?F��Y(&�@�����ٿ�6J���@ϵ!
��3@��}ճ�!?F��Y(&�@�����ٿ�6J���@ϵ!
��3@��}ճ�!?F��Y(&�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@O[`�ÞٿÈ��Ö�@$�Q;�3@<ȿY��!?�Y\�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@�O�X�ٿZH߄%�@�P��
�3@a���!?��J��H�@:b�ݣٿ�g��@�te�G�3@#�%���!?�8\a��@:b�ݣٿ�g��@�te�G�3@#�%���!?�8\a��@�Qe�R�ٿ�¬�:�@��M�S�3@JL���!?�nJ���@��3Q��ٿ��ԋh�@o�����3@f����!?�w��wJ�@��3Q��ٿ��ԋh�@o�����3@f����!?�w��wJ�@��3Q��ٿ��ԋh�@o�����3@f����!?�w��wJ�@��3Q��ٿ��ԋh�@o�����3@f����!?�w��wJ�@&m0�ٿ����0�@4[*���3@s_
��!?��ˑz�@&m0�ٿ����0�@4[*���3@s_
��!?��ˑz�@&m0�ٿ����0�@4[*���3@s_
��!?��ˑz�@��՛�ٿ���|9��@��!���3@N����!?3��E��@�M-Ȧٿ����@�g���3@�km��!?��7�0O�@�M-Ȧٿ����@�g���3@�km��!?��7�0O�@�M-Ȧٿ����@�g���3@�km��!?��7�0O�@�<��F�ٿ�'�V���@��b%��3@7<41ǐ!?Ί����@�<��F�ٿ�'�V���@��b%��3@7<41ǐ!?Ί����@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��W�(�ٿB��k��@9Ix���3@g!��ݐ!?36��(�@��b�ٿNIf\���@�����3@s��(Ӑ!?p�h���@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@���L�ٿ��|.}$�@����1�3@ߵ+��!?п����@�? 2��ٿ�߇����@�_՗��3@|�܇ؐ!?R��>��@�? 2��ٿ�߇����@�_՗��3@|�܇ؐ!?R��>��@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@ŭk�g�ٿ�=�I�@�����3@W���Ő!?�Y{d���@o�(u�ٿ6�W�$��@qN��3@6�/$z�!? 0p�+�@o�(u�ٿ6�W�$��@qN��3@6�/$z�!? 0p�+�@o�(u�ٿ6�W�$��@qN��3@6�/$z�!? 0p�+�@�Gm�ٿ0��}�@�P��X�3@��Ī�!?����{J�@�Gm�ٿ0��}�@�P��X�3@��Ī�!?����{J�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@XԿ���ٿ]�{Z��@YH/���3@/h�e��!?����,b�@�	HM�ٿ�N�P�@�p_���3@��,}�!?V3 .!��@�	HM�ٿ�N�P�@�p_���3@��,}�!?V3 .!��@bj��ӡٿ�-%@ڄ�@/e�$�3@��,n��!?�?����@bj��ӡٿ�-%@ڄ�@/e�$�3@��,n��!?�?����@��uiաٿ@���0�@�Q�ʷ�3@�_�Mې!?k�i�a�@��uiաٿ@���0�@�Q�ʷ�3@�_�Mې!?k�i�a�@��uiաٿ@���0�@�Q�ʷ�3@�_�Mې!?k�i�a�@B�e���ٿр���@��9ݕ�3@��uǴ�!?v.��`��@b\�+�ٿh���@Τ��3@�3�~ؐ!?�9�88&�@��]���ٿ�V��#�@�>Q�9�3@2�%��!?)j��C�@��]���ٿ�V��#�@�>Q�9�3@2�%��!?)j��C�@��]���ٿ�V��#�@�>Q�9�3@2�%��!?)j��C�@�Y���ٿ���}�P�@D�@�3@;AKwĐ!?W=U��@�Y���ٿ���}�P�@D�@�3@;AKwĐ!?W=U��@�Y���ٿ���}�P�@D�@�3@;AKwĐ!?W=U��@�Y���ٿ���}�P�@D�@�3@;AKwĐ!?W=U��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@Ub���ٿ�E�I��@��K�3@D���Đ!?��<�w��@^©F��ٿc���@�J�x�3@�K�
�!?��?���@@`h�A�ٿc"�T1�@"�$S��3@�T�!?b� k��@@`h�A�ٿc"�T1�@"�$S��3@�T�!?b� k��@@`h�A�ٿc"�T1�@"�$S��3@�T�!?b� k��@@`h�A�ٿc"�T1�@"�$S��3@�T�!?b� k��@?F�>��ٿnlHSY��@�EPv��3@/���!?�D�8vu�@?F�>��ٿnlHSY��@�EPv��3@/���!?�D�8vu�@�gAg=�ٿtۘ����@*��G��3@;[Ɛ!?_͟��8�@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@� �I�ٿ6�5R�@dJ���3@"��ِ!?������@s[z�|�ٿ������@��,zL�3@C���!?�Lܲ�	�@s[z�|�ٿ������@��,zL�3@C���!?�Lܲ�	�@s[z�|�ٿ������@��,zL�3@C���!?�Lܲ�	�@Wr�)8�ٿ� ��\�@r<�u�3@¯���!?�P���H�@'�����ٿU"�T/6�@Rĉ�D�3@�+��!?���2��@'�����ٿU"�T/6�@Rĉ�D�3@�+��!?���2��@'�����ٿU"�T/6�@Rĉ�D�3@�+��!?���2��@'�����ٿU"�T/6�@Rĉ�D�3@�+��!?���2��@A���F�ٿ#���@�@
Fx��3@�J����!?W��+��@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@깩�٢ٿw����@-%ۖ�3@�B�|�!?�����@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@�#.OH�ٿڄ1�$]�@f�P��3@��[m�!?(s��;��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@��O���ٿ�Ǚr��@�SVE/�3@��3�!?���A��@{�I��ٿ�����@2��i�3@�_�ː!?�$p��@{�I��ٿ�����@2��i�3@�_�ː!?�$p��@�Y�)�ٿ~g`�W�@7�a��3@���U�!?u.��%�@�Y�)�ٿ~g`�W�@7�a��3@���U�!?u.��%�@2B\[Q�ٿY]�M��@[�p��3@���pZ�!?��d��!�@@��n3�ٿ��U��@Rww�k�3@�R�3F�!?A,PW��@@��n3�ٿ��U��@Rww�k�3@�R�3F�!?A,PW��@@��n3�ٿ��U��@Rww�k�3@�R�3F�!?A,PW��@@��n3�ٿ��U��@Rww�k�3@�R�3F�!?A,PW��@@��n3�ٿ��U��@Rww�k�3@�R�3F�!?A,PW��@`�z�ٿ������@��-���3@z �+�!?�Sm|���@`�z�ٿ������@��-���3@z �+�!?�Sm|���@`�z�ٿ������@��-���3@z �+�!?�Sm|���@`�z�ٿ������@��-���3@z �+�!?�Sm|���@`�z�ٿ������@��-���3@z �+�!?�Sm|���@`�z�ٿ������@��-���3@z �+�!?�Sm|���@��0їٿ���ݿY�@3@��3@n����!?"��ן}�@��0їٿ���ݿY�@3@��3@n����!?"��ן}�@��:��ٿ�K&ë�@
0J�K�3@&ɠ�Q�!?���B� �@L󺜂�ٿ�k�@Rϳ��3@p3�_)�!?HsqJ�@��%���ٿחz�V��@.8���3@�8zkɐ!?��7�&C�@��%���ٿחz�V��@.8���3@�8zkɐ!?��7�&C�@��%���ٿחz�V��@.8���3@�8zkɐ!?��7�&C�@��%���ٿחz�V��@.8���3@�8zkɐ!?��7�&C�@��%���ٿחz�V��@.8���3@�8zkɐ!?��7�&C�@z@=�ٿ�̸��@̥"p9�3@��n'��!?H���N��@z@=�ٿ�̸��@̥"p9�3@��n'��!?H���N��@z@=�ٿ�̸��@̥"p9�3@��n'��!?H���N��@z@=�ٿ�̸��@̥"p9�3@��n'��!?H���N��@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@��<9�ٿ���'��@pG�z�3@A�`���!?/��W���@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@k�L���ٿ]`�Ÿq�@�Bv*�3@ْ8.�!?�j�yA�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@���S�ٿ�����@��d���3@�XԦ�!?��(&�;�@�+���ٿ���+�@3r`�(�3@ơӞ�!?��@N��@��+3�ٿ&���'��@0=E�f�3@)*��!?>H>b`��@��+3�ٿ&���'��@0=E�f�3@)*��!?>H>b`��@��+3�ٿ&���'��@0=E�f�3@)*��!?>H>b`��@��+3�ٿ&���'��@0=E�f�3@)*��!?>H>b`��@����ٿ2�UbA��@w!���3@�_�g��!?6���>��@����ٿ2�UbA��@w!���3@�_�g��!?6���>��@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@�P�U��ٿagbk���@v,���3@�I�_��!?33�8���@��~Z�ٿ4G��T�@>��p��3@�ѥ���!?���R���@��~Z�ٿ4G��T�@>��p��3@�ѥ���!?���R���@��~Z�ٿ4G��T�@>��p��3@�ѥ���!?���R���@��~Z�ٿ4G��T�@>��p��3@�ѥ���!?���R���@��~Z�ٿ4G��T�@>��p��3@�ѥ���!?���R���@2$5��ٿ��z���@~��b�3@7L�|�!?���&�@���}�ٿ5О�)2�@�a�M@�3@Y�EI��!?�)�o��@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��� �ٿ�pU��@8���R�3@�k�)�!?fv�q8�@��69�ٿ�+�#S�@�B�%�3@ �ǡ�!?��'�iX�@��69�ٿ�+�#S�@�B�%�3@ �ǡ�!?��'�iX�@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@����ٿ"4���:�@��E�p�3@��x��!?��7����@��)꘡ٿӎ��r��@�*���3@6��Aɐ!?�V�$P��@��)꘡ٿӎ��r��@�*���3@6��Aɐ!?�V�$P��@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�F�l�ٿ�^�,��@a&��3@����!?>�u�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@�m/�I�ٿs?���@[E1�1�3@eCȫe�!?�5��I�@P"f���ٿ��|��@�5~o�3@t�$�!?������@P"f���ٿ��|��@�5~o�3@t�$�!?������@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@�c1扞ٿ��d���@�?�)<�3@^
ᛐ!? ����e�@��M�E�ٿ�h4�s�@����I�3@'8z���!?�V(vw�@	>��ٿD�-���@���N��3@��-��!?^�h�jI�@	>��ٿD�-���@���N��3@��-��!?^�h�jI�@	>��ٿD�-���@���N��3@��-��!?^�h�jI�@	>��ٿD�-���@���N��3@��-��!?^�h�jI�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@,
��ʟٿ>�ʊ�@�V���3@��s��!?�(�/�@CǙǶ�ٿA7�K�!�@d�6��3@m�E��!?����@CǙǶ�ٿA7�K�!�@d�6��3@m�E��!?����@CǙǶ�ٿA7�K�!�@d�6��3@m�E��!?����@�b���ٿ11�u��@�M����3@�@y �!?�6��C)�@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@���(7�ٿ��Ҫ3B�@���;��3@Q%���!?G�����@����ǜٿ��׵���@��Ş�3@�7�y�!?Ciz0��@����ǜٿ��׵���@��Ş�3@�7�y�!?Ciz0��@����ǜٿ��׵���@��Ş�3@�7�y�!?Ciz0��@+/�ٿ"7����@�R�~u�3@�k����!?+\�����@+/�ٿ"7����@�R�~u�3@�k����!?+\�����@�����ٿv[�7�9�@�y��c�3@��p8��!?��3��@�����ٿv[�7�9�@�y��c�3@��p8��!?��3��@�����ٿ�oD�l�@_z�F��3@� h��!?˕��@�����ٿ�oD�l�@_z�F��3@� h��!?˕��@�����ٿ�oD�l�@_z�F��3@� h��!?˕��@�����ٿ�oD�l�@_z�F��3@� h��!?˕��@4�%
�ٿ9(Zcdx�@+�DA*�3@�0����!?�W�;]��@4�%
�ٿ9(Zcdx�@+�DA*�3@�0����!?�W�;]��@4�%
�ٿ9(Zcdx�@+�DA*�3@�0����!?�W�;]��@4�%
�ٿ9(Zcdx�@+�DA*�3@�0����!?�W�;]��@4�%
�ٿ9(Zcdx�@+�DA*�3@�0����!?�W�;]��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@w�����ٿ-��{�v�@,�t�3@�e\�!?���;��@��l�L�ٿ&ߋ�:�@\�0��3@�={n�!?*S��#�@��K�ٿ�b��@�<I�3@�Z�m��!?�\�5�@��K�ٿ�b��@�<I�3@�Z�m��!?�\�5�@�t>���ٿ��.�J�@`�xU�3@/����!?*�OSo��@�t>���ٿ��.�J�@`�xU�3@/����!?*�OSo��@ּ?�+�ٿ���.���@�-96�3@�khŞ�!?�Uŝ.��@ּ?�+�ٿ���.���@�-96�3@�khŞ�!?�Uŝ.��@ּ?�+�ٿ���.���@�-96�3@�khŞ�!?�Uŝ.��@ּ?�+�ٿ���.���@�-96�3@�khŞ�!?�Uŝ.��@ּ?�+�ٿ���.���@�-96�3@�khŞ�!?�Uŝ.��@Z�+M�ٿ�PѢ�@�&`�Z�3@/P�
��!?V�QN&o�@�Z=Z�ٿ���OFL�@v�r�}�3@�/��!?�[�ї�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@[x�-��ٿ8���Q�@2�e�r�3@_����!?��:��C�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@�֕�[�ٿA�����@��C�3@�hJײ�!?Le�):�@���x�ٿ��q�M��@!~C��3@ifj���!?�9ο���@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@�q��ٿᨾ�V��@ �zc��3@6!�a��!?�abZ�T�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@4���ˣٿo��9	�@�LW��3@�����!?��0�X�@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@�T�ٿܫgH�D�@�����3@[��!?֔��Q��@ �R8�ٿ:��q�@^���3@�7��!?!ȋ�'��@Eo��ٿh�W���@��ø��3@��� ��!?��'f��@Eo��ٿh�W���@��ø��3@��� ��!?��'f��@�����ٿ���N#��@Ħp3�3@(��!?l$��V��@�����ٿ���N#��@Ħp3�3@(��!?l$��V��@�����ٿ���N#��@Ħp3�3@(��!?l$��V��@9,0�ٿ��;�B�@T�Q��3@�n����!?������@Dx��ۡٿp�MN���@/����3@��Þ�!?5�V����@Dx��ۡٿp�MN���@/����3@��Þ�!?5�V����@Dx��ۡٿp�MN���@/����3@��Þ�!?5�V����@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@������ٿ��
���@��L=�3@6�����!? %Q-�H�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@q�i
1�ٿ�����,�@Z�\qi�3@��-�!? �}�"A�@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@N�h
��ٿ�ĭ�!@�@��E�3@�L��א!?#����@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@9h���ٿQ��=N��@/�
W�3@$K\j��!?�o���@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@�?�*�ٿ0�E�\L�@��3@]�؏�!?Y�����@m�-Нٿ���đ/�@�(K�X�3@;/@f��!?&U����@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@��Z�ٿ�a��X�@E�:t�3@�?�W��!?����	a�@�Z��ٿ!�1�
Q�@;Wo��3@K����!?�M�Y$��@�SQ�ٿ��'��@	����3@�_���!?�Rޟ�@��B���ٿ���+,Z�@,�M�3@ms�
��!?���c	�@f5=Ĩ�ٿ�U��U�@o͕��3@��a�!?:w�H�@f5=Ĩ�ٿ�U��U�@o͕��3@��a�!?:w�H�@f5=Ĩ�ٿ�U��U�@o͕��3@��a�!?:w�H�@ǵ���ٿD ����@F�H�Z�3@�ᡏ��!?&�����@ǵ���ٿD ����@F�H�Z�3@�ᡏ��!?&�����@�&
̝ٿ4�d�J=�@�Y�5j�3@I�G��!?�Y��s��@�&
̝ٿ4�d�J=�@�Y�5j�3@I�G��!?�Y��s��@���l�ٿc�����@W�+�3@���[�!?�WN�˞�@3��h�ٿ߲q�SL�@y^��"�3@T���g�!?�%����@��Bw�ٿ3�Z��@R~�,s�3@�j�*�!?�<$R�@��Bw�ٿ3�Z��@R~�,s�3@�j�*�!?�<$R�@��Bw�ٿ3�Z��@R~�,s�3@�j�*�!?�<$R�@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@�*?L��ٿ���y�@x3K��3@]�amݐ!?o�5��@%��.�ٿM�7����@^�߽�3@�Z䁩�!?�7����@%��.�ٿM�7����@^�߽�3@�Z䁩�!?�7����@%��.�ٿM�7����@^�߽�3@�Z䁩�!?�7����@%��.�ٿM�7����@^�߽�3@�Z䁩�!?�7����@%��.�ٿM�7����@^�߽�3@�Z䁩�!?�7����@��[*F�ٿ�w�N��@���V�3@�qtd��!?Se	�b�@��[*F�ٿ�w�N��@���V�3@�qtd��!?Se	�b�@��[*F�ٿ�w�N��@���V�3@�qtd��!?Se	�b�@����ٿ�[d| :�@6-xٚ�3@�ux��!?�t�0�R�@����ٿ�[d| :�@6-xٚ�3@�ux��!?�t�0�R�@f�iUz�ٿ�D=����@;ֵv�3@��NO��!?�Dإ5��@f�iUz�ٿ�D=����@;ֵv�3@��NO��!?�Dإ5��@f�iUz�ٿ�D=����@;ֵv�3@��NO��!?�Dإ5��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@u�����ٿ�$mmy��@������3@`�����!?��_��@��Z�G�ٿH�K�cT�@�v���3@��LQ��!?�V����@��Z�G�ٿH�K�cT�@�v���3@��LQ��!?�V����@����ٿ�~��*K�@��1E�3@���"Q�!?M˂�0�@�W�}��ٿd�n�@}_G��3@��s6d�!?sT�8��@�W�}��ٿd�n�@}_G��3@��s6d�!?sT�8��@�W�}��ٿd�n�@}_G��3@��s6d�!?sT�8��@�W�}��ٿd�n�@}_G��3@��s6d�!?sT�8��@�W�}��ٿd�n�@}_G��3@��s6d�!?sT�8��@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@9k����ٿ0s�F��@��D��3@�vb�А!?4� �6�@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@���V�ٿ7�v�@ �H���3@ Zy�Ő!?H�-���@i�D���ٿ�*���@��܊�3@��rÿ�!?��Y?n��@i�D���ٿ�*���@��܊�3@��rÿ�!?��Y?n��@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@	�����ٿ�|{?�@� ��b�3@���!?� �ly�@�;�{��ٿ)pP�1�@l� ]v�3@�ER�!?$�
m���@��ٿ{To���@��u-9�3@�t�`��!?���͸��@��ٿ{To���@��u-9�3@�t�`��!?���͸��@��ٿ{To���@��u-9�3@�t�`��!?���͸��@��ٿ{To���@��u-9�3@�t�`��!?���͸��@��ٿ{To���@��u-9�3@�t�`��!?���͸��@��ٿ{To���@��u-9�3@�t�`��!?���͸��@I_�(�ٿ�#�e]�@e�U
l�3@�C�}��!?��6A6�@��I��ٿ,���7b�@2�Aw�3@_h,E��!?<o�����@��I��ٿ,���7b�@2�Aw�3@_h,E��!?<o�����@��I��ٿ,���7b�@2�Aw�3@_h,E��!?<o�����@��I��ٿ,���7b�@2�Aw�3@_h,E��!?<o�����@��I��ٿ,���7b�@2�Aw�3@_h,E��!?<o�����@�%�Ө�ٿ�T�e���@�t2���3@�$���!?,#ŗϑ�@�%�Ө�ٿ�T�e���@�t2���3@�$���!?,#ŗϑ�@�%�Ө�ٿ�T�e���@�t2���3@�$���!?,#ŗϑ�@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@]��	\�ٿ��=rO�@��x���3@��}�А!?��w����@'��s�ٿ��3��@e�c_��3@��
~�!?k�[��@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@����}�ٿ�&�t;��@a!��3@%n���!?`�P�Ⱦ�@��߱b�ٿ_��Y���@�2U?O�3@t`����!?g�����@��߱b�ٿ_��Y���@�2U?O�3@t`����!?g�����@��߱b�ٿ_��Y���@�2U?O�3@t`����!?g�����@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@lV篨ٿV�e$��@F22yH�3@oaw��!?\:Ix�@���f�ٿ��%}W��@�?�8/�3@X�;1��!?F�
[w��@���f�ٿ��%}W��@�?�8/�3@X�;1��!?F�
[w��@d�8ܣٿ��R���@*�/rK�3@u.T�!?��Ƨ3�@d�8ܣٿ��R���@*�/rK�3@u.T�!?��Ƨ3�@d�8ܣٿ��R���@*�/rK�3@u.T�!?��Ƨ3�@���,��ٿ�\(���@[r�r��3@�*�\��!?�$
4C�@���,��ٿ�\(���@[r�r��3@�*�\��!?�$
4C�@���,��ٿ�\(���@[r�r��3@�*�\��!?�$
4C�@���,��ٿ�\(���@[r�r��3@�*�\��!?�$
4C�@?�2}�ٿ�j��@�C����3@�@�E�!?P����@?�2}�ٿ�j��@�C����3@�@�E�!?P����@?�2}�ٿ�j��@�C����3@�@�E�!?P����@?�2}�ٿ�j��@�C����3@�@�E�!?P����@lyBS.�ٿ#G�5��@tz�|-�3@ <W.�!?h� k���@lyBS.�ٿ#G�5��@tz�|-�3@ <W.�!?h� k���@lyBS.�ٿ#G�5��@tz�|-�3@ <W.�!?h� k���@lyBS.�ٿ#G�5��@tz�|-�3@ <W.�!?h� k���@e�:F��ٿ˄�B=C�@*��3@;�C���!?v$��W�@e�:F��ٿ˄�B=C�@*��3@;�C���!?v$��W�@)3I�z�ٿ�s��v�@�T�O�3@�geP��!?RU)�P�@)3I�z�ٿ�s��v�@�T�O�3@�geP��!?RU)�P�@)3I�z�ٿ�s��v�@�T�O�3@�geP��!?RU)�P�@)3I�z�ٿ�s��v�@�T�O�3@�geP��!?RU)�P�@)3I�z�ٿ�s��v�@�T�O�3@�geP��!?RU)�P�@��Z��ٿF��B�@S�Y4��3@͕��Ő!?�I+ &�@�1�{�ٿ"]�D��@\ 5���3@�X=֐!?p�2��@�1�{�ٿ"]�D��@\ 5���3@�X=֐!?p�2��@�1�{�ٿ"]�D��@\ 5���3@�X=֐!?p�2��@�1�{�ٿ"]�D��@\ 5���3@�X=֐!?p�2��@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@�\߀��ٿ�3z��@�А�3@�7S��!?�T���@,"���ٿ�j�9���@oh�f��3@�f��ʐ!?�����I�@,"���ٿ�j�9���@oh�f��3@�f��ʐ!?�����I�@NϣХٿݵp�_�@��z�+�3@ۼ�~�!?z ��@NϣХٿݵp�_�@��z�+�3@ۼ�~�!?z ��@4�A3�ٿ@�v����@�kW���3@�ڽ��!?�d0���@4�A3�ٿ@�v����@�kW���3@�ڽ��!?�d0���@4�A3�ٿ@�v����@�kW���3@�ڽ��!?�d0���@VK�1��ٿ�@/y�
�@�i��e�3@f��gÐ!?����@VK�1��ٿ�@/y�
�@�i��e�3@f��gÐ!?����@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@�fO��ٿ]���X��@�[�c�3@̈�C��!?��C��@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��j?�ٿ��S�/�@����3@��i���!?�u��5u�@��|��ٿ�DzRX��@�+ӯr�3@���qѐ!?9���W��@ ����ٿw�`�\w�@�}�a�3@��2Ő!?,�J�@m����ٿ�,J�
�@�X����3@�lŸ�!?��G���@Ҟ���ٿ�\E���@�f�g�3@���5�!?""nT��@Ҟ���ٿ�\E���@�f�g�3@���5�!?""nT��@B�sV�ٿ㼀J��@)J��Z�3@��'��!?�RfJ3�@�
���ٿfrW\���@�����3@},����!?]���4�@i�Q^ݜٿ�d�����@���6U�3@�;MkƐ!?�P���@��q{
�ٿv�#��D�@�ș#��3@��[�Ð!?��/z�@��q{
�ٿv�#��D�@�ș#��3@��[�Ð!?��/z�@��q{
�ٿv�#��D�@�ș#��3@��[�Ð!?��/z�@��q{
�ٿv�#��D�@�ș#��3@��[�Ð!?��/z�@%���ٿǛ����@;��]�3@{}3��!?d/�3�@%���ٿǛ����@;��]�3@{}3��!?d/�3�@%���ٿǛ����@;��]�3@{}3��!?d/�3�@%���ٿǛ����@;��]�3@{}3��!?d/�3�@5�D�ٿX�?#*��@\�����3@�Z��!?��a�A��@5�D�ٿX�?#*��@\�����3@�Z��!?��a�A��@5�D�ٿX�?#*��@\�����3@�Z��!?��a�A��@5�D�ٿX�?#*��@\�����3@�Z��!?��a�A��@��u3��ٿ�j ����@���I:�3@R�] ��!?j�˼�@��u3��ٿ�j ����@���I:�3@R�] ��!?j�˼�@��u3��ٿ�j ����@���I:�3@R�] ��!?j�˼�@��u3��ٿ�j ����@���I:�3@R�] ��!?j�˼�@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@/iUp�ٿ���%f�@�aa��3@�ǋ�Ɛ!?�����@� ��ڡٿ����9�@��#^�3@��s�!?9�i����@'��u$�ٿU�y��k�@T�>ɉ�3@��?�!?�dm3�@'��u$�ٿU�y��k�@T�>ɉ�3@��?�!?�dm3�@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@�F<u�ٿƥ�9c�@�j�\��3@���
�!?��M����@y�(�.�ٿ��6*x<�@��#�3@�C���!?}��1!�@y�(�.�ٿ��6*x<�@��#�3@�C���!?}��1!�@�`)5��ٿ�E���@���`��3@[���!?�\�>�:�@Z��ٿ���S�/�@:��e�3@rU�Ő!?�y����@�e��ٿ1�%����@@�'6�3@�b����!?�����a�@�e��ٿ1�%����@@�'6�3@�b����!?�����a�@�e��ٿ1�%����@@�'6�3@�b����!?�����a�@U��j�ٿ�����@_�R��3@LJ���!?�O�\�@U��j�ٿ�����@_�R��3@LJ���!?�O�\�@U��j�ٿ�����@_�R��3@LJ���!?�O�\�@]�3H�ٿ{�p����@;8���3@Z}��~�!?���^��@]�3H�ٿ{�p����@;8���3@Z}��~�!?���^��@#����ٿ�l���@�xmF�3@��5���!?X1���5�@#����ٿ�l���@�xmF�3@��5���!?X1���5�@#����ٿ�l���@�xmF�3@��5���!?X1���5�@��⇡ٿ����v��@���O��3@���7�!?8��d��@��⇡ٿ����v��@���O��3@���7�!?8��d��@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@'w��Ǥٿ�w�͓��@��'��3@%�����!?4�����@ƶ�8\�ٿG�K@_�@�Ճm��3@։/"�!?^9��7��@ƶ�8\�ٿG�K@_�@�Ճm��3@։/"�!?^9��7��@ƶ�8\�ٿG�K@_�@�Ճm��3@։/"�!?^9��7��@��mԥٿK��>�D�@�����3@P� �(�!?���_�@��mԥٿK��>�D�@�����3@P� �(�!?���_�@{��ƥٿs�E��@��R���3@�����!?37'�~�@{��ƥٿs�E��@��R���3@�����!?37'�~�@{��ƥٿs�E��@��R���3@�����!?37'�~�@{��ƥٿs�E��@��R���3@�����!?37'�~�@�n����ٿY lmPF�@�c��3@�$vY�!?l�*�nQ�@�n����ٿY lmPF�@�c��3@�$vY�!?l�*�nQ�@�n����ٿY lmPF�@�c��3@�$vY�!?l�*�nQ�@�n����ٿY lmPF�@�c��3@�$vY�!?l�*�nQ�@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@�\ȭ�ٿ8i���@�Yo)��3@������!?�Ŋ����@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@]�� ��ٿ���V�@]�Wc��3@�_s���!?�c�nP��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@!��_�ٿQF�0�\�@�IX�U�3@�|���!?��a��@1/"#�ٿ��A;�@��|~�3@���"g�!?l�GM��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@Y��ٿ�dc0`6�@J{Ϫ�3@Δ���!?e�w_��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@���̟ٿ�܋i�@Kc���3@	���!?ph�^K��@՜��ٿ�`"���@}�w)}�3@�粈�!?PG؄��@՜��ٿ�`"���@}�w)}�3@�粈�!?PG؄��@՜��ٿ�`"���@}�w)}�3@�粈�!?PG؄��@w2����ٿ�� ���@,�R���3@�jА!?��3��M�@w2����ٿ�� ���@,�R���3@�jА!?��3��M�@w2����ٿ�� ���@,�R���3@�jА!?��3��M�@w2����ٿ�� ���@,�R���3@�jА!?��3��M�@w2����ٿ�� ���@,�R���3@�jА!?��3��M�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X�{�_�ٿz��T-4�@�I��3@a��&��!?���L�@X����ٿ��&n�@OP@��3@P&9T�!?�:��h�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@/�\��ٿ��o����@�8�Y��3@:}f��!?sΆ8�@+	D$K�ٿ�?+�P�@�
߃��3@'ѰV��!?	x�҄��@+	D$K�ٿ�?+�P�@�
߃��3@'ѰV��!?	x�҄��@+	D$K�ٿ�?+�P�@�
߃��3@'ѰV��!?	x�҄��@+	D$K�ٿ�?+�P�@�
߃��3@'ѰV��!?	x�҄��@&���h�ٿY�q&��@^�����3@ʟ� �!?�2���@&���h�ٿY�q&��@^�����3@ʟ� �!?�2���@&���h�ٿY�q&��@^�����3@ʟ� �!?�2���@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@ߚ��ٿYT����@|� Q��3@�nf�͐!?<-uƺ �@oalÝٿ�� R��@�3�0��3@���.א!?CL��@��ȡ��ٿ~�0�S�@VN���3@L�����!?�0l��@��ȡ��ٿ~�0�S�@VN���3@L�����!?�0l��@�u{��ٿ�1Qߐ9�@��V:�3@��,*�!?R�����@�u{��ٿ�1Qߐ9�@��V:�3@��,*�!?R�����@�u{��ٿ�1Qߐ9�@��V:�3@��,*�!?R�����@�u{��ٿ�1Qߐ9�@��V:�3@��,*�!?R�����@�u{��ٿ�1Qߐ9�@��V:�3@��,*�!?R�����@��N%��ٿ������@���] �3@���J�!?Y��;�@W��Ûٿ��"�R�@#�r�3@��j#�!?b�r���@W��Ûٿ��"�R�@#�r�3@��j#�!?b�r���@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@K)��ٿ�}r5�@o>xJ��3@�ѐ!?m�1�q�@��f3�ٿ N1��@���#��3@����ؐ!?��\���@��f3�ٿ N1��@���#��3@����ؐ!?��\���@��f3�ٿ N1��@���#��3@����ؐ!?��\���@��f3�ٿ N1��@���#��3@����ؐ!?��\���@��f3�ٿ N1��@���#��3@����ؐ!?��\���@FTaC��ٿ�3Z����@�H�j�3@~��!?MvQ#��@FTaC��ٿ�3Z����@�H�j�3@~��!?MvQ#��@FTaC��ٿ�3Z����@�H�j�3@~��!?MvQ#��@s�6r�ٿ�ϸr�@\��͋�3@�.��!?�8ę,��@s�6r�ٿ�ϸr�@\��͋�3@�.��!?�8ę,��@s�6r�ٿ�ϸr�@\��͋�3@�.��!?�8ę,��@���r��ٿR�'���@�4�"�3@@�	�ǐ!?���I�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@���߄�ٿ:�5�@'岰�3@�,����!?�in�67�@h�H��ٿFJy��@*����3@=�hې!?O)C��$�@h�H��ٿFJy��@*����3@=�hې!?O)C��$�@h�H��ٿFJy��@*����3@=�hې!?O)C��$�@�(}��ٿ#<hP��@(��B��3@G���ߐ!?c#Ӊ��@�(}��ٿ#<hP��@(��B��3@G���ߐ!?c#Ӊ��@����ٿ���W���@> :5��3@��+Š�!?#��	���@����ٿ���W���@> :5��3@��+Š�!?#��	���@����ٿ���W���@> :5��3@��+Š�!?#��	���@�l̃��ٿz��|2q�@�n0(�3@�Q1{��!?/��V��@�l̃��ٿz��|2q�@�n0(�3@�Q1{��!?/��V��@�l̃��ٿz��|2q�@�n0(�3@�Q1{��!?/��V��@�l̃��ٿz��|2q�@�n0(�3@�Q1{��!?/��V��@��?W�ٿh��'�@a���2�3@�-h��!?*z��	�@\oO�@�ٿ��Nuf��@�0؎��3@j�+��!?D�"��H�@\oO�@�ٿ��Nuf��@�0؎��3@j�+��!?D�"��H�@^Kq<4�ٿ���ê9�@<�7��3@�®Ő!?��Lq�M�@^Kq<4�ٿ���ê9�@<�7��3@�®Ő!?��Lq�M�@^Kq<4�ٿ���ê9�@<�7��3@�®Ő!?��Lq�M�@^�e��ٿ�t/J���@��1���3@\���!?�z����@x��ٿ�r`I���@*Tؔ�3@�H�?�!?z�V~�s�@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@]#�|��ٿ�jx{ �@�~�w�3@&�]s%�!?ѭ�'���@�ju�ٿ�A��(�@G��@�3@�#��?�!?��GR�,�@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@c���ٿu7��W.�@	��F��3@Q1��!?�����@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@2�L���ٿ���C�@`_���3@���Ԑ!?	,Z�N�@�Q�	�ٿ�A�@,b!7�3@�8Ð!?>�i({{�@�Q�	�ٿ�A�@,b!7�3@�8Ð!?>�i({{�@�Q�	�ٿ�A�@,b!7�3@�8Ð!?>�i({{�@�Q�	�ٿ�A�@,b!7�3@�8Ð!?>�i({{�@i��.�ٿ������@�X$hW�3@1C��ϐ!?Pg��?�@i��.�ٿ������@�X$hW�3@1C��ϐ!?Pg��?�@i��.�ٿ������@�X$hW�3@1C��ϐ!?Pg��?�@i��.�ٿ������@�X$hW�3@1C��ϐ!?Pg��?�@i��.�ٿ������@�X$hW�3@1C��ϐ!?Pg��?�@��O>�ٿ�6ޕ1�@x!���3@�[�RƐ!?'��b�@�\�bǣٿT!
y���@��A�`�3@q�q� �!?����@�\�bǣٿT!
y���@��A�`�3@q�q� �!?����@�\�bǣٿT!
y���@��A�`�3@q�q� �!?����@a���@�ٿ�o����@�1#^�3@j��!?<�U���@a���@�ٿ�o����@�1#^�3@j��!?<�U���@a���@�ٿ�o����@�1#^�3@j��!?<�U���@a���@�ٿ�o����@�1#^�3@j��!?<�U���@[����ٿ��د�@����3@�+��!?j vA�"�@[����ٿ��د�@����3@�+��!?j vA�"�@[����ٿ��د�@����3@�+��!?j vA�"�@�U�t3�ٿ�Ga�\��@����3@)mV� �!?x��6��@�P���ٿ[V�jɺ�@��j[�3@pN@�!?<!��A�@�P���ٿ[V�jɺ�@��j[�3@pN@�!?<!��A�@�a�?�ٿ2<h����@v���3@�*{��!?��u�L"�@�a�?�ٿ2<h����@v���3@�*{��!?��u�L"�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@p�B�àٿ�a�����@^w{$�3@��u��!?�Ȓ]v%�@0�P�q�ٿ쿝(r��@K]�+�3@�� �x�!?;g߰)=�@0�P�q�ٿ쿝(r��@K]�+�3@�� �x�!?;g߰)=�@���b�ٿ�y�\ �@E�x��3@�SM3v�!?!"/����@���b�ٿ�y�\ �@E�x��3@�SM3v�!?!"/����@���b�ٿ�y�\ �@E�x��3@�SM3v�!?!"/����@���b�ٿ�y�\ �@E�x��3@�SM3v�!?!"/����@���b�ٿ�y�\ �@E�x��3@�SM3v�!?!"/����@~��#�ٿ��z)�@:��w]�3@>���!?�PLI1�@~��#�ٿ��z)�@:��w]�3@>���!?�PLI1�@~��#�ٿ��z)�@:��w]�3@>���!?�PLI1�@~��#�ٿ��z)�@:��w]�3@>���!?�PLI1�@��<s!�ٿqGb���@�=�U�3@&5!5�!?e�VP�'�@̞%���ٿЏ����@Rm<��3@�r��!?�l��Li�@̞%���ٿЏ����@Rm<��3@�r��!?�l��Li�@̞%���ٿЏ����@Rm<��3@�r��!?�l��Li�@����#�ٿG*1̶�@N�c�>�3@���vX�!?[jٸC �@����#�ٿG*1̶�@N�c�>�3@���vX�!?[jٸC �@����#�ٿG*1̶�@N�c�>�3@���vX�!?[jٸC �@����#�ٿG*1̶�@N�c�>�3@���vX�!?[jٸC �@����#�ٿG*1̶�@N�c�>�3@���vX�!?[jٸC �@�ۨ5�ٿ�t�";�@c.�=*�3@6ؕ�!?գ>߷��@�i�"�ٿ���Y�@`�	��3@���zb�!?9j�N�'�@�t�ŝ�ٿJ+S����@";`�3@h	
��!?��qϬ�@�t�ŝ�ٿJ+S����@";`�3@h	
��!?��qϬ�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@Bw��Ǣٿ�����@[z�3@��r��!?2�v�8�@����՛ٿ.�pj<��@�ԛ�h�3@�Lځ��!?�n�H�F�@����՛ٿ.�pj<��@�ԛ�h�3@�Lځ��!?�n�H�F�@����՛ٿ.�pj<��@�ԛ�h�3@�Lځ��!?�n�H�F�@����՛ٿ.�pj<��@�ԛ�h�3@�Lځ��!?�n�H�F�@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@Օ�@�ٿ����e��@Щ ��3@���ڐ!?��t&���@�w���ٿWi�a��@��|&�3@��$@ΐ!?�/��Y�@�w���ٿWi�a��@��|&�3@��$@ΐ!?�/��Y�@�w���ٿWi�a��@��|&�3@��$@ΐ!?�/��Y�@�5�$��ٿu��NA��@���x��3@�oP���!?�����@�5�$��ٿu��NA��@���x��3@�oP���!?�����@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@>��W�ٿK�Q��'�@�3 n�3@'�˔�!?��0A���@��|zY�ٿ�c��Th�@6ٞ�u�3@���x�!?Y�6@��@��|zY�ٿ�c��Th�@6ٞ�u�3@���x�!?Y�6@��@��|zY�ٿ�c��Th�@6ٞ�u�3@���x�!?Y�6@��@��|zY�ٿ�c��Th�@6ٞ�u�3@���x�!?Y�6@��@S�ٿ��(����@����3@xH����!?�;�oL��@S�ٿ��(����@����3@xH����!?�;�oL��@S�ٿ��(����@����3@xH����!?�;�oL��@��Y�Шٿ���OC�@�{����3@��c��!?<�|@�@��ƵP�ٿE��Dw#�@Wm�D�3@a�Hڐ!?�G�hq�@��ƵP�ٿE��Dw#�@Wm�D�3@a�Hڐ!?�G�hq�@��ƵP�ٿE��Dw#�@Wm�D�3@a�Hڐ!?�G�hq�@��ƵP�ٿE��Dw#�@Wm�D�3@a�Hڐ!?�G�hq�@��ƵP�ٿE��Dw#�@Wm�D�3@a�Hڐ!?�G�hq�@u�]L��ٿ;Ű��@S�	H��3@���8��!?6���Jq�@u�]L��ٿ;Ű��@S�	H��3@���8��!?6���Jq�@u�]L��ٿ;Ű��@S�	H��3@���8��!?6���Jq�@u�]L��ٿ;Ű��@S�	H��3@���8��!?6���Jq�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@��.�ԟٿp������@��c�x�3@lUM���!?l]à�@�`9K�ٿ���F�@_���@�3@J�p�!?:B*0���@�`9K�ٿ���F�@_���@�3@J�p�!?:B*0���@
����ٿ}�W��@j`يh�3@������!?v����@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@}��۠ٿx�w�>�@0R;z��3@r��ڐ!?	"�w��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�cߟ�ٿ�֒��@+Q$�3@�����!?Z��E��@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@�ഗ�ٿк�~�O�@����3@�f�Ð!?jh���V�@!	��6�ٿ�I�q\2�@�����3@x|ؐ!?�eY9��@!	��6�ٿ�I�q\2�@�����3@x|ؐ!?�eY9��@P� K�ٿ��0����@S�S���3@���wӐ!?A�'P��@P� K�ٿ��0����@S�S���3@���wӐ!?A�'P��@P� K�ٿ��0����@S�S���3@���wӐ!?A�'P��@P� K�ٿ��0����@S�S���3@���wӐ!?A�'P��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�{0V��ٿ�^9G#�@p���3@X�r��!?N��&��@�k���ٿ�J�EC2�@��z��3@���ֹ�!?��E���@�k���ٿ�J�EC2�@��z��3@���ֹ�!?��E���@�E���ٿ�9x��@ցÏ��3@]�
���!?"�:���@�E���ٿ�9x��@ցÏ��3@]�
���!?"�:���@�E���ٿ�9x��@ցÏ��3@]�
���!?"�:���@U��K��ٿ������@6\����3@���	ې!?�|��j��@�$t�؛ٿo�\��@Oϑ���3@��_��!?�蒲NY�@�$t�؛ٿo�\��@Oϑ���3@��_��!?�蒲NY�@�S���ٿ"�#����@���]�3@r�*7��!?���@�S���ٿ"�#����@���]�3@r�*7��!?���@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@�d�.��ٿ74�A��@v�o�3@Rj1���!?1��Ǹ�@^�	UZ�ٿXV>�F�@�;����3@�`Ր!?S�Ժ��@^�	UZ�ٿXV>�F�@�;����3@�`Ր!?S�Ժ��@��
*��ٿ5�E��@"���x�3@��~���!?!������@��
*��ٿ5�E��@"���x�3@��~���!?!������@��
*��ٿ5�E��@"���x�3@��~���!?!������@��
*��ٿ5�E��@"���x�3@��~���!?!������@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@��k	�ٿd������@M*F�3@'?z���!?叡�7�@F�0ݠٿ�S��17�@�IN�`�3@mjU��!?0C�.�@F�0ݠٿ�S��17�@�IN�`�3@mjU��!?0C�.�@F�0ݠٿ�S��17�@�IN�`�3@mjU��!?0C�.�@��g��ٿ	��A��@-F�A��3@��ѐ!?�OC3<��@��g��ٿ	��A��@-F�A��3@��ѐ!?�OC3<��@��g��ٿ	��A��@-F�A��3@��ѐ!?�OC3<��@��g��ٿ	��A��@-F�A��3@��ѐ!?�OC3<��@��g��ٿ	��A��@-F�A��3@��ѐ!?�OC3<��@�-�.��ٿ�����@��k=��3@@%nrѐ!?�:���@{��hD�ٿ]>�����@���5�3@T��V�!?�WYX*�@{��hD�ٿ]>�����@���5�3@T��V�!?�WYX*�@{��hD�ٿ]>�����@���5�3@T��V�!?�WYX*�@{��hD�ٿ]>�����@���5�3@T��V�!?�WYX*�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@E>%҈�ٿ䬵 ��@���j��3@ݳ�y�!?�q��<b�@�>�_��ٿ��c"ۧ�@x*����3@n�iꛐ!?Oq�Av�@�>�_��ٿ��c"ۧ�@x*����3@n�iꛐ!?Oq�Av�@�>�_��ٿ��c"ۧ�@x*����3@n�iꛐ!?Oq�Av�@�>�_��ٿ��c"ۧ�@x*����3@n�iꛐ!?Oq�Av�@.�HC��ٿ-k}��y�@!�~��3@����!?�N���@.�HC��ٿ-k}��y�@!�~��3@����!?�N���@�W�+��ٿ>E*���@���0z�3@�0�(`�!?O(@��@�W�+��ٿ>E*���@���0z�3@�0�(`�!?O(@��@�W�+��ٿ>E*���@���0z�3@�0�(`�!?O(@��@��o쩧ٿ�H����@A���3@R)A���!?��G�$��@��o쩧ٿ�H����@A���3@R)A���!?��G�$��@�4��	�ٿ�o�/�@5ڄ�;�3@|�+x��!?�<tL4�@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@x-XCX�ٿ�Z��l�@嚴���3@��2���!?e��w���@ƴ�?B�ٿ��fT_��@y-8���3@)+9%��!?�y�����@����ٿpOF���@� Ԯ��3@�<x{�!?L��Kg�@����ٿpOF���@� Ԯ��3@�<x{�!?L��Kg�@����ٿpOF���@� Ԯ��3@�<x{�!?L��Kg�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@Ҏfk"�ٿU- )5��@v����3@��
��!?;��b�F�@(�ʒ��ٿ�PH4���@��_`�3@XI_��!?�2n��@�"C�ٿ4����@Џ��J�3@�	)��!?ˊA|��@�"C�ٿ4����@Џ��J�3@�	)��!?ˊA|��@D^�8؟ٿ���#}I�@~n5���3@�w����!?'
��Z��@M�m�ؠٿ&�B�,��@5�(Z��3@Y{�K��!?��)����@M�m�ؠٿ&�B�,��@5�(Z��3@Y{�K��!?��)����@M�m�ؠٿ&�B�,��@5�(Z��3@Y{�K��!?��)����@M�m�ؠٿ&�B�,��@5�(Z��3@Y{�K��!?��)����@r��z�ٿ�G�@q���&�3@4��Ɛ!?�����@r��z�ٿ�G�@q���&�3@4��Ɛ!?�����@r��z�ٿ�G�@q���&�3@4��Ɛ!?�����@r��z�ٿ�G�@q���&�3@4��Ɛ!?�����@N�`�ٿ�׈K
�@���#��3@L ��А!?x@�_���@N�`�ٿ�׈K
�@���#��3@L ��А!?x@�_���@N�`�ٿ�׈K
�@���#��3@L ��А!?x@�_���@N�`�ٿ�׈K
�@���#��3@L ��А!?x@�_���@N�`�ٿ�׈K
�@���#��3@L ��А!?x@�_���@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@*!�P �ٿDtVFe��@�+#t��3@7S�:�!?j?[����@�����ٿ������@6=�`�3@DA��!?�uLν�@�����ٿ������@6=�`�3@DA��!?�uLν�@e��
=�ٿ,�	B5��@��n$��3@�IU��!?ʷ�����@e��
=�ٿ,�	B5��@��n$��3@�IU��!?ʷ�����@	��ٿ�h[+�@�R���3@eI���!?���Ɉ�@	��ٿ�h[+�@�R���3@eI���!?���Ɉ�@	��ٿ�h[+�@�R���3@eI���!?���Ɉ�@	��ٿ�h[+�@�R���3@eI���!?���Ɉ�@U���h�ٿD�U`���@D׶��3@��J��!?L'�
�C�@U���h�ٿD�U`���@D׶��3@��J��!?L'�
�C�@���ٿ.�Hf��@�$m��3@b����!?j�� H��@���ٿ.�Hf��@�$m��3@b����!?j�� H��@���ٿ.�Hf��@�$m��3@b����!?j�� H��@���ٿ.�Hf��@�$m��3@b����!?j�� H��@�/�q�ٿ&0��@�����3@����!?S��N��@�/�q�ٿ&0��@�����3@����!?S��N��@cI���ٿ�_��I�@=�N�3@������!?5퓑���@$Z�y�ٿ��0r�x�@�t(�3@��ы�!?#7ˑ���@$Z�y�ٿ��0r�x�@�t(�3@��ы�!?#7ˑ���@4�} ��ٿ��y�U��@�y���3@jA{�!?hF��!��@4�} ��ٿ��y�U��@�y���3@jA{�!?hF��!��@4�} ��ٿ��y�U��@�y���3@jA{�!?hF��!��@ XE���ٿ�`db�@t��)��3@r�ǐ!?�v��j�@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@ߖ�-��ٿ[�V�%��@��j/#�3@�Yk缐!?w�k"���@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@�3�8�ٿn�zؼ�@�/=�3@'��>��!?j��k�K�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@nj�t	�ٿ_�%����@ݵ�}��3@���wؐ!?��/�jO�@ ����ٿ�[���]�@Hu���3@{���Ӑ!?�H�/�u�@ ����ٿ�[���]�@Hu���3@{���Ӑ!?�H�/�u�@ ����ٿ�[���]�@Hu���3@{���Ӑ!?�H�/�u�@�O����ٿZt�*q�@�=��5�3@�V��ؐ!?d�\�Gy�@-N^dR�ٿι�෡�@O5��3@p��a�!?��y�r��@-N^dR�ٿι�෡�@O5��3@p��a�!?��y�r��@-N^dR�ٿι�෡�@O5��3@p��a�!?��y�r��@-N^dR�ٿι�෡�@O5��3@p��a�!?��y�r��@  �S�ٿ�1.-F1�@|)��^�3@[L?�p�!?
�����@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@
�DȨ�ٿ��I����@Z�yR�3@|ಢ��!?���F���@����U�ٿtJ�^0l�@�4���3@��0&_�!?�s�u�4�@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@!}��ٿ]3pxh�@lS�Iu�3@x�|Լ�!?�����@� ��ٿJI%���@U�����3@���e��!?r�ӓa�@� ��ٿJI%���@U�����3@���e��!?r�ӓa�@� ��ٿJI%���@U�����3@���e��!?r�ӓa�@� ��ٿJI%���@U�����3@���e��!?r�ӓa�@�Vs�ٿ�4wRs�@�x�۳�3@JNk��!?B�s'�@8^Zv~�ٿĢW�=�@���ˮ�3@���~��!? v&<#�@8^Zv~�ٿĢW�=�@���ˮ�3@���~��!? v&<#�@�V�Q�ٿ!^��!��@�@����3@9㖽�!?��^�m��@�V�Q�ٿ!^��!��@�@����3@9㖽�!?��^�m��@�V�Q�ٿ!^��!��@�@����3@9㖽�!?��^�m��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@�Pvp��ٿ�7��@wf�N�3@�®�А!?����k��@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@Iӣ��ٿ�ɛK���@|�=��3@��`��!?uR^���@�`�	��ٿ|���s��@1�:%��3@�b�D�!?Eߵ#���@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@���U��ٿ�5�F���@��8:��3@�ls�!?D�D[��@\!�3�ٿ�d�(K��@4x����3@y��	�!?�ᬢ��@\!�3�ٿ�d�(K��@4x����3@y��	�!?�ᬢ��@�~TߝٿŤR$^��@BjTus�3@�/8�ʐ!?��)%�8�@�~TߝٿŤR$^��@BjTus�3@�/8�ʐ!?��)%�8�@�~TߝٿŤR$^��@BjTus�3@�/8�ʐ!?��)%�8�@�a\ǚٿ� W%��@�s6O$�3@D��ڭ�!?�z�R�<�@�wu6��ٿ�Q~�~��@���s�3@�l�А!?L���>�@�wu6��ٿ�Q~�~��@���s�3@�l�А!?L���>�@�wu6��ٿ�Q~�~��@���s�3@�l�А!?L���>�@I��\̛ٿك�,D�@�?��6�3@�$�7��!?�I�d�L�@R���ޣٿ�%���@p����3@��x Ð!?��l�@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@b��$�ٿjbB���@j�����3@
-'"А!?,!IqW��@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@x2J~Ģٿ�6��x��@OZ�'?�3@VD���!?�E����@��॥ٿ��?&+C�@cz��q�3@��Ő!?��\���@��॥ٿ��?&+C�@cz��q�3@��Ő!?��\���@��॥ٿ��?&+C�@cz��q�3@��Ő!?��\���@�;�ϧٿEu���@�c��3@��Ά��!?�t�3�h�@�;�ϧٿEu���@�c��3@��Ά��!?�t�3�h�@ȭ8K٤ٿ4��(���@�h����3@�� �ϐ!?��4����@ȭ8K٤ٿ4��(���@�h����3@�� �ϐ!?��4����@ȭ8K٤ٿ4��(���@�h����3@�� �ϐ!?��4����@����|�ٿ|�����@J�[�/�3@�ݶ�!?8��yL�@����|�ٿ|�����@J�[�/�3@�ݶ�!?8��yL�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@sK��=�ٿ��_��@0�'��3@d����!?o�_p�1�@Z3A��ٿ���K�Q�@����3@������!?u����@Z3A��ٿ���K�Q�@����3@������!?u����@Z3A��ٿ���K�Q�@����3@������!?u����@Z3A��ٿ���K�Q�@����3@������!?u����@Z3A��ٿ���K�Q�@����3@������!?u����@Z3A��ٿ���K�Q�@����3@������!?u����@Xxq�ݣٿN�8��@���X-�3@��R�ߐ!?�"C�7.�@Xxq�ݣٿN�8��@���X-�3@��R�ߐ!?�"C�7.�@Xxq�ݣٿN�8��@���X-�3@��R�ߐ!?�"C�7.�@Xxq�ݣٿN�8��@���X-�3@��R�ߐ!?�"C�7.�@VPܸ��ٿ�~�@���@��$��3@�:[�ِ!?������@VPܸ��ٿ�~�@���@��$��3@�:[�ِ!?������@VPܸ��ٿ�~�@���@��$��3@�:[�ِ!?������@:�߉-�ٿ��J>��@�I�2��3@ut�!?���K��@:�߉-�ٿ��J>��@�I�2��3@ut�!?���K��@:�߉-�ٿ��J>��@�I�2��3@ut�!?���K��@��5��ٿzw�PP��@����]�3@�򼎬�!?�^1O�@��5��ٿzw�PP��@����]�3@�򼎬�!?�^1O�@��5��ٿzw�PP��@����]�3@�򼎬�!?�^1O�@��5��ٿzw�PP��@����]�3@�򼎬�!?�^1O�@��5��ٿzw�PP��@����]�3@�򼎬�!?�^1O�@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@CF�g�ٿ�+G��@e�:
��3@��Ր!?�4�Eo��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��t��ٿ�u���@�W�3@����ِ!?��5,��@��YZ�ٿ��$^���@�H����3@W���Ɛ!?=�����@�g��ßٿ�������@A2���3@ 50��!?%�ִ��@�g��ßٿ�������@A2���3@ 50��!?%�ִ��@�g��ßٿ�������@A2���3@ 50��!?%�ִ��@��!TS�ٿ��8��@�T�3@[z
���!?܏�0Hj�@�c�ٿ$N��͵�@���8L�3@�5�%�!?A������@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@#ކv��ٿec��$�@�˧5��3@���+��!?WO�f��@'���ٿXbt\S��@=R��f�3@��8�!?p���#�@'���ٿXbt\S��@=R��f�3@��8�!?p���#�@'���ٿXbt\S��@=R��f�3@��8�!?p���#�@'���ٿXbt\S��@=R��f�3@��8�!?p���#�@t�x���ٿ���!��@���^[�3@��!��!?m�1�$�@t�x���ٿ���!��@���^[�3@��!��!?m�1�$�@t�x���ٿ���!��@���^[�3@��!��!?m�1�$�@t�x���ٿ���!��@���^[�3@��!��!?m�1�$�@t�x���ٿ���!��@���^[�3@��!��!?m�1�$�@�QI�ٿE�d� �@;�3���3@o�Ă�!?up����@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@�!!%�ٿ��F�@�r���3@t.��!?+�v���@J|W�ٿ�S�ny�@,0�y�3@(���!?z�n0�$�@J|W�ٿ�S�ny�@,0�y�3@(���!?z�n0�$�@J|W�ٿ�S�ny�@,0�y�3@(���!?z�n0�$�@J|W�ٿ�S�ny�@,0�y�3@(���!?z�n0�$�@"��'�ٿ������@ޡ�r��3@xsߐ!?A�$?��@���|N�ٿ/t�8-E�@@wTiJ�3@M����!?�Κ�1�@���|N�ٿ/t�8-E�@@wTiJ�3@M����!?�Κ�1�@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@W�s��ٿ��Q���@+�%K�3@�w���!?�iB���@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@mC��ٿ��FT�T�@���x��3@isS$�!?S�����@�|���ٿ���^�$�@�Z�@��3@�e!Z�!?|D���=�@�|���ٿ���^�$�@�Z�@��3@�e!Z�!?|D���=�@�|���ٿ���^�$�@�Z�@��3@�e!Z�!?|D���=�@oAyJ%�ٿ��>���@�7@��3@%�m+�!?������@����љٿf�f�^�@�19�3@���*>�!?�ӻ�Rv�@4:\ߞٿa��Wؙ�@�xa3B�3@�����!? �*ҷ*�@4:\ߞٿa��Wؙ�@�xa3B�3@�����!? �*ҷ*�@4:\ߞٿa��Wؙ�@�xa3B�3@�����!? �*ҷ*�@t�.m�ٿŕar��@�s'���3@�2�R��!?�:���M�@t�.m�ٿŕar��@�s'���3@�2�R��!?�:���M�@$��9q�ٿӟ���@�K�3@�sc��!?�����@$��9q�ٿӟ���@�K�3@�sc��!?�����@$��9q�ٿӟ���@�K�3@�sc��!?�����@$��9q�ٿӟ���@�K�3@�sc��!?�����@$��9q�ٿӟ���@�K�3@�sc��!?�����@$��9q�ٿӟ���@�K�3@�sc��!?�����@/]C){�ٿ�'���@�-M�j�3@����!?ld����@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@eѲ��ٿ��+0���@��+���3@��E�ǐ!?BЕBP��@"	�ٿ`NP����@�c���3@��^���!?Ž�/�@"	�ٿ`NP����@�c���3@��^���!?Ž�/�@"	�ٿ`NP����@�c���3@��^���!?Ž�/�@4�;e�ٿF�9���@]R�8V�3@-�QG��!?�+��@4�;e�ٿF�9���@]R�8V�3@-�QG��!?�+��@4�;e�ٿF�9���@]R�8V�3@-�QG��!?�+��@4�;e�ٿF�9���@]R�8V�3@-�QG��!?�+��@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@l�J�ٿ�����@GIҴ�3@U�7�!?9=�����@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@���9Q�ٿ��&\���@	�G�\�3@�8��!?f4���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@�A�>r�ٿ!��:�@��b!�3@��*��!?�:�2���@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@A��'�ٿ0ύz���@놉z�3@�,���!?�K�:5�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@��h��ٿ�"�:dg�@�����3@[e�Z��!?1���X�@u,��ٿ-�Q�to�@�Ee���3@�Վ�!?��$>��@u,��ٿ-�Q�to�@�Ee���3@�Վ�!?��$>��@u,��ٿ-�Q�to�@�Ee���3@�Վ�!?��$>��@u,��ٿ-�Q�to�@�Ee���3@�Վ�!?��$>��@���u�ٿKX+�x�@��8���3@ayrʐ!?��A�@@��̜ٿ&��=��@��v��3@˟�!?������@@��̜ٿ&��=��@��v��3@˟�!?������@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@��O&�ٿ!\���#�@�Q aK�3@5c���!?(((�Zt�@�ZC��ٿ����@V��K�3@;�_��!?j�@\��@�ZC��ٿ����@V��K�3@;�_��!?j�@\��@�ZC��ٿ����@V��K�3@;�_��!?j�@\��@��
�H�ٿ�"O=b��@[��q�3@�-T	�!?9S�M�@��
�H�ٿ�"O=b��@[��q�3@�-T	�!?9S�M�@��
�H�ٿ�"O=b��@[��q�3@�-T	�!?9S�M�@����ٿm�o�L`�@
����3@���	��!?��E��Y�@����ٿm�o�L`�@
����3@���	��!?��E��Y�@��ZWJ�ٿP��jy��@<D���3@ʲ±��!?��A�@��ZWJ�ٿP��jy��@<D���3@ʲ±��!?��A�@��ZWJ�ٿP��jy��@<D���3@ʲ±��!?��A�@��ZWJ�ٿP��jy��@<D���3@ʲ±��!?��A�@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@��+��ٿߵ����@񙗇^�3@�z
V!?�a���@!ٜٿh�B�i�@�X����3@|����!?qi0a��@�l��ٿ��-���@qZ��^�3@��'Ñ�!?��L�r�@�l��ٿ��-���@qZ��^�3@��'Ñ�!?��L�r�@�l��ٿ��-���@qZ��^�3@��'Ñ�!?��L�r�@�l��ٿ��-���@qZ��^�3@��'Ñ�!?��L�r�@�l��ٿ��-���@qZ��^�3@��'Ñ�!?��L�r�@vYM���ٿ���^��@�mD9_�3@�ݢ;m�!?��ǋ��@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@�W���ٿ��ą��@f���e�3@��s��!?�߬��O�@���A�ٿK�|�I�@{ԬC�3@���.��!?�?��A�@���A�ٿK�|�I�@{ԬC�3@���.��!?�?��A�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@Y�;9#�ٿ�Z�-��@��}q��3@D�U�Ő!?���,/�@���m�ٿ��&��@�4�3@�Ov��!?�7���@���m�ٿ��&��@�4�3@�Ov��!?�7���@���m�ٿ��&��@�4�3@�Ov��!?�7���@���m�ٿ��&��@�4�3@�Ov��!?�7���@���m�ٿ��&��@�4�3@�Ov��!?�7���@���m�ٿ��&��@�4�3@�Ov��!?�7���@��J؊�ٿ�_X
%��@�c��3@R9p���!?'�$\�@�����ٿ�	"I�@�.|S�3@㟇��!?=�')`��@�����ٿ�	"I�@�.|S�3@㟇��!?=�')`��@�����ٿ�	"I�@�.|S�3@㟇��!?=�')`��@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@S�ſ��ٿ���r��@Ǖ�O��3@�%@���!?&����@<�}�ٿ��fS�4�@�:�}��3@��ݯ��!?\a��@<�}�ٿ��fS�4�@�:�}��3@��ݯ��!?\a��@<�}�ٿ��fS�4�@�:�}��3@��ݯ��!?\a��@��r;�ٿ*�PM�@4Jl��3@�kA��!?D������@��r;�ٿ*�PM�@4Jl��3@�kA��!?D������@�yEp��ٿz��64�@ޅ����3@�Q�"Ɛ!?���)5��@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@=��
�ٿ{F�}�@��U�4�3@k1�!?���g7�@����I�ٿ�����@.�P&�3@�lP��!?�R��nx�@3U���ٿ���4��@�Ѐ��3@rouŐ!?n�|޸�@3U���ٿ���4��@�Ѐ��3@rouŐ!?n�|޸�@3U���ٿ���4��@�Ѐ��3@rouŐ!?n�|޸�@3U���ٿ���4��@�Ѐ��3@rouŐ!?n�|޸�@q!�˝ٿ"p$����@+!�ئ�3@�b�@�!?���M�
�@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@=D�$C�ٿ������@	�B{�3@�tݐ!?Ac~���@1L&��ٿ�bY/�@��n��3@�� 4Ɛ!?h�-���@�:�]أٿ� ��1�@:�����3@��1�Ð!?}��6�@�:�]أٿ� ��1�@:�����3@��1�Ð!?}��6�@�:�]أٿ� ��1�@:�����3@��1�Ð!?}��6�@�����ٿ-U;R3�@'��W��3@zmi廐!?��^����@u�#��ٿ��:9���@ k��[�3@�[þ�!?����
�@u�#��ٿ��:9���@ k��[�3@�[þ�!?����
�@u�#��ٿ��:9���@ k��[�3@�[þ�!?����
�@7S^��ٿ�ɻs���@����2�3@4e���!?y������@7S^��ٿ�ɻs���@����2�3@4e���!?y������@7S^��ٿ�ɻs���@����2�3@4e���!?y������@7S^��ٿ�ɻs���@����2�3@4e���!?y������@��sRơٿr�>�_�@~ۖs��3@D"!�ʐ!? rT;4��@��sRơٿr�>�_�@~ۖs��3@D"!�ʐ!? rT;4��@�cS��ٿ���F���@5M��L�3@0*�(��!?�,����@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@#�Lݧٿ�P'I���@�Y$ֲ�3@6@�ؐ!?IW;���@t�H�*�ٿ��J)�@h��'�3@LPV���!?�m���@t�H�*�ٿ��J)�@h��'�3@LPV���!?�m���@t�H�*�ٿ��J)�@h��'�3@LPV���!?�m���@t�H�*�ٿ��J)�@h��'�3@LPV���!?�m���@t�H�*�ٿ��J)�@h��'�3@LPV���!?�m���@l�D	.�ٿsI�
�@
�M��3@�����!?�VuԘ��@l�D	.�ٿsI�
�@
�M��3@�����!?�VuԘ��@l�D	.�ٿsI�
�@
�M��3@�����!?�VuԘ��@l�D	.�ٿsI�
�@
�M��3@�����!?�VuԘ��@l�D	.�ٿsI�
�@
�M��3@�����!?�VuԘ��@gNf�ٿER�o��@��E��3@�^?:]�!?�*�>�@gNf�ٿER�o��@��E��3@�^?:]�!?�*�>�@gNf�ٿER�o��@��E��3@�^?:]�!?�*�>�@gNf�ٿER�o��@��E��3@�^?:]�!?�*�>�@����ٿ8�h�y�@W�6�3@����!?�P�x��@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@�:�?��ٿ-c�*	a�@�|4��3@n��Ų�!?3�)����@��ߋ�ٿ�l4����@��!��3@�fϐ!?KE0���@��ߋ�ٿ�l4����@��!��3@�fϐ!?KE0���@��ߋ�ٿ�l4����@��!��3@�fϐ!?KE0���@��
��ٿ���7n��@(.H��3@ǡ'��!?��(���@��
��ٿ���7n��@(.H��3@ǡ'��!?��(���@��
��ٿ���7n��@(.H��3@ǡ'��!?��(���@�I׀W�ٿud�Ť��@����3@��н�!?��q}���@^���ٿm�^B�L�@:�P��3@=��.�!??�ѣx�@��At�ٿ�,�,VX�@�ދ%��3@�CG�ɐ!?P�zUH��@��At�ٿ�,�,VX�@�ދ%��3@�CG�ɐ!?P�zUH��@��At�ٿ�,�,VX�@�ދ%��3@�CG�ɐ!?P�zUH��@ZZ��ٿc��4)%�@�3�5�3@an!���!?��1�o��@ZZ��ٿc��4)%�@�3�5�3@an!���!?��1�o��@ZZ��ٿc��4)%�@�3�5�3@an!���!?��1�o��@ZZ��ٿc��4)%�@�3�5�3@an!���!?��1�o��@ZZ��ٿc��4)%�@�3�5�3@an!���!?��1�o��@�ה�ٿ�\ز���@)~3���3@D���!?y�[r���@�ה�ٿ�\ز���@)~3���3@D���!?y�[r���@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@��E�ٿ��0ϚB�@��{G�3@����!?pt��s��@]��|�ٿ���T�@�7����3@�X�!?p[3�k�@]��|�ٿ���T�@�7����3@�X�!?p[3�k�@3]|�S�ٿS������@{E1,�3@g�(���!?�����@3]|�S�ٿS������@{E1,�3@g�(���!?�����@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@��;�ؤٿ��p���@�����3@:*��!?e���:q�@�2��&�ٿ��0��@�)��3@�3�Đ!?�)���@���je�ٿQ�[;&�@"���3@�IkQ�!?N�3����@���je�ٿQ�[;&�@"���3@�IkQ�!?N�3����@�Q���ٿ�9�YG�@�&���3@7�,z�!?㒹V��@�Q���ٿ�9�YG�@�&���3@7�,z�!?㒹V��@�Q���ٿ�9�YG�@�&���3@7�,z�!?㒹V��@g����ٿG�N��=�@N*�<!�3@ͩ���!?���gB�@g����ٿG�N��=�@N*�<!�3@ͩ���!?���gB�@g����ٿG�N��=�@N*�<!�3@ͩ���!?���gB�@g����ٿG�N��=�@N*�<!�3@ͩ���!?���gB�@5u�n�ٿLO9�r�@��l�3@v_N��!?`��1�@5u�n�ٿLO9�r�@��l�3@v_N��!?`��1�@�l"5��ٿ�aVp��@ӆO�o�3@������!?ӷ����@�l"5��ٿ�aVp��@ӆO�o�3@������!?ӷ����@�l"5��ٿ�aVp��@ӆO�o�3@������!?ӷ����@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@o	3Кٿ�T+a���@cqT �3@�RT&�!?͸|)�*�@쨓�F�ٿn���Ǌ�@,�+5'�3@y�-Xː!?��r��@쨓�F�ٿn���Ǌ�@,�+5'�3@y�-Xː!?��r��@�]�oÞٿ�D�h�@K���3@ڼZ��!?�1R�\��@�]�oÞٿ�D�h�@K���3@ڼZ��!?�1R�\��@��.e��ٿ���O�@%��3@��߶�!?G�E��@��ܟٿ����"�@���6p�3@�Y�ͥ�!?�^���L�@���V��ٿ�΢!�`�@.�q���3@{�G��!?,i��j�@���V��ٿ�΢!�`�@.�q���3@{�G��!?,i��j�@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@���ܞ�ٿ:�����@X�|��3@���!?9	��S��@�U/���ٿ��*��@��$�=�3@�w,�!?�e����@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@ɂ!�q�ٿoΖ\���@�~lt�3@�U����!?�P�匃�@le�ןٿ�&���@ȧk�!�3@��+TŐ!?(�ڭÈ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@ʒ�,�ٿ"Oi�� �@=�J�3@ 	@ڐ!?LoؑQ�@���W�ٿ&ᠸ~��@	Ro�:�3@S�_�!?��w&���@���W�ٿ&ᠸ~��@	Ro�:�3@S�_�!?��w&���@��)?�ٿ�žo��@J� �3�3@C�R�ݐ!?<��tg�@��)?�ٿ�žo��@J� �3�3@C�R�ݐ!?<��tg�@w�g�u�ٿ��P���@nJ�u��3@\,�!?8��qB��@w�g�u�ٿ��P���@nJ�u��3@\,�!?8��qB��@��<�ٿ++2Z��@OX�4�3@����!?]p`m��@��<�ٿ++2Z��@OX�4�3@����!?]p`m��@î���ٿZ�(�|�@/�B�J�3@�7�ϐ!?&$�(��@î���ٿZ�(�|�@/�B�J�3@�7�ϐ!?&$�(��@��6.ƣٿ��;o��@��]� �3@�(Eh��!?LH.AL��@��6.ƣٿ��;o��@��]� �3@�(Eh��!?LH.AL��@��6.ƣٿ��;o��@��]� �3@�(Eh��!?LH.AL��@�E�V��ٿ�}2��@1�X��3@?�&뤐!?�6�B�@�E�V��ٿ�}2��@1�X��3@?�&뤐!?�6�B�@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@�LI�ٿ��S��@H�F�z�3@�l���!?ʋ`����@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@;s�s�ٿ#a~���@<�,���3@=�>a��!?� ��M��@4i͢ٿ,{Jd�!�@t3&��3@�s�:l�!?l~FlK��@4i͢ٿ,{Jd�!�@t3&��3@�s�:l�!?l~FlK��@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��"�ٿrưw4��@�)�y�3@u[W���!?�9�M�@��,㷡ٿ|f�pJy�@US����3@�=����!?Vm�� +�@��,㷡ٿ|f�pJy�@US����3@�=����!?Vm�� +�@��,㷡ٿ|f�pJy�@US����3@�=����!?Vm�� +�@��,㷡ٿ|f�pJy�@US����3@�=����!?Vm�� +�@^����ٿs ��2��@������3@�5�y�!?�$�,s3�@^����ٿs ��2��@������3@�5�y�!?�$�,s3�@^����ٿs ��2��@������3@�5�y�!?�$�,s3�@^����ٿs ��2��@������3@�5�y�!?�$�,s3�@���n�ٿ&����\�@�+[�W�3@��@ⷐ!?m-o���@���n�ٿ&����\�@�+[�W�3@��@ⷐ!?m-o���@���n�ٿ&����\�@�+[�W�3@��@ⷐ!?m-o���@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�6�ٿ�;��'�@���/x�3@|PhQ��!?TG��"S�@�m����ٿ~��:�@G<��"�3@��1�ؐ!?���|�@��u��ٿ�֬��Z�@������3@_W�Ɛ!?^�'����@��u��ٿ�֬��Z�@������3@_W�Ɛ!?^�'����@��u��ٿ�֬��Z�@������3@_W�Ɛ!?^�'����@g�����ٿ�����@-�;���3@��֐!?�(B����@��:�	�ٿJDr�(�@��L�'�3@5�L0��!?��[���@��:�	�ٿJDr�(�@��L�'�3@5�L0��!?��[���@��:�	�ٿJDr�(�@��L�'�3@5�L0��!?��[���@��:�	�ٿJDr�(�@��L�'�3@5�L0��!?��[���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@Ez�B�ٿ���5���@KAqD�3@�u!�!?"2y���@���	�ٿ�Y$0��@���i�3@�3#�!?�r#���@���	�ٿ�Y$0��@���i�3@�3#�!?�r#���@�o���ٿ��Ǣ��@wݱ���3@�;)�Ґ!?vN��k�@�o���ٿ��Ǣ��@wݱ���3@�;)�Ґ!?vN��k�@�o���ٿ��Ǣ��@wݱ���3@�;)�Ґ!?vN��k�@'�#�ٿs����@#\�_�3@v�r� �!?��!�@y���ٿ��L���@�gR�3@W�����!?;�A��@y���ٿ��L���@�gR�3@W�����!?;�A��@y���ٿ��L���@�gR�3@W�����!?;�A��@y���ٿ��L���@�gR�3@W�����!?;�A��@y���ٿ��L���@�gR�3@W�����!?;�A��@�ECs��ٿ1P�4c�@��$��3@�jB�!?�͸x���@������ٿI��L$��@&<c�3@ٯC��!?Mt]�z�@������ٿI��L$��@&<c�3@ٯC��!?Mt]�z�@�����ٿ�y�f��@џ�`�3@3�O�!?����Y��@�����ٿ�y�f��@џ�`�3@3�O�!?����Y��@�����ٿ�y�f��@џ�`�3@3�O�!?����Y��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@����ٿ����n��@CA��3@$]L�ސ!?Ձ��K��@������ٿ:k�o�}�@A����3@
�4�!?a2.}ʤ�@������ٿ:k�o�}�@A����3@
�4�!?a2.}ʤ�@������ٿ:k�o�}�@A����3@
�4�!?a2.}ʤ�@������ٿ:k�o�}�@A����3@
�4�!?a2.}ʤ�@������ٿ:k�o�}�@A����3@
�4�!?a2.}ʤ�@{�M�ٿ�z#�z�@guA���3@��}�ǐ!?c~�7�p�@{�M�ٿ�z#�z�@guA���3@��}�ǐ!?c~�7�p�@{�M�ٿ�z#�z�@guA���3@��}�ǐ!?c~�7�p�@{�M�ٿ�z#�z�@guA���3@��}�ǐ!?c~�7�p�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�n</��ٿ�O{ņ��@ʧ%4D�3@���iĐ!?pn"{JZ�@�{�+q�ٿ���-R(�@��K�3@kԛRq�!?�͸.���@�{�+q�ٿ���-R(�@��K�3@kԛRq�!?�͸.���@�{�+q�ٿ���-R(�@��K�3@kԛRq�!?�͸.���@��Y��ٿhky.���@�*Ո�3@zӎ��!?w0	'��@��Y��ٿhky.���@�*Ո�3@zӎ��!?w0	'��@��Y��ٿhky.���@�*Ո�3@zӎ��!?w0	'��@��Y��ٿhky.���@�*Ո�3@zӎ��!?w0	'��@RÒ�Q�ٿ�,L#�$�@�s$[>�3@7;���!?���S��@RÒ�Q�ٿ�,L#�$�@�s$[>�3@7;���!?���S��@RÒ�Q�ٿ�,L#�$�@�s$[>�3@7;���!?���S��@RÒ�Q�ٿ�,L#�$�@�s$[>�3@7;���!?���S��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@���V��ٿ��W�R �@�4���3@E��Đ!?��J9��@	�^�ٿ��jV�@�;o���3@<�u��!?��'d9��@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@BjG �ٿ��Q�i��@�T����3@0X���!?��:���@��g^A�ٿ��*��@�V���3@�,^���!?�Zĭ��@��g^A�ٿ��*��@�V���3@�,^���!?�Zĭ��@��g^A�ٿ��*��@�V���3@�,^���!?�Zĭ��@��g^A�ٿ��*��@�V���3@�,^���!?�Zĭ��@��g^A�ٿ��*��@�V���3@�,^���!?�Zĭ��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@��D�ٿ���Y7�@�q��3@s>���!?��aGH��@Q�	&I�ٿ�<�x��@{��3@�eA;ؐ!?9A���*�@Q�	&I�ٿ�<�x��@{��3@�eA;ؐ!?9A���*�@Q�	&I�ٿ�<�x��@{��3@�eA;ؐ!?9A���*�@
�*d�ٿ�v��y�@3�Zl�3@e���!?�Ri4���@
�*d�ٿ�v��y�@3�Zl�3@e���!?�Ri4���@�t�	�ٿnA����@-�$�@�3@�	�!?3��c[�@O����ٿ��R���@�j(��3@��#� �!?��]�y�@<q"�ߜٿY���t��@��e��3@ӥR*��!?�pB��1�@<q"�ߜٿY���t��@��e��3@ӥR*��!?�pB��1�@<q"�ߜٿY���t��@��e��3@ӥR*��!?�pB��1�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ&l����@F.kY[�3@I��!?vtϭ�S�@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@����ٿ��Rt]��@A���3@�@<]��!?¸�h���@w�P�8�ٿif�^��@�MB�r�3@=Ğh��!?V��P��@w�P�8�ٿif�^��@�MB�r�3@=Ğh��!?V��P��@�3��D�ٿ�z�2e�@��pZ�3@�^]@��!?��^b��@�3��D�ٿ�z�2e�@��pZ�3@�^]@��!?��^b��@�3��D�ٿ�z�2e�@��pZ�3@�^]@��!?��^b��@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@,�Dѥٿ|���-�@M����3@X�k�Ő!?b�o���@%�H�ٿ`�u��@�c޼�3@\�^��!?{yj�A��@%�H�ٿ`�u��@�c޼�3@\�^��!?{yj�A��@��ŝٿ�oz�g��@{h	!#�3@.�h=��!?�.���@��ŝٿ�oz�g��@{h	!#�3@.�h=��!?�.���@��ŝٿ�oz�g��@{h	!#�3@.�h=��!?�.���@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@�9b�x�ٿkl�t=R�@��B�3@�.��!?�u��D�@T��ٿKT��;�@�,㚝�3@h@ipƐ!?H*�]�@T��ٿKT��;�@�,㚝�3@h@ipƐ!?H*�]�@�iIN1�ٿ�ef�<��@Fba���3@���ǐ!?U����@�k��ٿ�30�N�@xŧ���3@�S�I��!?[P9�#��@�k��ٿ�30�N�@xŧ���3@�S�I��!?[P9�#��@�k��ٿ�30�N�@xŧ���3@�S�I��!?[P9�#��@�k��ٿ�30�N�@xŧ���3@�S�I��!?[P9�#��@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@�c�ʟٿ+����@(���K�3@B�C���!?���f�F�@���Y�ٿ�]#��@��Ӭ��3@�@�KА!?d��]��@���Y�ٿ�]#��@��Ӭ��3@�@�KА!?d��]��@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@�!Λٿ����@�j�0�3@ۢ���!?��7G�S�@� /��ٿ4�q��@��
(�3@�%����!?sŗj)�@lVX�ٿ
$��j�@4�(s��3@෤ɳ�!?N&r���@lVX�ٿ
$��j�@4�(s��3@෤ɳ�!?N&r���@lVX�ٿ
$��j�@4�(s��3@෤ɳ�!?N&r���@lVX�ٿ
$��j�@4�(s��3@෤ɳ�!?N&r���@lVX�ٿ
$��j�@4�(s��3@෤ɳ�!?N&r���@�m����ٿ�=潝u�@�աO�3@ڜz��!?:+[��@�@�m����ٿ�=潝u�@�աO�3@ڜz��!?:+[��@�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@��Rd�ٿYH1���@��9�3@[B�_��!?�����#�@)�qS\�ٿ�$ë�0�@w���
�3@����!?;�\���@)�qS\�ٿ�$ë�0�@w���
�3@����!?;�\���@)�qS\�ٿ�$ë�0�@w���
�3@����!?;�\���@)�qS\�ٿ�$ë�0�@w���
�3@����!?;�\���@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@m⭬�ٿ��Àl�@e0?���3@�����!?I����e�@��/�ٿ�0�_���@�#�>6�3@��,�!?5v��mw�@��/�ٿ�0�_���@�#�>6�3@��,�!?5v��mw�@U6C1�ٿc�@��@O���3@��^X(�!?��v竴�@��	��ٿk�7O�V�@زzP�3@���� �!?|=x �-�@��	��ٿk�7O�V�@زzP�3@���� �!?|=x �-�@��	��ٿk�7O�V�@زzP�3@���� �!?|=x �-�@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@̡�?�ٿ�i���K�@ă{6�3@�ݸb�!?��e�:��@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@(̥��ٿg�sX)��@�AaR��3@׈d�Ð!?G�|���@e���0�ٿ�L����@��+�3@���D�!?B�	���@�	^�ڛٿ@o6�x2�@|SPs_�3@a��o�!?i�N/���@�t�ٿ͛Wơ�@?�;�3@��J���!?O��H���@�q�i�ٿ(�W��6�@�W��3@#E�|��!?WD*I'��@�q�i�ٿ(�W��6�@�W��3@#E�|��!?WD*I'��@�q�i�ٿ(�W��6�@�W��3@#E�|��!?WD*I'��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@M��>�ٿ��C5u��@�bE��3@�6�Cy�!?3B�P��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@z��A�ٿ�K�h�~�@�����3@�@k㉐!?Aw*�1��@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@�oÛ��ٿz�,}�@��*;�3@���Y�!?+���ϋ�@��4o�ٿ�!�4��@���z�3@�ߡ�!?3s��U�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�"
{��ٿ��=#�@XzK%@�3@��Vڐ!?����W�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�ERx��ٿ�f�	 a�@pKm�h�3@ ��x��!?���z�@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@�7�Mx�ٿ���)���@L�����3@ �hӐ!?�"�����@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@L�*�ٿ[tܾW|�@�WXp�3@�G7!?0,�-�@�Ct��ٿ	y�����@��{��3@��C��!?��i��.�@�Ct��ٿ	y�����@��{��3@��C��!?��i��.�@��9�ٿ���+�@W~[:�3@��Zߐ!?��}u9r�@��9�ٿ���+�@W~[:�3@��Zߐ!?��}u9r�@��9�ٿ���+�@W~[:�3@��Zߐ!?��}u9r�@��>h�ٿ,|�ݨ�@tx�G��3@c�!?W��C��@��>h�ٿ,|�ݨ�@tx�G��3@c�!?W��C��@��>h�ٿ,|�ݨ�@tx�G��3@c�!?W��C��@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@�>�?��ٿ�ȹ�m�@N	��3@7����!?�NR���@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@%��ѡٿ=&
e:�@s��&a�3@��a���!?�P/�)�@��ؼ�ٿ�g��ny�@�DK��3@�R=%��!?��$��/�@խ�Sv�ٿ���=���@�ɧ
��3@�i���!?�햴��@խ�Sv�ٿ���=���@�ɧ
��3@�i���!?�햴��@խ�Sv�ٿ���=���@�ɧ
��3@�i���!?�햴��@խ�Sv�ٿ���=���@�ɧ
��3@�i���!?�햴��@�}��T�ٿ��T7q�@�Q���3@���!?�7W����@�}��T�ٿ��T7q�@�Q���3@���!?�7W����@�}��T�ٿ��T7q�@�Q���3@���!?�7W����@�}��T�ٿ��T7q�@�Q���3@���!?�7W����@�Q���ٿ�����@�Ð���3@��َې!?&H�n��@=M۸�ٿ�J��l��@� ���3@,7<�Đ!?��̫���@=M۸�ٿ�J��l��@� ���3@,7<�Đ!?��̫���@G��6�ٿ5�$��@����3@�x���!?���&��@��۩��ٿ��פ���@��f,�3@Z
ӫ�!?�Y�����@��۩��ٿ��פ���@��f,�3@Z
ӫ�!?�Y�����@��۩��ٿ��פ���@��f,�3@Z
ӫ�!?�Y�����@��۩��ٿ��פ���@��f,�3@Z
ӫ�!?�Y�����@��۩��ٿ��פ���@��f,�3@Z
ӫ�!?�Y�����@n�6��ٿ箄��@���g�3@彵���!?���9o�@6a$�ٿ���E�@)��K�3@;�d���!?�낶���@6a$�ٿ���E�@)��K�3@;�d���!?�낶���@6a$�ٿ���E�@)��K�3@;�d���!?�낶���@@X� �ٿT9�|�@-���n�3@�˼��!?��o�i�@����ͧٿ�ꨲ��@��(j��3@�ۢa�!?�X�4sO�@����ͧٿ�ꨲ��@��(j��3@�ۢa�!?�X�4sO�@h/ș	�ٿ9	�5�0�@Tn�p��3@�R�֐!?�C%��=�@h/ș	�ٿ9	�5�0�@Tn�p��3@�R�֐!?�C%��=�@h/ș	�ٿ9	�5�0�@Tn�p��3@�R�֐!?�C%��=�@h/ș	�ٿ9	�5�0�@Tn�p��3@�R�֐!?�C%��=�@h/ș	�ٿ9	�5�0�@Tn�p��3@�R�֐!?�C%��=�@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@������ٿJ�H��@M�r{�3@��Ȑ!?��90���@�O'��ٿ�C�8�@�!m�S�3@�R�֐!?�N#����@�O'��ٿ�C�8�@�!m�S�3@�R�֐!?�N#����@�O'��ٿ�C�8�@�!m�S�3@�R�֐!?�N#����@�O'��ٿ�C�8�@�!m�S�3@�R�֐!?�N#����@�'�s9�ٿo1����@�?��X�3@ڈñ��!?Zw�C��@�'�s9�ٿo1����@�?��X�3@ڈñ��!?Zw�C��@�'�s9�ٿo1����@�?��X�3@ڈñ��!?Zw�C��@�'�s9�ٿo1����@�?��X�3@ڈñ��!?Zw�C��@�#��ٿ�y����@�MM��3@�eS�!?K�Sě�@�#��ٿ�y����@�MM��3@�eS�!?K�Sě�@�#��ٿ�y����@�MM��3@�eS�!?K�Sě�@�#��ٿ�y����@�MM��3@�eS�!?K�Sě�@Յn��ٿ)���r��@�x�&�3@@#iR
�!?�f�{ڹ�@(��5��ٿ�����@FB���3@��J�!?�M��j��@(��5��ٿ�����@FB���3@��J�!?�M��j��@θֆv�ٿW?7��@_��$��3@݊��!?`ᘮ���@θֆv�ٿW?7��@_��$��3@݊��!?`ᘮ���@θֆv�ٿW?7��@_��$��3@݊��!?`ᘮ���@θֆv�ٿW?7��@_��$��3@݊��!?`ᘮ���@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�	P�R�ٿwYk�S�@�;�l��3@���Ր!?�{Ofad�@�\��k�ٿ]V�$���@������3@<��ŧ�!?��xt�Y�@�p3��ٿ:�(���@Z�ϋ#�3@Ǥ4�ѐ!?���K�@�{�E�ٿ�~2��*�@w�ğ��3@y
�T�!?��� ��@2t�?��ٿ�P̂�@��@��3@s�Oz��!?>XH����@��Q@�ٿ�&~Q�@�6�T��3@�q��!?Za��z��@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@��\쯠ٿ4����@މ�G�3@��u⺐!?��Ѫ�@�`��}�ٿ$>�]`��@d�IU�3@�9�!?w�&H��@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@���Y*�ٿ�~ɢ�@ߋr>��3@{�Y� �!?\d���@��Hv.�ٿaO:-R��@��4�8�3@��"��!?�n��;��@��Hv.�ٿaO:-R��@��4�8�3@��"��!?�n��;��@��Hv.�ٿaO:-R��@��4�8�3@��"��!?�n��;��@^W��H�ٿ��kܺ	�@��ܫ��3@�1U|��!?�ZD}�@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@w3�Vw�ٿ.��<��@`L�L*�3@m����!?������@쨝&�ٿ�Q�v��@��(1�3@ NK�!?[:�/��@쨝&�ٿ�Q�v��@��(1�3@ NK�!?[:�/��@8p�E�ٿ�g8��5�@��uQ��3@���W��!?�#�H���@8p�E�ٿ�g8��5�@��uQ��3@���W��!?�#�H���@[=6ϟٿ�H�X���@���Zy�3@�Kw��!?Sp����@��X�5�ٿ���k��@�#�r�3@�D���!?̠���t�@��X�5�ٿ���k��@�#�r�3@�D���!?̠���t�@��X�5�ٿ���k��@�#�r�3@�D���!?̠���t�@��X�5�ٿ���k��@�#�r�3@�D���!?̠���t�@��X�5�ٿ���k��@�#�r�3@�D���!?̠���t�@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@W���ٿ�\:w���@_�]�_�3@�@��!?y*z4��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�����ٿ��Y2�@}j��3@a0df��!?��k��@�A�1��ٿubt���@�k�i�3@֗�nȐ!?u3m�5�@�A�1��ٿubt���@�k�i�3@֗�nȐ!?u3m�5�@�A�1��ٿubt���@�k�i�3@֗�nȐ!?u3m�5�@���8Ϡٿ��"�/^�@�W�a�3@	���!?�/I�I��@���8Ϡٿ��"�/^�@�W�a�3@	���!?�/I�I��@���8Ϡٿ��"�/^�@�W�a�3@	���!?�/I�I��@���})�ٿtS�&�5�@�w?1��3@	����!?���:�@���})�ٿtS�&�5�@�w?1��3@	����!?���:�@���})�ٿtS�&�5�@�w?1��3@	����!?���:�@���})�ٿtS�&�5�@�w?1��3@	����!?���:�@���})�ٿtS�&�5�@�w?1��3@	����!?���:�@`0h�b�ٿp���Z�@���3@���!?�Ha���@`0h�b�ٿp���Z�@���3@���!?�Ha���@Y��5z�ٿ�k�@��@�3Ԓ�3@�a{�Ր!?���|h�@Y��5z�ٿ�k�@��@�3Ԓ�3@�a{�Ր!?���|h�@fy�K�ٿ,��p���@�QE�I�3@6V�_��!?��;���@fy�K�ٿ,��p���@�QE�I�3@6V�_��!?��;���@fy�K�ٿ,��p���@�QE�I�3@6V�_��!?��;���@fy�K�ٿ,��p���@�QE�I�3@6V�_��!?��;���@T�Xc��ٿ��L��`�@�+B^&�3@
��+��!?	tq$��@��qۑ�ٿ�|9d �@ ��3��3@� ؐ!?8�����@��qۑ�ٿ�|9d �@ ��3��3@� ؐ!?8�����@��qۑ�ٿ�|9d �@ ��3��3@� ؐ!?8�����@��qۑ�ٿ�|9d �@ ��3��3@� ؐ!?8�����@(L̑�ٿ���.��@Y���3@)(���!?��"��z�@(L̑�ٿ���.��@Y���3@)(���!?��"��z�@(L̑�ٿ���.��@Y���3@)(���!?��"��z�@ws���ٿ�&���M�@��^�3@*���!?9.�2}�@1�N��ٿZJU���@�q�f�3@ڟ�	�!?՞~g#n�@�Lޛ��ٿGAg,s�@3^�t �3@�[���!?ns����@��Q6�ٿ�8SR���@�a5�$�3@����!?54��B��@��Q6�ٿ�8SR���@�a5�$�3@����!?54��B��@���<��ٿ�ר��@j�N![�3@�0(�Ő!?/�z�H�@���<��ٿ�ר��@j�N![�3@�0(�Ő!?/�z�H�@���/�ٿ��fxz7�@�����3@��7𢡄!?,�����@���/�ٿ��fxz7�@�����3@��7𢡄!?,�����@���/�ٿ��fxz7�@�����3@��7𢡄!?,�����@���/�ٿ��fxz7�@�����3@��7𢡄!?,�����@���/�ٿ��fxz7�@�����3@��7𢡄!?,�����@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�oTU�ٿ�S�
b%�@x��3@v�!��!?��w׻�@�a �ٿ���+F��@~�
��3@Ǩ����!?�Y����@�a �ٿ���+F��@~�
��3@Ǩ����!?�Y����@�a �ٿ���+F��@~�
��3@Ǩ����!?�Y����@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@��*~��ٿ�����`�@��1��3@5�'�n�!?q��`a��@YX��h�ٿ2��Կ�@M��3@���a}�!?=C��7#�@YX��h�ٿ2��Կ�@M��3@���a}�!?=C��7#�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@TSrlo�ٿ�OP
��@c.śg�3@�kN���!?HK��G�@R��^�ٿο��	��@��7.8�3@!x�֐!?�&��?�@R��^�ٿο��	��@��7.8�3@!x�֐!?�&��?�@R��^�ٿο��	��@��7.8�3@!x�֐!?�&��?�@R��^�ٿο��	��@��7.8�3@!x�֐!?�&��?�@h���ٿ(I�U��@��B6�3@����!?�S�#���@h���ٿ(I�U��@��B6�3@����!?�S�#���@ZMZ6@�ٿ�^�ۢ��@�0���3@c���!?�jH��@ZMZ6@�ٿ�^�ۢ��@�0���3@c���!?�jH��@�V���ٿ��Qs���@
��"��3@�E4-!?�Mu&�@�:F�t�ٿ��h��(�@0�V��3@`!�V��!?���:���@�:F�t�ٿ��h��(�@0�V��3@`!�V��!?���:���@*�6�P�ٿ�w#�]��@>y�q�3@=��rl�!?��^�eK�@*�6�P�ٿ�w#�]��@>y�q�3@=��rl�!?��^�eK�@*�6�P�ٿ�w#�]��@>y�q�3@=��rl�!?��^�eK�@*�6�P�ٿ�w#�]��@>y�q�3@=��rl�!?��^�eK�@*�6�P�ٿ�w#�]��@>y�q�3@=��rl�!?��^�eK�@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@p�]�ٿg8�����@���>��3@�T$��!?��P�2��@�"QW��ٿ��M�֞�@����3@q�*�!?�5AV�@�"QW��ٿ��M�֞�@����3@q�*�!?�5AV�@�"QW��ٿ��M�֞�@����3@q�*�!?�5AV�@��F�B�ٿ����Z�@�R��3�3@E0:1$�!?/��<���@��F�B�ٿ����Z�@�R��3�3@E0:1$�!?/��<���@��F�B�ٿ����Z�@�R��3�3@E0:1$�!?/��<���@��F�B�ٿ����Z�@�R��3�3@E0:1$�!?/��<���@dh����ٿE�T���@������3@|7m��!?�R�	'�@dh����ٿE�T���@������3@|7m��!?�R�	'�@dh����ٿE�T���@������3@|7m��!?�R�	'�@dh����ٿE�T���@������3@|7m��!?�R�	'�@�`3�ٿ:��c\h�@���#�3@o"e��!?2�Jި��@��?�r�ٿ*2��j�@��~��3@����ؐ!?+lX.��@ۿ E�ٿ2����/�@�<,z�3@]�b��!?�N\#��@ۿ E�ٿ2����/�@�<,z�3@]�b��!?�N\#��@ۿ E�ٿ2����/�@�<,z�3@]�b��!?�N\#��@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�38m4�ٿ!����@��'�3@)�T�!?��S:=�@�.�b$�ٿ$76��@51�X��3@�\t\q�!?���0y�@�.�b$�ٿ$76��@51�X��3@�\t\q�!?���0y�@�.�b$�ٿ$76��@51�X��3@�\t\q�!?���0y�@�.�b$�ٿ$76��@51�X��3@�\t\q�!?���0y�@�����ٿ�����H�@~>#���3@�Ǵ~�!?�~��2�@�����ٿ���@$�@��Y#� 4@Sl����!?uK�P�[�@�����ٿ���@$�@��Y#� 4@Sl����!?uK�P�[�@�����ٿ���@$�@��Y#� 4@Sl����!?uK�P�[�@�����ٿ���@$�@��Y#� 4@Sl����!?uK�P�[�@�����ٿ���@$�@��Y#� 4@Sl����!?uK�P�[�@��ٲ�ٿ�tU���@)�����3@UU&�!?L
I���@��ٲ�ٿ�tU���@)�����3@UU&�!?L
I���@��ٲ�ٿ�tU���@)�����3@UU&�!?L
I���@"s�&�ٿ%v7�|��@b���3@D���!?�<�_�@"s�&�ٿ%v7�|��@b���3@D���!?�<�_�@k���r�ٿY���~2�@�.\�3@�f7��!?Cb�;/�@k���r�ٿY���~2�@�.\�3@�f7��!?Cb�;/�@k���r�ٿY���~2�@�.\�3@�f7��!?Cb�;/�@.��c�ٿ����@�|I	#�3@_d&���!?�3����@.��c�ٿ����@�|I	#�3@_d&���!?�3����@.��c�ٿ����@�|I	#�3@_d&���!?�3����@.��c�ٿ����@�|I	#�3@_d&���!?�3����@`5d�G�ٿa"3�=��@L�+?�3@W5�ګ�!?��5DYF�@x̵���ٿ(L�:���@ާ����3@D�S#�!?�i��o�@x̵���ٿ(L�:���@ާ����3@D�S#�!?�i��o�@x̵���ٿ(L�:���@ާ����3@D�S#�!?�i��o�@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@z�."�ٿ)e��u�@͖ly�3@��xT+�!?�����@*��Q_�ٿ���S�@��{��3@�?eT0�!?8\t�@&yk=�ٿ�Pn�r��@��xCq�3@��Đ!?c�M�@&yk=�ٿ�Pn�r��@��xCq�3@��Đ!?c�M�@&yk=�ٿ�Pn�r��@��xCq�3@��Đ!?c�M�@&yk=�ٿ�Pn�r��@��xCq�3@��Đ!?c�M�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@����ٿ�9�K[��@����3@�O`IА!?�8���}�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@]lK��ٿ]����@x2�0�3@�"(ސ!?��� �{�@��j  �ٿ@�Y�_�@��J@C�3@��ҳ��!?��}�Q��@���P��ٿ������@��Z2M�3@Gs��!?S�@����@���P��ٿ������@��Z2M�3@Gs��!?S�@����@\�̕��ٿ]��P���@Qj��3@Ӵ��!?�X�J(�@\�̕��ٿ]��P���@Qj��3@Ӵ��!?�X�J(�@\�̕��ٿ]��P���@Qj��3@Ӵ��!?�X�J(�@\�̕��ٿ]��P���@Qj��3@Ӵ��!?�X�J(�@\�̕��ٿ]��P���@Qj��3@Ӵ��!?�X�J(�@h^���ٿ�#ظ��@��6��3@\���!?�L�|P��@Ef�>�ٿ�
�qO�@5�p���3@�x�5ݐ!?��'m��@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@���#�ٿ��a�U��@adXa��3@���\Ґ!?Е[���@.���ٿ+�\��U�@�b��g�3@�>���!?naA���@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@���詢ٿ��	_�@���7�3@,�f-��!?�Z��Lm�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@��<�+�ٿ�W|��J�@��f�*�3@w,`|�!?5s�S/�@nVPEm�ٿ~��ܥ��@������3@y��!?��Z�a9�@nVPEm�ٿ~��ܥ��@������3@y��!?��Z�a9�@nVPEm�ٿ~��ܥ��@������3@y��!?��Z�a9�@nVPEm�ٿ~��ܥ��@������3@y��!?��Z�a9�@nVPEm�ٿ~��ܥ��@������3@y��!?��Z�a9�@$�W�-�ٿ��e�S��@de�a�3@����<�!?�_���@$�W�-�ٿ��e�S��@de�a�3@����<�!?�_���@$�W�-�ٿ��e�S��@de�a�3@����<�!?�_���@$�W�-�ٿ��e�S��@de�a�3@����<�!?�_���@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@�mAJ��ٿ���@6�.2C�3@��^��!?��)��@&�����ٿm�%oC�@��\q��3@p {W��!?�?�v�@&�����ٿm�%oC�@��\q��3@p {W��!?�?�v�@8��0�ٿ",X�u��@1a�'��3@��fn��!?�rap�5�@8��0�ٿ",X�u��@1a�'��3@��fn��!?�rap�5�@xdM:C�ٿ:ܵHHK�@V�}���3@|9����!?�s#�)��@�6�&x�ٿ2���Rt�@-�h�y�3@�9>�ڐ!?R���`V�@��O�ġٿOf�;���@�
|���3@5?�g�!?���+���@��O�ġٿOf�;���@�
|���3@5?�g�!?���+���@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@)	"�ףٿ-�b��@�)���3@�0ʖ�!?�6�آ��@�L �ٿ}Ŝu�)�@^����3@wI�[��!?�].���@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�L20�ٿa�Ӳs�@r���3@5�<��!?��h�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@�҈�ٿ�Mk�i�@��LY��3@�.�Ȑ!?ĜH�9�@��-��ٿ�}��C�@8?�s��3@�_�f��!?e��@��-��ٿ�}��C�@8?�s��3@�_�f��!?e��@��-��ٿ�}��C�@8?�s��3@�_�f��!?e��@��-��ٿ�}��C�@8?�s��3@�_�f��!?e��@��-��ٿ�}��C�@8?�s��3@�_�f��!?e��@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�F�	ʜٿ��:4Q��@4��!��3@��ߐ!?T6�~�@�a�D�ٿ�*��"w�@=ܬ�j�3@gN4c�!?��y��@��؛ٿ�>}�_x�@��M�3@�B��!?i&I��R�@��؛ٿ�>}�_x�@��M�3@�B��!?i&I��R�@��؛ٿ�>}�_x�@��M�3@�B��!?i&I��R�@{�i�p�ٿP�3Vb�@h�G�\�3@�w����!?3/]~��@{�i�p�ٿP�3Vb�@h�G�\�3@�w����!?3/]~��@J΁S�ٿŝ�f�@27�ԇ�3@y�]3�!?I&4��!�@J΁S�ٿŝ�f�@27�ԇ�3@y�]3�!?I&4��!�@J΁S�ٿŝ�f�@27�ԇ�3@y�]3�!?I&4��!�@J΁S�ٿŝ�f�@27�ԇ�3@y�]3�!?I&4��!�@����a�ٿ�Gݡ�X�@�Bk`�3@���'�!?���v�@����a�ٿ�Gݡ�X�@�Bk`�3@���'�!?���v�@����a�ٿ�Gݡ�X�@�Bk`�3@���'�!?���v�@��e�ٞٿC'���T�@f�D���3@�S{r��!?yK�ܥX�@��e�ٞٿC'���T�@f�D���3@�S{r��!?yK�ܥX�@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@���5�ٿ�w3�z �@�.��3@͏r�Ȑ!?�����@��v�4�ٿi�?z�$�@���(�3@薉���!?K����s�@Y���F�ٿ��y�_(�@�<&�8�3@�xT��!?�yÍ���@Y���F�ٿ��y�_(�@�<&�8�3@�xT��!?�yÍ���@�|����ٿ�Q����@��G��3@�7���!?r`���{�@�|����ٿ�Q����@��G��3@�7���!?r`���{�@L@�D��ٿ�yg�T�@�V"���3@��TȐ!?�=	VH�@L@�D��ٿ�yg�T�@�V"���3@��TȐ!?�=	VH�@��t{}�ٿO�&x�O�@;���)�3@��؁�!?Xi�KW�@�ĺ��ٿb��Av�@@`jV�3@������!?���8%��@�ĺ��ٿb��Av�@@`jV�3@������!?���8%��@�ĺ��ٿb��Av�@@`jV�3@������!?���8%��@�ĺ��ٿb��Av�@@`jV�3@������!?���8%��@��9��ٿ�e�[N�@�����3@��h谐!?n�����@��9��ٿ�e�[N�@�����3@��h谐!?n�����@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�=֯��ٿo©E/�@?�.�� 4@��m��!?EIn1w�@�QD��ٿ��@�b��@�Qm��4@���IZ�!?@��9��@w�wХٿ���l}�@�ou|��3@�Ve�!?h��%��@�����ٿ�|n�F�@d�m4@�	��^�!?e��0�@�����ٿ�|n�F�@d�m4@�	��^�!?e��0�@�����ٿ�|n�F�@d�m4@�	��^�!?e��0�@�����ٿ�|n�F�@d�m4@�	��^�!?e��0�@�����ٿ�|n�F�@d�m4@�	��^�!?e��0�@3h�Ћ�ٿ�I/����@�ި�C�3@�8��!?y%����@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@�ć��ٿ5mf�w�@p�3L\�3@:�G}ѐ!?�{��b��@A\a��ٿ�ȏڑ�@�6|��3@THTې!?g�u���@A\a��ٿ�ȏڑ�@�6|��3@THTې!?g�u���@�j�M3�ٿ4�].��@��DH�3@�.ͮ�!?��h�H��@�j�M3�ٿ4�].��@��DH�3@�.ͮ�!?��h�H��@�j�M3�ٿ4�].��@��DH�3@�.ͮ�!?��h�H��@���ֆ�ٿJm�S�@y�g8}�3@�7 �d�!?̀�5���@���ֆ�ٿJm�S�@y�g8}�3@�7 �d�!?̀�5���@���ֆ�ٿJm�S�@y�g8}�3@�7 �d�!?̀�5���@��8e �ٿ��u
��@�+���3@��0�!?`+���@��8e �ٿ��u
��@�+���3@��0�!?`+���@��8e �ٿ��u
��@�+���3@��0�!?`+���@��8e �ٿ��u
��@�+���3@��0�!?`+���@��8e �ٿ��u
��@�+���3@��0�!?`+���@�@n�@�ٿ�]JE��@o�yx�3@�pP�S�!?������@�@n�@�ٿ�]JE��@o�yx�3@�pP�S�!?������@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@1sÆN�ٿdMYa�@y�ƀ�3@�x��A�!?	��93��@�x�h�ٿ��n�iG�@���>�3@��ț��!?�������@�x�h�ٿ��n�iG�@���>�3@��ț��!?�������@��@��ٿ@Y�M��@^�<Y(�3@�`Au�!?�o�ӎ/�@��@��ٿ@Y�M��@^�<Y(�3@�`Au�!?�o�ӎ/�@윊�C�ٿ`��\�>�@#�$���3@�1�А!?���$�^�@윊�C�ٿ`��\�>�@#�$���3@�1�А!?���$�^�@윊�C�ٿ`��\�>�@#�$���3@�1�А!?���$�^�@윊�C�ٿ`��\�>�@#�$���3@�1�А!?���$�^�@윊�C�ٿ`��\�>�@#�$���3@�1�А!?���$�^�@��zg�ٿ6�8
���@c�
��3@s�A0��!?�[&yʸ�@��zg�ٿ6�8
���@c�
��3@s�A0��!?�[&yʸ�@��zg�ٿ6�8
���@c�
��3@s�A0��!?�[&yʸ�@��zg�ٿ6�8
���@c�
��3@s�A0��!?�[&yʸ�@��zg�ٿ6�8
���@c�
��3@s�A0��!?�[&yʸ�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@y݇���ٿ������@5�� �3@�<��{�!?Pe2)sp�@*�n]��ٿ�>�H���@��>�3@�E	Þ�!?c�uDd��@jMX�ٿv � ���@��F_�3@�)*��!?�/
�b��@jMX�ٿv � ���@��F_�3@�)*��!?�/
�b��@jMX�ٿv � ���@��F_�3@�)*��!?�/
�b��@��y�0�ٿ|��R��@8��]�3@gϼ'��!?�\k��<�@��y�0�ٿ|��R��@8��]�3@gϼ'��!?�\k��<�@��y�0�ٿ|��R��@8��]�3@gϼ'��!?�\k��<�@��y�0�ٿ|��R��@8��]�3@gϼ'��!?�\k��<�@��y�0�ٿ|��R��@8��]�3@gϼ'��!?�\k��<�@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@G�<ǟٿ���%�@9�О��3@�q`?�!?#x�M��@CT��Οٿg��l3��@Vd�%�3@Q {Ð!?@>�Hu�@CT��Οٿg��l3��@Vd�%�3@Q {Ð!?@>�Hu�@���<�ٿ-KH�-"�@6�i�3@�[ָ��!?J.��@���<�ٿ-KH�-"�@6�i�3@�[ָ��!?J.��@���<�ٿ-KH�-"�@6�i�3@�[ָ��!?J.��@���<�ٿ-KH�-"�@6�i�3@�[ָ��!?J.��@���<�ٿ-KH�-"�@6�i�3@�[ָ��!?J.��@�߰4�ٿ�����@*�T
��3@E��~�!?��*�Z�@�߰4�ٿ�����@*�T
��3@E��~�!?��*�Z�@�߰4�ٿ�����@*�T
��3@E��~�!?��*�Z�@�߰4�ٿ�����@*�T
��3@E��~�!?��*�Z�@��E[��ٿfx3C�(�@���LR�3@޹aC�!? 4����@��E[��ٿfx3C�(�@���LR�3@޹aC�!? 4����@��E[��ٿfx3C�(�@���LR�3@޹aC�!? 4����@�D�&��ٿ��	��@�v�*�3@��x`�!?�u�w F�@�D�&��ٿ��	��@�v�*�3@��x`�!?�u�w F�@�D�&��ٿ��	��@�v�*�3@��x`�!?�u�w F�@��W�ٿ	b��@\h7C��3@���fi�!?\�[�W�@��W�ٿ	b��@\h7C��3@���fi�!?\�[�W�@��W�ٿ	b��@\h7C��3@���fi�!?\�[�W�@v�Cr�ٿT�&K��@`g,Ef�3@��═!?�n2��\�@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@��, �ٿ־~�f5�@�
AƎ�3@���tѐ!?�&�ٗ��@ �;��ٿ�'� �@6�>�3@�YѺ*�!?δ��2�@ �;��ٿ�'� �@6�>�3@�YѺ*�!?δ��2�@ �;��ٿ�'� �@6�>�3@�YѺ*�!?δ��2�@ �;��ٿ�'� �@6�>�3@�YѺ*�!?δ��2�@˪���ٿ�?��n#�@S\�K�3@�Iv��!?{�Łpx�@˪���ٿ�?��n#�@S\�K�3@�Iv��!?{�Łpx�@˪���ٿ�?��n#�@S\�K�3@�Iv��!?{�Łpx�@˪���ٿ�?��n#�@S\�K�3@�Iv��!?{�Łpx�@˪���ٿ�?��n#�@S\�K�3@�Iv��!?{�Łpx�@�9�s�ٿ'YX(��@B��j��3@�0�Đ!?�{����@�9�s�ٿ'YX(��@B��j��3@�0�Đ!?�{����@�9�s�ٿ'YX(��@B��j��3@�0�Đ!?�{����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@n�h��ٿ2�ǨTH�@qd��3@�'a��!?�+�����@]j�&�ٿ=�Ryg�@�:V�r�3@��r���!?��k�]h�@jJބ�ٿ�9�s�+�@,�!�3@!��/��!?�UK�j�@��\Üٿ�Y�=�@�FjCe�3@�q맡�!?�t7T�@��\Üٿ�Y�=�@�FjCe�3@�q맡�!?�t7T�@��\Üٿ�Y�=�@�FjCe�3@�q맡�!?�t7T�@��\Üٿ�Y�=�@�FjCe�3@�q맡�!?�t7T�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@����ٿ��L�@�Sڅf�3@��׆ؐ!?y�<�zL�@��7
�ٿ ο?��@���CU�3@f����!?���Y<p�@��7
�ٿ ο?��@���CU�3@f����!?���Y<p�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�؇���ٿk���`z�@�����3@�:͏�!?ΘŊ_�@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@�f���ٿ���,��@:����3@\W�	А!?�������@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@���ر�ٿ�B�n��@w�#��3@V!l��!?bm��Gq�@�8a���ٿ٪��]��@� ���3@�sxaː!?��4mh�@�8a���ٿ٪��]��@� ���3@�sxaː!?��4mh�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@9���ٿj|@s��@).+���3@XL�踐!?��	�t�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@U�9V��ٿt����@5�n,�3@�v�Jɐ!?:K��&�@�ЮBޗٿ �b��@��/�3@OWF�Ր!?�؅��t�@�ЮBޗٿ �b��@��/�3@OWF�Ր!?�؅��t�@�ЮBޗٿ �b��@��/�3@OWF�Ր!?�؅��t�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@ka�H�ٿ�DXg��@SP#r�3@m��@Ӑ!?�S�)r�@`�6�ٿ��T�)�@<����3@X���!?� ����@`�6�ٿ��T�)�@<����3@X���!?� ����@>R2�>�ٿ�j7,�{�@7ʈP4@6_����!?���w!��@
)?��ٿ;��w{�@E�~��3@'��\��!?�5���@
)?��ٿ;��w{�@E�~��3@'��\��!?�5���@
)?��ٿ;��w{�@E�~��3@'��\��!?�5���@���C�ٿ��w��Q�@{�0�3@V��U�!?f��X'�@K@���ٿ�T�O��@u{SҀ�3@ݣA��!?jS��@K@���ٿ�T�O��@u{SҀ�3@ݣA��!?jS��@.7?sܛٿ�֎;2��@�\5<��3@�����!?�c����@.7?sܛٿ�֎;2��@�\5<��3@�����!?�c����@.7?sܛٿ�֎;2��@�\5<��3@�����!?�c����@��xD��ٿ�����@8xA?��3@tE��!?���
��@��xD��ٿ�����@8xA?��3@tE��!?���
��@��xD��ٿ�����@8xA?��3@tE��!?���
��@1܍�=�ٿ$6�ׅ�@��0�3@�����!?�-��@1܍�=�ٿ$6�ׅ�@��0�3@�����!?�-��@1܍�=�ٿ$6�ׅ�@��0�3@�����!?�-��@e�����ٿ��1�@&!�f��3@^�k��!?�$Q���@e�����ٿ��1�@&!�f��3@^�k��!?�$Q���@e�����ٿ��1�@&!�f��3@^�k��!?�$Q���@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@k�)}�ٿ��=c#%�@ڥM&c�3@Ґ�A��!?d`?��{�@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@Tā�ٿ��X��'�@��-z�3@TLf��!?tԧv���@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@���䜘ٿ2y����@#g5u�3@�m��!?[9��3��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@-�0�G�ٿ�s�	��@��x�E�3@
�J��!?@\�B��@������ٿp�&R��@ƟK��3@�A��!?<�����@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@��X�ٿ�lBqĔ�@�R	L,�3@��i��!?y���]��@&?�4�ٿ����ķ�@,RY��3@2�\�'�!?���@=Kї;�ٿ���X?[�@����W�3@�7$��!?H*Չ��@�j'��ٿ�n�{�@��|��3@�����!?k�ER!��@�j'��ٿ�n�{�@��|��3@�����!?k�ER!��@���wW�ٿ}z��h�@�L1��3@Js�ڐ!?�u}^s��@��)�ϡٿ�0����@��C�3@����!?	�����@��)�ϡٿ�0����@��C�3@����!?	�����@��)�ϡٿ�0����@��C�3@����!?	�����@��)�ϡٿ�0����@��C�3@����!?	�����@��)�ϡٿ�0����@��C�3@����!?	�����@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�s)|U�ٿɂ��M^�@����3@|>��Ґ!?��)���@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�rm~�ٿ6�����@*H���3@=�Jt�!?��:�t�@�`�;�ٿ�j�#���@�KI*��3@4̐!?5}���B�@�`�;�ٿ�j�#���@�KI*��3@4̐!?5}���B�@�`�;�ٿ�j�#���@�KI*��3@4̐!?5}���B�@�`�;�ٿ�j�#���@�KI*��3@4̐!?5}���B�@�� E�ٿ�!��
O�@���n�3@��S�!?W�^��)�@�� E�ٿ�!��
O�@���n�3@��S�!?W�^��)�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@	F��բٿzQ�����@������3@%�y�Ԑ!?d�v!Ο�@OQED�ٿ��V�*��@. �<��3@�b��!?�oLs�@OQED�ٿ��V�*��@. �<��3@�b��!?�oLs�@�?Q�ٿ���$L�@G�bP�3@ↄA��!?���K���@�?Q�ٿ���$L�@G�bP�3@ↄA��!?���K���@�t1ꥥٿ��' nX�@�v���3@d�`��!?T�L8��@�t1ꥥٿ��' nX�@�v���3@d�`��!?T�L8��@���9�ٿĩ��|�@���%@�3@FY�a�!?�tJ ��@���{�ٿP����T�@�O�zN�3@'o9�s�!?�4��+�@3�.���ٿ��(Y(��@��!x�3@�u�#��!?Q�$�|��@3�.���ٿ��(Y(��@��!x�3@�u�#��!?Q�$�|��@3�.���ٿ��(Y(��@��!x�3@�u�#��!?Q�$�|��@3�M]աٿO�2���@_o#t5�3@S~Dv�!?R�[l�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@EpW	�ٿq�P��e�@���C��3@��|�!?h��<�d�@@����ٿ��Q��"�@��Ũ��3@QJ@Ɛ!?n~߃�@@����ٿ��Q��"�@��Ũ��3@QJ@Ɛ!?n~߃�@(�R�ٿ��xw�@s�ݬ2�3@���$�!?4.w=�@(�R�ٿ��xw�@s�ݬ2�3@���$�!?4.w=�@(�R�ٿ��xw�@s�ݬ2�3@���$�!?4.w=�@(�R�ٿ��xw�@s�ݬ2�3@���$�!?4.w=�@�AҺ͟ٿ�;���B�@�l����3@>Y��ݐ!?�r4aQ�@�AҺ͟ٿ�;���B�@�l����3@>Y��ݐ!?�r4aQ�@��X�ٿ��4jE��@\�g�J�3@9��\Ր!?�Wm�0�@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@���ٿ��w��@�& ��3@�IA榐!?�۷���@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@ʻ�0�ٿ:K�b�@?~W���3@��}��!?z��!M�@&��2:�ٿ@�w]��@	>�5��3@1p7^r�!?�2l��P�@&��2:�ٿ@�w]��@	>�5��3@1p7^r�!?�2l��P�@&��2:�ٿ@�w]��@	>�5��3@1p7^r�!?�2l��P�@&��2:�ٿ@�w]��@	>�5��3@1p7^r�!?�2l��P�@��]?�ٿ�ux�4�@֜�W��3@`�7k�!?,���uF�@��]?�ٿ�ux�4�@֜�W��3@`�7k�!?,���uF�@��]?�ٿ�ux�4�@֜�W��3@`�7k�!?,���uF�@$��G�ٿO(i��@x�i@��3@��Љ�!?��ƫ_�@$��G�ٿO(i��@x�i@��3@��Љ�!?��ƫ_�@$��G�ٿO(i��@x�i@��3@��Љ�!?��ƫ_�@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@V(.��ٿ��'�@	%݉X�3@�; �!?�Ϻ���@��1В�ٿv��	�;�@��V�3@��w��!?�o�c���@��1В�ٿv��	�;�@��V�3@��w��!?�o�c���@��1В�ٿv��	�;�@��V�3@��w��!?�o�c���@��1В�ٿv��	�;�@��V�3@��w��!?�o�c���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@�����ٿe����@A
l�C�3@�F
�!?�ĖC���@䒺E��ٿ�:�WP;�@���(�3@=�pd��!?�����@!t$��ٿ(i�D���@?�SF�3@�mo��!?&�_��a�@X��u�ٿ���ȇ�@�;y|��3@Z��oܐ!?��,|l�@X��u�ٿ���ȇ�@�;y|��3@Z��oܐ!?��,|l�@X��u�ٿ���ȇ�@�;y|��3@Z��oܐ!?��,|l�@z�]�ٿ|�E&��@@?��3@�5�n�!?P�>�U��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@�̲mY�ٿ*�@LSZ�@\%��3@���y�!?<�*RQ��@����+�ٿ}�c��@o0ph��3@l�P��!?���[��@���V�ٿ�/L�e�@��z�3@����!?�P��ܰ�@x�>���ٿ���ʎ�@��N�{�3@w����!?!�Ot��@�����ٿA&���@�-u��3@���!?����]��@�����ٿA&���@�-u��3@���!?����]��@Gtjу�ٿ���o�@հO�w�3@C�x��!?������@Gtjу�ٿ���o�@հO�w�3@C�x��!?������@Gtjу�ٿ���o�@հO�w�3@C�x��!?������@"FlK|�ٿ�ّ�f�@��yX��3@��~�!?��-'��@"FlK|�ٿ�ّ�f�@��yX��3@��~�!?��-'��@qB:�ʜٿ�ئ	:�@ �uP��3@��&�!?B��|��@qB:�ʜٿ�ئ	:�@ �uP��3@��&�!?B��|��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�^���ٿ��]Y�@bބ���3@�[����!?��Ñ+��@�S�Y��ٿw������@���3@��U3��!?�q͓��@�S�Y��ٿw������@���3@��U3��!?�q͓��@�P|ףٿ���5:�@�I&��3@�^F��!?�ϻ�*��@]OF��ٿ�Ȱ����@������3@���"ѐ!?��Kvc�@(Ң(�ٿ_쫾���@�0G�^�3@$X����!?��K�@(Ң(�ٿ_쫾���@�0G�^�3@$X����!?��K�@(Ң(�ٿ_쫾���@�0G�^�3@$X����!?��K�@(Ң(�ٿ_쫾���@�0G�^�3@$X����!?��K�@(Ң(�ٿ_쫾���@�0G�^�3@$X����!?��K�@��C�ۧٿ����}�@�2����3@y��y�!?B��M���@��C�ۧٿ����}�@�2����3@y��y�!?B��M���@xI���ٿu�l:/��@T�+��3@,go�Q�!?ȓ����@���z�ٿi|ˤs�@8�����3@�vf�!?:��@�ٿd������@����H�3@�I�2��!?] \�O�@�ٿd������@����H�3@�I�2��!?] \�O�@T�o���ٿ�������@+Y&���3@�wxא!?����@-���@�ٿ��<���@�/�Rj�3@!^����!?�����@-���@�ٿ��<���@�/�Rj�3@!^����!?�����@-���@�ٿ��<���@�/�Rj�3@!^����!?�����@-���@�ٿ��<���@�/�Rj�3@!^����!?�����@-���@�ٿ��<���@�/�Rj�3@!^����!?�����@V+ZK|�ٿ�Y�����@��T��3@�\7��!?ڄY�i�@V+ZK|�ٿ�Y�����@��T��3@�\7��!?ڄY�i�@V+ZK|�ٿ�Y�����@��T��3@�\7��!?ڄY�i�@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@�~Iԡٿ�M![,�@P�ofZ�3@I���!?��+#���@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@��V7�ٿj����@@���;�3@��*��!?/���h�@�]٦ٿ�z2x�9�@�ܹ[N�3@Z��B��!?F`��6�@�b��}�ٿ��ڣ0�@������3@x��e2�!?O)%H���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�����ٿ���JG��@���3@�eY�!?M��*���@�Z]o�ٿ�Zoh9�@���rs�3@P��!?�$v@2��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@/dJ	v�ٿ��sO��@���l�3@��Iǐ!?�e[A��@�j����ٿ���T,r�@�L$j8�3@�K����!?�n{5q9�@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@tN����ٿ�f۰y5�@�}����3@(v���!?�`y��@Y���S�ٿ�����@2���3@�;[8Ԑ!?������@Y���S�ٿ�����@2���3@�;[8Ԑ!?������@Y���S�ٿ�����@2���3@�;[8Ԑ!?������@Y���S�ٿ�����@2���3@�;[8Ԑ!?������@qѳ��ٿ�8�x+�@�w_�V�3@uL�M�!?EP�ew�@qѳ��ٿ�8�x+�@�w_�V�3@uL�M�!?EP�ew�@qѳ��ٿ�8�x+�@�w_�V�3@uL�M�!?EP�ew�@qѳ��ٿ�8�x+�@�w_�V�3@uL�M�!?EP�ew�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@�o]0�ٿ�W,:��@/lW���3@��:ِ!?K%y�~l�@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@Q!���ٿ�r��,;�@�}j��3@2�����!?J�����@C���L�ٿ� #��@�X�>�3@E��j�!?����A��@C���L�ٿ� #��@�X�>�3@E��j�!?����A��@C���L�ٿ� #��@�X�>�3@E��j�!?����A��@n�cҡٿB���R�@۸�3�3@$�)��!?��)\_�@n�cҡٿB���R�@۸�3�3@$�)��!?��)\_�@LV_���ٿ��=����@��P�3@�g͐!?��BoXC�@LV_���ٿ��=����@��P�3@�g͐!?��BoXC�@LV_���ٿ��=����@��P�3@�g͐!?��BoXC�@LV_���ٿ��=����@��P�3@�g͐!?��BoXC�@LV_���ٿ��=����@��P�3@�g͐!?��BoXC�@����ٿ�驶���@ǩ��w�3@�y�͐!?���C�@����ٿ�驶���@ǩ��w�3@�y�͐!?���C�@s����ٿ��_���@+V�3@$Bj>��!?2�-;#�@s����ٿ��_���@+V�3@$Bj>��!?2�-;#�@Y7)�ٿFS3��@�׆|%�3@*3�g��!?u�bpG��@n��'h�ٿv�m���@�]�ߵ�3@T)-�ؐ!?U���)�@Z���ٿC��?
�@ȝG�o�3@餡�!?P&xk��@Z���ٿC��?
�@ȝG�o�3@餡�!?P&xk��@Z���ٿC��?
�@ȝG�o�3@餡�!?P&xk��@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�ð�k�ٿ����o\�@�%8���3@���_��!?��/�@�.�IL�ٿ�!����@�0�RT�3@K4솢�!?��[(�@�.�IL�ٿ�!����@�0�RT�3@K4솢�!?��[(�@�.�IL�ٿ�!����@�0�RT�3@K4솢�!?��[(�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@�2n��ٿ��b ��@�cs�3@�U�4��!?l��p�@Mb&-�ٿ�^ٳsW�@�Y?���3@ yH͐!?.r~�h�@Mb&-�ٿ�^ٳsW�@�Y?���3@ yH͐!?.r~�h�@Mb&-�ٿ�^ٳsW�@�Y?���3@ yH͐!?.r~�h�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�~/�ٿ!fX��@޻e(�3@>�d2��!?{���%�@�܌W�ٿ�yzΨ�@�R�'�3@����!?Q�H԰��@�����ٿ%s,��]�@�ޭ6'�3@Y���ǐ!?��f$���@�����ٿ%s,��]�@�ޭ6'�3@Y���ǐ!?��f$���@�����ٿ%s,��]�@�ޭ6'�3@Y���ǐ!?��f$���@� 2��ٿ*ch��x�@e�c���3@�g�l��!?�'��\��@� 2��ٿ*ch��x�@e�c���3@�g�l��!?�'��\��@-�-�ٿ����Q�@�����3@��b>��!?����@-�-�ٿ����Q�@�����3@��b>��!?����@-�-�ٿ����Q�@�����3@��b>��!?����@-�-�ٿ����Q�@�����3@��b>��!?����@awR(%�ٿf~�m!��@~ہ�V�3@N��V��!?���g�@awR(%�ٿf~�m!��@~ہ�V�3@N��V��!?���g�@H��ol�ٿݱ�6���@X3b�}�3@B$wj�!?���S��@cX�.��ٿ�sm���@:�±��3@�=����!?��"QWb�@cX�.��ٿ�sm���@:�±��3@�=����!?��"QWb�@cX�.��ٿ�sm���@:�±��3@�=����!?��"QWb�@cX�.��ٿ�sm���@:�±��3@�=����!?��"QWb�@�?f�تٿ/�ż���@�,�h�3@���T�!?1�zO���@�?f�تٿ/�ż���@�,�h�3@���T�!?1�zO���@#)Ҟ��ٿ��ұN�@��3@�w��N�!?8��C���@�_Q��ٿ=8���l�@l\����3@�G&�!?8���S�@�_Q��ٿ=8���l�@l\����3@�G&�!?8���S�@�_Q��ٿ=8���l�@l\����3@�G&�!?8���S�@�� k�ٿ���+�@�^�b��3@8��"�!?����h��@���iv�ٿ��8C���@������3@��'���!?��}�4�@���P�ٿ��W	���@�1��3@�
?F�!?�����@���P�ٿ��W	���@�1��3@�
?F�!?�����@���P�ٿ��W	���@�1��3@�
?F�!?�����@���P�ٿ��W	���@�1��3@�
?F�!?�����@��J�ٿ;$/��`�@�=}�j�3@�"�P�!?��ٚ-$�@��J�ٿ;$/��`�@�=}�j�3@�"�P�!?��ٚ-$�@��J�ٿ;$/��`�@�=}�j�3@�"�P�!?��ٚ-$�@��J�ٿ;$/��`�@�=}�j�3@�"�P�!?��ٚ-$�@��J�ٿ;$/��`�@�=}�j�3@�"�P�!?��ٚ-$�@q�*��ٿ�0�Xt��@d�^R�3@� ۰��!?e�%���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@�����ٿ�-X�D(�@�{�%�3@��{ߐ!?�
�i���@���ٿ)��O�@���$(�3@,�p\a�!?��E��@���ٿ)��O�@���$(�3@,�p\a�!?��E��@��qc�ٿ�=�!��@��)�3@8B���!?s��<��@��qc�ٿ�=�!��@��)�3@8B���!?s��<��@�p�ON�ٿg�Key�@NӥZ��3@�;��!?��Đm��@�p�ON�ٿg�Key�@NӥZ��3@�;��!?��Đm��@�p�ON�ٿg�Key�@NӥZ��3@�;��!?��Đm��@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@��!�,�ٿ�	��e��@�P����3@�,k���!?y����~�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@QK���ٿ�j[d���@�|U�I�3@�GG*ʐ!?~����,�@$�6�o�ٿ��ʼ���@	�����3@����!?[cv�*�@$�6�o�ٿ��ʼ���@	�����3@����!?[cv�*�@,Ġ� �ٿ,��� v�@:��L�3@�L[K͐!?d! <K��@,Ġ� �ٿ,��� v�@:��L�3@�L[K͐!?d! <K��@,Ġ� �ٿ,��� v�@:��L�3@�L[K͐!?d! <K��@n:�,{�ٿ�{:B���@XH�g��3@��ݐ!?;���@'��"��ٿ�C��,o�@լ".��3@H%��!?���0�@�^:��ٿܭ��c�@B<��3@$Sן�!?�'�~���@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@uI^�ٿ|��7���@���Ķ�3@��	mސ!?�U���f�@z�*U�ٿm���ZF�@z���3@y,�
'�!?1)���@M�V¡ٿ_1p�@�r�t4�3@��6G��!?#��u@W�@M�V¡ٿ_1p�@�r�t4�3@��6G��!?#��u@W�@M�V¡ٿ_1p�@�r�t4�3@��6G��!?#��u@W�@%�]�d�ٿ��X�K�@��և��3@>ϫ��!?U!�&��@%�]�d�ٿ��X�K�@��և��3@>ϫ��!?U!�&��@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@#���ٿ�V��@q�3�[�3@�5���!?Y�B�D�@k���e�ٿM�&�@�ʣg��3@m�n<�!?}��L�@k���e�ٿM�&�@�ʣg��3@m�n<�!?}��L�@k���e�ٿM�&�@�ʣg��3@m�n<�!?}��L�@k���e�ٿM�&�@�ʣg��3@m�n<�!?}��L�@ov�s'�ٿ{z�S�`�@�B��3@�F1�,�!?~*�7~�@ܵ��ӟٿ,�:]5�@��T�3@:�ue	�!?�#�=¥�@ܵ��ӟٿ,�:]5�@��T�3@:�ue	�!?�#�=¥�@ܵ��ӟٿ,�:]5�@��T�3@:�ue	�!?�#�=¥�@ܵ��ӟٿ,�:]5�@��T�3@:�ue	�!?�#�=¥�@ܵ��ӟٿ,�:]5�@��T�3@:�ue	�!?�#�=¥�@J�}�ٿ9�D*��@��x�3@��Č�!?�:�=��@�[#]��ٿ�X\C�N�@�m�>��3@x���!?��p�@�[#]��ٿ�X\C�N�@�m�>��3@x���!?��p�@�'9ޡٿ ���@^HOs�3@U��ː!?'{�=��@�'9ޡٿ ���@^HOs�3@U��ː!?'{�=��@�'9ޡٿ ���@^HOs�3@U��ː!?'{�=��@�'9ޡٿ ���@^HOs�3@U��ː!?'{�=��@�'9ޡٿ ���@^HOs�3@U��ː!?'{�=��@�zL
�ٿ_o�����@���.K�3@4�ů�!?{>p���@�zL
�ٿ_o�����@���.K�3@4�ů�!?{>p���@�zL
�ٿ_o�����@���.K�3@4�ů�!?{>p���@�zL
�ٿ_o�����@���.K�3@4�ů�!?{>p���@
(�m�ٿ���KU�@��ѫ�3@ymW,p�!?�IT{�X�@
(�m�ٿ���KU�@��ѫ�3@ymW,p�!?�IT{�X�@
(�m�ٿ���KU�@��ѫ�3@ymW,p�!?�IT{�X�@[�t��ٿ|��Ym��@��=��3@p�n�Ő!?:�I8G��@[�t��ٿ|��Ym��@��=��3@p�n�Ő!?:�I8G��@l�V�ƥٿOU�6��@mk���3@z{�f��!?`�e��@c�1���ٿ ��A��@���h��3@-!iy�!?gk�����@c�1���ٿ ��A��@���h��3@-!iy�!?gk�����@c�1���ٿ ��A��@���h��3@-!iy�!?gk�����@�F�!�ٿ���c9�@��	]�3@U��篐!?����~�@�F�!�ٿ���c9�@��	]�3@U��篐!?����~�@qq�F�ٿ���%1�@B��eG�3@�,����!?��ǌ��@g�����ٿ �`����@G.�J��3@�s��!?��њ�)�@5'p���ٿj?¼���@!|J(�3@@� U��!?�����G�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@�U���ٿ�x�5?�@�����3@[6�ِ!?�x;��#�@:��	ȟٿfv�f�3�@���w��3@"N�R�!?�ķ`���@:��	ȟٿfv�f�3�@���w��3@"N�R�!?�ķ`���@:��	ȟٿfv�f�3�@���w��3@"N�R�!?�ķ`���@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�$~�W�ٿ a��?r�@��:o�3@t�8ΐ!?�	��~�@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@�����ٿ�Ni�_�@��1�3@^��x�!?vy�DO��@���is�ٿ��xf8l�@l$�8��3@�~Z�z�!?�����|�@���is�ٿ��xf8l�@l$�8��3@�~Z�z�!?�����|�@���is�ٿ��xf8l�@l$�8��3@�~Z�z�!?�����|�@�o��ٿ��h�D �@~
��3@�$��^�!?s�Ę�;�@�o��ٿ��h�D �@~
��3@�$��^�!?s�Ę�;�@�d���ٿ�W��@�2֡��3@ι�i��!?�]K�K��@�d���ٿ�W��@�2֡��3@ι�i��!?�]K�K��@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@�0�!�ٿ�[�G��@��Ϝ{�3@��-攐!?/���J]�@����ٿ���M�@����3@�D(	|�!?����(g�@������ٿ��W�J�@���E�3@s~�j��!?���+�2�@������ٿ��W�J�@���E�3@s~�j��!?���+�2�@������ٿ��W�J�@���E�3@s~�j��!?���+�2�@\�nˤٿzr�gH�@���3@<"(��!?��ӝ�@\�nˤٿzr�gH�@���3@<"(��!?��ӝ�@\�nˤٿzr�gH�@���3@<"(��!?��ӝ�@\�nˤٿzr�gH�@���3@<"(��!?��ӝ�@�Tk�ٿB������@gm����3@��ۺĐ!?�W,�=�@�Tk�ٿB������@gm����3@��ۺĐ!?�W,�=�@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@�pt��ٿ�CBm"�@7�M��3@����!?ɬ�O���@l<�ln�ٿ㝎As��@%�Be�3@U�a��!?D��m��@l<�ln�ٿ㝎As��@%�Be�3@U�a��!?D��m��@Q.wBP�ٿE0:e�`�@4EF��3@K�x��!?p�/���@Q.wBP�ٿE0:e�`�@4EF��3@K�x��!?p�/���@!�$,��ٿ����U%�@�(\�3@���v��!??����*�@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@���ҡٿ�k��Ȯ�@-P=�,�3@�E�]��!?7�����@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@T���g�ٿL	T�`Z�@#5� ��3@.2d���!?��ݸ��@��u���ٿ����ٮ�@`q�a.�3@���+�!?�żt�S�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�dK���ٿ�?�+���@B O�7�3@�/��!?��1��,�@�XsШٿ�����@��e���3@`��)�!?-Ζ{c��@�XsШٿ�����@��e���3@`��)�!?-Ζ{c��@�XsШٿ�����@��e���3@`��)�!?-Ζ{c��@�XsШٿ�����@��e���3@`��)�!?-Ζ{c��@�XsШٿ�����@��e���3@`��)�!?-Ζ{c��@�˟4�ٿ)�$N�"�@�8�̎�3@�����!?r�wp�@�)��=�ٿ\���F��@9����3@��Ґ!?y���s��@�)��=�ٿ\���F��@9����3@��Ґ!?y���s��@�)��=�ٿ\���F��@9����3@��Ґ!?y���s��@�)��=�ٿ\���F��@9����3@��Ґ!?y���s��@rz�Šٿt����@�0�x��3@:�9\��!?Ns��@���z�ٿ�v��@b��>��3@������!?*��^��@���z�ٿ�v��@b��>��3@������!?*��^��@���z�ٿ�v��@b��>��3@������!?*��^��@���z�ٿ�v��@b��>��3@������!?*��^��@��x=�ٿ|^<T˝�@	�{���3@rF��p�!?1q�V��@��x=�ٿ|^<T˝�@	�{���3@rF��p�!?1q�V��@��x=�ٿ|^<T˝�@	�{���3@rF��p�!?1q�V��@��x=�ٿ|^<T˝�@	�{���3@rF��p�!?1q�V��@G��&�ٿ� �<ɔ�@�9�Al�3@��=��!?�,a��@G��&�ٿ� �<ɔ�@�9�Al�3@��=��!?�,a��@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@����ٿ�3�^���@"S���3@�+*���!? 3�2���@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@3�Q��ٿ"p;���@]H4<�3@~��t��!?:�Mr��@5s��\�ٿ����0|�@���i�3@�H���!?U������@5s��\�ٿ����0|�@���i�3@�H���!?U������@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@&�d�ٿ���Z��@TI`?T�3@��׿Đ!?��/o���@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@�s�t�ٿ����@���O�3@ƲxGԐ!?,֩�p��@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@��n�ٿ6V%��1�@����3@ �fې!?�э҈X�@�����ٿs�0�;�@ͣ(��3@z_�4��!?�)�rV��@�����ٿs�0�;�@ͣ(��3@z_�4��!?�)�rV��@�����ٿs�0�;�@ͣ(��3@z_�4��!?�)�rV��@؋ŊD�ٿ �����@f��fV�3@_�� ��!?Z�֠'�@؋ŊD�ٿ �����@f��fV�3@_�� ��!?Z�֠'�@؋ŊD�ٿ �����@f��fV�3@_�� ��!?Z�֠'�@����ٿI��$u�@�n��l�3@�����!?8A�����@����ٿI��$u�@�n��l�3@�����!?8A�����@�d�]��ٿv�����@�����3@�r��!?��g�+�@	�S�ٿ^]�`�?�@+�&@�3@���0�!?�ӹ=�Z�@	�S�ٿ^]�`�?�@+�&@�3@���0�!?�ӹ=�Z�@	�S�ٿ^]�`�?�@+�&@�3@���0�!?�ӹ=�Z�@	�S�ٿ^]�`�?�@+�&@�3@���0�!?�ӹ=�Z�@�'��	�ٿY���t�@�d��3@F�"��!?fc���@�'��	�ٿY���t�@�d��3@F�"��!?fc���@�'��	�ٿY���t�@�d��3@F�"��!?fc���@2��9�ٿtE@&<�@^��3@0햘�!?��q���@2��9�ٿtE@&<�@^��3@0햘�!?��q���@2��9�ٿtE@&<�@^��3@0햘�!?��q���@�.*��ٿ&h��.��@�L�t�3@�Y���!?���2��@�.*��ٿ&h��.��@�L�t�3@�Y���!?���2��@�.*��ٿ&h��.��@�L�t�3@�Y���!?���2��@���V�ٿՅ����@�EW�3@"�7Ő!?D�@}��@���V�ٿՅ����@�EW�3@"�7Ő!?D�@}��@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@ݔ:Рٿ�R3�m�@�Kɘ��3@�u�	��!?��07bb�@���|�ٿޢ�^���@^]�=��3@��d�!?��g���@���|�ٿޢ�^���@^]�=��3@��d�!?��g���@�2�X#�ٿ��To��@��-i�3@�:�K��!?�~￁��@zrmW~�ٿI�����@�f�Z�3@���9��!?������@�l�s�ٿ*�W�7r�@ k���3@`���e�!?#��5U��@�l�s�ٿ*�W�7r�@ k���3@`���e�!?#��5U��@�l�s�ٿ*�W�7r�@ k���3@`���e�!?#��5U��@�l�s�ٿ*�W�7r�@ k���3@`���e�!?#��5U��@�j��ٿ�eۯ��@�^댠�3@�a�PU�!?<u�a��@�j��ٿ�eۯ��@�^댠�3@�a�PU�!?<u�a��@�j��ٿ�eۯ��@�^댠�3@�a�PU�!?<u�a��@�j��ٿ�eۯ��@�^댠�3@�a�PU�!?<u�a��@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@'%Nq�ٿa1���>�@���q��3@�@%�P�!?���9���@�)Vl�ٿ�`����@�3'��3@�]n���!?-��9�@�)Vl�ٿ�`����@�3'��3@�]n���!?-��9�@�)Vl�ٿ�`����@�3'��3@�]n���!?-��9�@�)Vl�ٿ�`����@�3'��3@�]n���!?-��9�@�)Vl�ٿ�`����@�3'��3@�]n���!?-��9�@��nDĦٿ�5��7�@����3@��6���!?��r,nT�@+��)�ٿrt��@{.O���3@���[v�!?��|{���@�mA��ٿx�R����@j�+�R�3@=7���!?��ӋuQ�@�mA��ٿx�R����@j�+�R�3@=7���!?��ӋuQ�@I�E
�ٿx1�����@A��s��3@z��WА!?�$�QK�@O��ٿM���T�@�[���3@�GC�G�!?9��>���@O��ٿM���T�@�[���3@�GC�G�!?9��>���@BF�ٿP�f�@K?Mg�3@(?��y�!?u=�
���@_��b.�ٿ��f�@OxZ�`�3@�(�q��!?�[g|�_�@_��b.�ٿ��f�@OxZ�`�3@�(�q��!?�[g|�_�@_��b.�ٿ��f�@OxZ�`�3@�(�q��!?�[g|�_�@_��b.�ٿ��f�@OxZ�`�3@�(�q��!?�[g|�_�@� ��2�ٿ{�k���@���(�3@��2�f�!?��z�1��@� ��2�ٿ{�k���@���(�3@��2�f�!?��z�1��@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@SC1!��ٿ�w��x�@����3@p�N�֐!?$���on�@Ѓ��n�ٿ���@�@KߪG�3@*�Ώ��!?~u4���@Ѓ��n�ٿ���@�@KߪG�3@*�Ώ��!?~u4���@Ѓ��n�ٿ���@�@KߪG�3@*�Ώ��!?~u4���@Ѓ��n�ٿ���@�@KߪG�3@*�Ώ��!?~u4���@8��ʟٿ��)��@��M$�3@���g�!?�t(W�a�@��1��ٿ��KVi�@��%��3@XV2�ϐ!?B��n���@��1��ٿ��KVi�@��%��3@XV2�ϐ!?B��n���@�V��'�ٿ���m�
�@:7���3@��]��!?&q~�7�@0o�M۞ٿ!с���@?.���3@y5ؙ�!? ׶�.�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@�m�J�ٿɿY2%�@��bq
�3@���Ӣ�!?��c�#�@>�{O�ٿ�<D"��@�E���3@6'�Ő!?������@�M����ٿ�iL@�@.�D�-�3@�*�(א!?�l��@�M����ٿ�iL@�@.�D�-�3@�*�(א!?�l��@�M����ٿ�iL@�@.�D�-�3@�*�(א!?�l��@�M����ٿ�iL@�@.�D�-�3@�*�(א!?�l��@��zF��ٿ�/����@��3=�3@I<w7��!?���N��@��zF��ٿ�/����@��3=�3@I<w7��!?���N��@��zF��ٿ�/����@��3=�3@I<w7��!?���N��@��zF��ٿ�/����@��3=�3@I<w7��!?���N��@��zF��ٿ�/����@��3=�3@I<w7��!?���N��@_Ҋ��ٿq�$�@��)��3@٘^��!?�҂��@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@;�퍞ٿK�.i��@��)���3@��!���!?j�lgQ�@�v���ٿ�l�����@c1�E�3@�0�+ �!?��B�|�@�v���ٿ�l�����@c1�E�3@�0�+ �!?��B�|�@�v���ٿ�l�����@c1�E�3@�0�+ �!?��B�|�@�v���ٿ�l�����@c1�E�3@�0�+ �!?��B�|�@��2�ٿ����"�@�"F�3@����ߐ!?����r�@�aV�ٿ�������@O��z�3@�j>�ݐ!?�-tr��@�U��ٿ������@����J�3@6��2ߐ!?cZ;���@�U��ٿ������@����J�3@6��2ߐ!?cZ;���@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@gg���ٿw�/3���@+���3@�EFD��!?��
�@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@�Bh�=�ٿo����@o"b�f�3@);Ɛ!?f�ߘp��@#�H���ٿ�c�W�@�:4��3@9��Oؐ!?�W�ǃ�@+[
��ٿ 6�
zI�@��@n�3@Ա[�͐!?�����@+[
��ٿ 6�
zI�@��@n�3@Ա[�͐!?�����@+[
��ٿ 6�
zI�@��@n�3@Ա[�͐!?�����@+[
��ٿ 6�
zI�@��@n�3@Ա[�͐!?�����@+[
��ٿ 6�
zI�@��@n�3@Ա[�͐!?�����@45��ٿ�8�tB�@�;r	��3@��ǳ��!?c���%�@��jg��ٿ��8���@)����3@;��;��!?�j���@��jg��ٿ��8���@)����3@;��;��!?�j���@��jg��ٿ��8���@)����3@;��;��!?�j���@��jg��ٿ��8���@)����3@;��;��!?�j���@��a�k�ٿ#��"	�@�k���3@���,��!?7s��kF�@��a�k�ٿ#��"	�@�k���3@���,��!?7s��kF�@��a�k�ٿ#��"	�@�k���3@���,��!?7s��kF�@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@'G����ٿ�J0�e�@�0��	�3@�G�ꡐ!?��^c��@IK(�ٿr��c���@�O3�I�3@�[�Ԡ�!?���A��@IK(�ٿr��c���@�O3�I�3@�[�Ԡ�!?���A��@��qw[�ٿ��!ĉ�@+��U�3@l_M7��!?N�*!C0�@��r$��ٿ-%_���@�?ĝ��3@%�J!?�����@Ձ�L��ٿ������@�����3@Bh � �!?��Xݿ�@a/*�ٿ·��@�n>�<�3@���!?�s/T���@a/*�ٿ·��@�n>�<�3@���!?�s/T���@�j��.�ٿ�h ��`�@��b��3@૧�>�!?��dRa�@BrٿG�µ��@B����3@�l�T�!?�.f"�@BrٿG�µ��@B����3@�l�T�!?�.f"�@BrٿG�µ��@B����3@�l�T�!?�.f"�@BrٿG�µ��@B����3@�l�T�!?�.f"�@BrٿG�µ��@B����3@�l�T�!?�.f"�@�)ԊP�ٿˠ˵��@�l2$\�3@D&�ސ!?{_ү�@�)ԊP�ٿˠ˵��@�l2$\�3@D&�ސ!?{_ү�@�)ԊP�ٿˠ˵��@�l2$\�3@D&�ސ!?{_ү�@�i��ٿus�0�m�@������3@�e�ߐ!?t&����@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@���a�ٿ$ډd�@R2���3@��wd�!?��%Y���@z�{��ٿf/�U�o�@�{6�Y�3@�Q�^�!?�_4/��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@����ٿ�?�:4x�@!ns��3@�Dl�a�!?���d��@$����ٿ�mZ}�@2�����3@�H~�c�!?������@$����ٿ�mZ}�@2�����3@�H~�c�!?������@$����ٿ�mZ}�@2�����3@�H~�c�!?������@8���u�ٿ�~�x���@I� ��3@��ː!?�4�t�@8���u�ٿ�~�x���@I� ��3@��ː!?�4�t�@��(�ߚٿ�)�Sj�@�추�3@����2�!?$��q���@VqB�ٿ��Q���@θ�=��3@Mz��͐!?C���C��@�p}B�ٿ�7��y5�@c:���3@:ժ�!?��aU��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@�,s�ٿ)�O�@ͺR3��3@O��6�!?xέ$z��@'�,��ٿ�~����@v�o���3@�8�Ő!?>�5��a�@'�,��ٿ�~����@v�o���3@�8�Ő!?>�5��a�@'�,��ٿ�~����@v�o���3@�8�Ő!?>�5��a�@'�,��ٿ�~����@v�o���3@�8�Ő!?>�5��a�@'�,��ٿ�~����@v�o���3@�8�Ő!?>�5��a�@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@������ٿRq���)�@�g��g�3@�L�H��!?���e���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@E���ٿ�E�H�@�b>��3@��7���!?P�k���@�J��ٿ����Qr�@��%�V�3@GFx��!?bD���@E?t���ٿ��S����@�	��3@�9(ю�!?u����@E?t���ٿ��S����@�	��3@�9(ю�!?u����@E?t���ٿ��S����@�	��3@�9(ю�!?u����@E?t���ٿ��S����@�	��3@�9(ю�!?u����@h�'ٿ��߸��@��z���3@<�� ��!?�F��b&�@h�'ٿ��߸��@��z���3@<�� ��!?�F��b&�@h�'ٿ��߸��@��z���3@<�� ��!?�F��b&�@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@Nq�%Ɲٿ��/g��@-��+�3@�A!Ԑ!?w��֮��@w�Ro��ٿ���CN��@��S:�3@XW���!?�QP�V�@bpjh�ٿa8�ķ��@�N��z�3@/*���!?�E�z�^�@bpjh�ٿa8�ķ��@�N��z�3@/*���!?�E�z�^�@bpjh�ٿa8�ķ��@�N��z�3@/*���!?�E�z�^�@酒�@�ٿ�������@,H���3@�� �5�!?F�YJc��@��4|�ٿ���9ھ�@�sJ��3@���#�!?=O�#I�@��4|�ٿ���9ھ�@�sJ��3@���#�!?=O�#I�@��4|�ٿ���9ھ�@�sJ��3@���#�!?=O�#I�@��4|�ٿ���9ھ�@�sJ��3@���#�!?=O�#I�@��X�U�ٿ���d��@4�ݧ�3@�q�f�!?(��6��@rH�	�ٿ>�R,44�@	ᡙ��3@�俐!?e�=��@h,�y��ٿ�� l���@7�6�8�3@�=`ʮ�!?�1�)���@h,�y��ٿ�� l���@7�6�8�3@�=`ʮ�!?�1�)���@h,�y��ٿ�� l���@7�6�8�3@�=`ʮ�!?�1�)���@h,�y��ٿ�� l���@7�6�8�3@�=`ʮ�!?�1�)���@�ھϖ�ٿ,��t��@2f؋�3@)�3�ǐ!?&��2)��@�ھϖ�ٿ,��t��@2f؋�3@)�3�ǐ!?&��2)��@�ھϖ�ٿ,��t��@2f؋�3@)�3�ǐ!?&��2)��@�ھϖ�ٿ,��t��@2f؋�3@)�3�ǐ!?&��2)��@��ܡٿ�Zs5��@�j;8#�3@x!-@��!?J]�^��@��ܡٿ�Zs5��@�j;8#�3@x!-@��!?J]�^��@��ܡٿ�Zs5��@�j;8#�3@x!-@��!?J]�^��@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@h:�/�ٿ��_WG��@z��'��3@��o�!?�#�8R�@�����ٿO���u?�@}!����3@HE���!?����Ѻ�@�����ٿO���u?�@}!����3@HE���!?����Ѻ�@��R1l�ٿag���@����_�3@�{;O�!?��~���@��R1l�ٿag���@����_�3@�{;O�!?��~���@P����ٿGF��Q�@N�5ߍ�3@��E>�!?�į��@P����ٿGF��Q�@N�5ߍ�3@��E>�!?�į��@�+N���ٿ?�����@*�|T��3@�Μ���!?��e+���@.�c9��ٿ�ɡ+Z�@rGd%�3@�߿I�!?�v��Y�@.�c9��ٿ�ɡ+Z�@rGd%�3@�߿I�!?�v��Y�@.�c9��ٿ�ɡ+Z�@rGd%�3@�߿I�!?�v��Y�@.�c9��ٿ�ɡ+Z�@rGd%�3@�߿I�!?�v��Y�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�Ҙ�j�ٿ_*��@���J��3@��[��!?r�.��:�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�V[,��ٿ2��`[A�@�gG(m�3@[��&ѐ!?���w�@�><�ٿ
��'k�@x\Ba��3@PSm��!?�	6 �@(5�K֗ٿI[�(��@&��3@��L���!?��(���@(5�K֗ٿI[�(��@&��3@��L���!?��(���@(5�K֗ٿI[�(��@&��3@��L���!?��(���@�Q�W��ٿK�"�H��@��0?��3@vI����!?߳:�H9�@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@Q7>Ҟٿx'n���@*�v�3@2"N��!?�L=c��@��N���ٿ����V��@Bת>��3@�T޸��!?aY��@��N���ٿ����V��@Bת>��3@�T޸��!?aY��@��N���ٿ����V��@Bת>��3@�T޸��!?aY��@��N���ٿ����V��@Bת>��3@�T޸��!?aY��@��N���ٿ����V��@Bת>��3@�T޸��!?aY��@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@ZlT>�ٿG��`!�@���/��3@���!?�-����@�b���ٿk~t����@��x8��3@������!?qMKx��@�b���ٿk~t����@��x8��3@������!?qMKx��@�DN��ٿ�q�gs��@AJ٧��3@�]U�֐!?�I�����@�DN��ٿ�q�gs��@AJ٧��3@�]U�֐!?�I�����@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@�'�o�ٿ�K�۠��@���(��3@m��א!?��$�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@`.7(S�ٿc����@���x�3@c�_a	�!?T�"�2�@�U�7��ٿ3%g~��@�>H�3@�1���!?I�Uu�@�U�7��ٿ3%g~��@�>H�3@�1���!?I�Uu�@�U�7��ٿ3%g~��@�>H�3@�1���!?I�Uu�@�U�7��ٿ3%g~��@�>H�3@�1���!?I�Uu�@�᰼�ٿ�Y)݆�@�0�r=�3@?W-�ϐ!?i����@�᰼�ٿ�Y)݆�@�0�r=�3@?W-�ϐ!?i����@�᰼�ٿ�Y)݆�@�0�r=�3@?W-�ϐ!?i����@�᰼�ٿ�Y)݆�@�0�r=�3@?W-�ϐ!?i����@�����ٿ9���@5k�Z�3@�tѐ!?��%����@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@w�@�U�ٿM��\~�@�>L4��3@˳���!?� /?[��@��OX�ٿT���@xs���3@�v'^��!?���'�@��OX�ٿT���@xs���3@�v'^��!?���'�@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@Q{P��ٿ�w�a��@	����3@�WH|ߐ!?3�v���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@ۤie�ٿ�h{e���@q�驮�3@�?�ِ!?�Ҟ���@;!���ٿh4"c���@���Y��3@K��jې!?n�T�t��@���t�ٿ7���I^�@��[�y�3@�o�^�!?�j��@���t�ٿ7���I^�@��[�y�3@�o�^�!?�j��@��xD��ٿ�VL�R�@��B+��3@�v���!?�q��F��@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@!_�ﴜٿQeQ0�t�@<\8�3@䫏o��!?��-���@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@R�\�ٿ�f>�s��@NԘ���3@r�P!��!?���x�<�@0�3N��ٿ(�Q�:�@י�R%�3@:�<§�!?��9j2�@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@E̢ٿ���B��@�(�B��3@��ԟ��!?��j��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@�`�b��ٿ@HZ�	��@&��V�3@OOq���!?�a��@���ݜٿe�^���@X�,���3@$#����!?7�v��@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@�܋��ٿ?e��P�@�����3@�{Q���!?������@Z�a��ٿ�L��hc�@4]�F��3@Kb7�!?�ۛ ֨�@Z�a��ٿ�L��hc�@4]�F��3@Kb7�!?�ۛ ֨�@Z�a��ٿ�L��hc�@4]�F��3@Kb7�!?�ۛ ֨�@�aM�M�ٿ@	2=��@�s��3@�/+�!?q��.=��@�aM�M�ٿ@	2=��@�s��3@�/+�!?q��.=��@�aM�M�ٿ@	2=��@�s��3@�/+�!?q��.=��@�aM�M�ٿ@	2=��@�s��3@�/+�!?q��.=��@�aM�M�ٿ@	2=��@�s��3@�/+�!?q��.=��@��ߚٿp��u&�@�Vd ��3@�K��!?238���@7tB^G�ٿ�=�O�*�@oG/y�3@�DՕ�!?T��$3�@�iXFӡٿJБ!iv�@P&�K��3@{3��!?��#����@�iXFӡٿJБ!iv�@P&�K��3@{3��!?��#����@^�ක�ٿH��{r��@?v���3@�:���!?(	�m���@^�ක�ٿH��{r��@?v���3@�:���!?(	�m���@�����ٿ��û��@
��j��3@Zݟ��!?�&�X�@�����ٿ��û��@
��j��3@Zݟ��!?�&�X�@7D�ٿ������@�]axf�3@4A�Ð!?�w�18�@7D�ٿ������@�]axf�3@4A�Ð!?�w�18�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@�T�!�ٿ����W�@�+QmH�3@��FŐ!?Rb�y�@[��~n�ٿ� ���@bF�Vo�3@k�N=��!?�s�m��@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@�e>=Z�ٿ�y�S��@M0�^�3@��|��!?�Ԯr�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Y�\N��ٿ��Kl ��@=����3@�cM��!?���"P�@Vn 86�ٿ^��G�u�@��F���3@K۾Z��!?VA�t��@Vn 86�ٿ^��G�u�@��F���3@K۾Z��!?VA�t��@����o�ٿD�Q�Â�@��
*>�3@T)5i��!?wP�'W�@����o�ٿD�Q�Â�@��
*>�3@T)5i��!?wP�'W�@����o�ٿD�Q�Â�@��
*>�3@T)5i��!?wP�'W�@����o�ٿD�Q�Â�@��
*>�3@T)5i��!?wP�'W�@�s�B.�ٿf����@7uVu��3@bg��Ő!?[�j���@�s�B.�ٿf����@7uVu��3@bg��Ő!?[�j���@��J��ٿ��VC�@�{g�3@׊�Yא!?��[��3�@��J��ٿ��VC�@�{g�3@׊�Yא!?��[��3�@��J��ٿ��VC�@�{g�3@׊�Yא!?��[��3�@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@_W�Z�ٿ���C�@=x����3@��"H̐!?<����@q��B9�ٿ%v*2t�@&C�<��3@��L�̐!?�q�t.�@q��B9�ٿ%v*2t�@&C�<��3@��L�̐!?�q�t.�@q��B9�ٿ%v*2t�@&C�<��3@��L�̐!?�q�t.�@�!�� �ٿ3�\�@/2�q�3@�<Đ!?�������@�!�� �ٿ3�\�@/2�q�3@�<Đ!?�������@�!�� �ٿ3�\�@/2�q�3@�<Đ!?�������@�!�� �ٿ3�\�@/2�q�3@�<Đ!?�������@�!�� �ٿ3�\�@/2�q�3@�<Đ!?�������@�D���ٿd�a���@�B�Q�3@��Ҩ��!?֮�oU��@�D���ٿd�a���@�B�Q�3@��Ҩ��!?֮�oU��@�D���ٿd�a���@�B�Q�3@��Ҩ��!?֮�oU��@�D���ٿd�a���@�B�Q�3@��Ҩ��!?֮�oU��@�D���ٿd�a���@�B�Q�3@��Ҩ��!?֮�oU��@4�>��ٿbGg/۽�@Λ ��3@��"�!?�<lZ��@4�>��ٿbGg/۽�@Λ ��3@��"�!?�<lZ��@m6���ٿw�#xφ�@������3@�紐!?J>{'є�@���C�ٿ0�4c��@n�J��3@�ɜ�ؐ!?v�27�@_5�i�ٿD�q�c�@QI��Y�3@�9���!?�/�T�@_5�i�ٿD�q�c�@QI��Y�3@�9���!?�/�T�@w����ٿ h[_�
�@��Z��3@m] �ɐ!?bN��v�@w����ٿ h[_�
�@��Z��3@m] �ɐ!?bN��v�@w����ٿ h[_�
�@��Z��3@m] �ɐ!?bN��v�@w����ٿ h[_�
�@��Z��3@m] �ɐ!?bN��v�@�M^���ٿ㳼�7u�@�C���3@?>gM��!?��X7=]�@����ٿ�{���t�@=�M"�3@6a�ݐ!?PF�@��@����ٿ�{���t�@=�M"�3@6a�ݐ!?PF�@��@����ٿ�{���t�@=�M"�3@6a�ݐ!?PF�@��@����ٿ�{���t�@=�M"�3@6a�ݐ!?PF�@��@����ٿ�{���t�@=�M"�3@6a�ݐ!?PF�@��@͵´	�ٿ�>y�WL�@O�?���3@�8�א!?�m�Q:�@͵´	�ٿ�>y�WL�@O�?���3@�8�א!?�m�Q:�@͵´	�ٿ�>y�WL�@O�?���3@�8�א!?�m�Q:�@͵´	�ٿ�>y�WL�@O�?���3@�8�א!?�m�Q:�@]c|-�ٿ�/@��@���{��3@c���ڐ!?�%��{�@]c|-�ٿ�/@��@���{��3@c���ڐ!?�%��{�@]c|-�ٿ�/@��@���{��3@c���ڐ!?�%��{�@]c|-�ٿ�/@��@���{��3@c���ڐ!?�%��{�@]c|-�ٿ�/@��@���{��3@c���ڐ!?�%��{�@0=�G��ٿ��a����@�ǳ��3@�����!?:�����@0=�G��ٿ��a����@�ǳ��3@�����!?:�����@&B�g�ٿ:{��0�@�/s���3@�%&�ѐ!?��'���@&B�g�ٿ:{��0�@�/s���3@�%&�ѐ!?��'���@&B�g�ٿ:{��0�@�/s���3@�%&�ѐ!?��'���@&B�g�ٿ:{��0�@�/s���3@�%&�ѐ!?��'���@&B�g�ٿ:{��0�@�/s���3@�%&�ѐ!?��'���@^�q�ٿ�?��H��@�xш�3@���a��!?� ,�+F�@^�q�ٿ�?��H��@�xш�3@���a��!?� ,�+F�@6���ڧٿwK���@��Vm�3@dB��ɐ!?���G8�@6���ڧٿwK���@��Vm�3@dB��ɐ!?���G8�@6���ڧٿwK���@��Vm�3@dB��ɐ!?���G8�@6���ڧٿwK���@��Vm�3@dB��ɐ!?���G8�@6���ڧٿwK���@��Vm�3@dB��ɐ!?���G8�@�����ٿ��*�Ft�@��$"/�3@�ⶉ$�!?¹P����@?�/�âٿ���]!6�@h񥙝�3@iC�A%�!?�I�8��@?�/�âٿ���]!6�@h񥙝�3@iC�A%�!?�I�8��@k㩨B�ٿ����8�@����3@����!?��u��#�@k㩨B�ٿ����8�@����3@����!?��u��#�@�*S��ٿe�^>�@��pZ��3@ׄ'`�!?�֓_f�@��5l;�ٿ=��7͓�@ua���3@�`5��!?���a���@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@۱.z�ٿ=x�=s�@Q T=��3@4yu��!?�S��/�@at\Ո�ٿJ��R��@.�$�N�3@�wu$��!?�In0��@at\Ո�ٿJ��R��@.�$�N�3@�wu$��!?�In0��@at\Ո�ٿJ��R��@.�$�N�3@�wu$��!?�In0��@at\Ո�ٿJ��R��@.�$�N�3@�wu$��!?�In0��@at\Ո�ٿJ��R��@.�$�N�3@�wu$��!?�In0��@ʨ�y��ٿ�;�Q��@����3@Ñ�%�!?w�y��@ʨ�y��ٿ�;�Q��@����3@Ñ�%�!?w�y��@ʨ�y��ٿ�;�Q��@����3@Ñ�%�!?w�y��@ʨ�y��ٿ�;�Q��@����3@Ñ�%�!?w�y��@{��`��ٿ��:�x��@�B<��3@�C�N�!?�~HN���@{��`��ٿ��:�x��@�B<��3@�C�N�!?�~HN���@{��`��ٿ��:�x��@�B<��3@�C�N�!?�~HN���@��u�ٿ����m�@��j�3@h�U�!?TEs{��@��u�ٿ����m�@��j�3@h�U�!?TEs{��@��u�ٿ����m�@��j�3@h�U�!?TEs{��@��u�ٿ����m�@��j�3@h�U�!?TEs{��@��u�ٿ����m�@��j�3@h�U�!?TEs{��@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@S�	А�ٿ>�OUT�@�7}L��3@gt_��!?�����@�9eg�ٿ-�8l}�@i{F	�3@�}�ؐ!?���WE�@���g�ٿ��+�o�@����Y�3@ߐ���!?��?��@���ٿlv$�s�@�x@D�3@�����!?�r��/��@�R�2Y�ٿ�`l�g�@"?7(5�3@r+�ΐ!?�������@�R�2Y�ٿ�`l�g�@"?7(5�3@r+�ΐ!?�������@�R�2Y�ٿ�`l�g�@"?7(5�3@r+�ΐ!?�������@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@�2�HѠٿ%F��J�@:��@��3@�����!?ˠ�6���@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@ڪf��ٿ�������@��^�3@����!?R��1��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@���k�ٿ�Ԏ'�@�mw��3@�G�D2�!?�"�Y��@a[�#�ٿXO^�k�@^��D�3@^V��ߐ!?�&={��@a[�#�ٿXO^�k�@^��D�3@^V��ߐ!?�&={��@a[�#�ٿXO^�k�@^��D�3@^V��ߐ!?�&={��@U�l�ٿ�A5��@� �N��3@��Ð!? j&S�'�@U�l�ٿ�A5��@� �N��3@��Ð!? j&S�'�@U�l�ٿ�A5��@� �N��3@��Ð!? j&S�'�@���Bp�ٿ���@!��@Iބ\�3@�j#N�!?G�(3C�@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@����z�ٿ�=�iX�@���p�3@b42h4�!?�QE{>��@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@��}Z�ٿ��3��*�@ך�ai�3@c�j�!?�ˢ��/�@0��*o�ٿ���Z���@W���k�3@
2N���!?�ަ�v]�@K��ٿߣ����@ �r�3@�c�!?!�,ɏ��@<�5ڴ�ٿ�)��]��@|�a��3@�y-Ր!?ʋSO��@<�5ڴ�ٿ�)��]��@|�a��3@�y-Ր!?ʋSO��@<�5ڴ�ٿ�)��]��@|�a��3@�y-Ր!?ʋSO��@<�5ڴ�ٿ�)��]��@|�a��3@�y-Ր!?ʋSO��@<�5ڴ�ٿ�)��]��@|�a��3@�y-Ր!?ʋSO��@2U%g�ٿN-�u�@9 ���3@�&?N�!?o�6�9�@2U%g�ٿN-�u�@9 ���3@�&?N�!?o�6�9�@2U%g�ٿN-�u�@9 ���3@�&?N�!?o�6�9�@	�V}*�ٿ� ���@�?���3@#~�$�!?�~]���@��
���ٿ�ӞH�#�@O�	��3@a��!?�C� #��@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@��j�ٿ3{�P�|�@$V��,�3@�S_���!?3�!W`�@���/�ٿ�$l{�@�늏��3@�"���!?-Lܯ��@S���ٿ�-P�@TԜw�3@|��2ѐ!?<籋���@S���ٿ�-P�@TԜw�3@|��2ѐ!?<籋���@S���ٿ�-P�@TԜw�3@|��2ѐ!?<籋���@S���ٿ�-P�@TԜw�3@|��2ѐ!?<籋���@S���ٿ�-P�@TԜw�3@|��2ѐ!?<籋���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@,��F�ٿ�7�e��@kKW���3@����͐!?S�C���@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@#Nz���ٿKk��kK�@��1�3@5�ΐ!?�)�Ł��@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�W��Y�ٿ��=Ԩ��@�A�0�3@�VbGƐ!?��w���@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@�h��-�ٿ�P��ߛ�@��/m1�3@Kj�罐!?~�(�!��@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@U�*�E�ٿ}����@�n�q�3@�"t��!?-�2f)�@��.^�ٿ�!I :�@Ď���3@	�A�!?�����@��.^�ٿ�!I :�@Ď���3@	�A�!?�����@��.^�ٿ�!I :�@Ď���3@	�A�!?�����@��.^�ٿ�!I :�@Ď���3@	�A�!?�����@����àٿSq?#�@�f���3@�C�`�!?FM�u��@����àٿSq?#�@�f���3@�C�`�!?FM�u��@a=��P�ٿ�:ӵV��@M���3@V�f��!?z@��gE�@a=��P�ٿ�:ӵV��@M���3@V�f��!?z@��gE�@a=��P�ٿ�:ӵV��@M���3@V�f��!?z@��gE�@^��V�ٿ &���,�@��+���3@~���!?������@^��V�ٿ &���,�@��+���3@~���!?������@�����ٿ�8{�h�@ݹ]���3@=�Gʐ!?ޭ����@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@q6��G�ٿ��p���@�ꤞ�3@i^{c��!?�Ɉ�q*�@T�乡ٿ��1� �@>��3@���!?H.7��%�@T�P� �ٿ���O�@8p�
�3@�M՚�!?�:��5��@T�P� �ٿ���O�@8p�
�3@�M՚�!?�:��5��@T�P� �ٿ���O�@8p�
�3@�M՚�!?�:��5��@T�P� �ٿ���O�@8p�
�3@�M՚�!?�:��5��@��{�i�ٿ,|�1�T�@Ӱp���3@���$ː!?$�C �@|K�j��ٿ�,�%��@��X��3@�ꤞ�!?�A�#"��@|K�j��ٿ�,�%��@��X��3@�ꤞ�!?�A�#"��@|K�j��ٿ�,�%��@��X��3@�ꤞ�!?�A�#"��@o���ٿ"�p�z�@<�Ԏ��3@�;Rq��!?CC�y�@o���ٿ"�p�z�@<�Ԏ��3@�;Rq��!?CC�y�@o���ٿ"�p�z�@<�Ԏ��3@�;Rq��!?CC�y�@o���ٿ"�p�z�@<�Ԏ��3@�;Rq��!?CC�y�@l\ �e�ٿ���L��@W�G�	�3@�vBп�!?�����S�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@�-Ǩ�ٿ�-�_��@B�)���3@���	��!?��Lܕ�@<�U⚠ٿ=���K@�@�W9�l�3@������!?����.��@<�U⚠ٿ=���K@�@�W9�l�3@������!?����.��@\�ϑ'�ٿN_/R�@ij�K|�3@�u����!?/�A���@\�ϑ'�ٿN_/R�@ij�K|�3@�u����!?/�A���@~=���ٿ�B����@u����3@��t�!?�5�����@~=���ٿ�B����@u����3@��t�!?�5�����@~=���ٿ�B����@u����3@��t�!?�5�����@~=���ٿ�B����@u����3@��t�!?�5�����@~=���ٿ�B����@u����3@��t�!?�5�����@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@rL�N�ٿ*LghU��@R~۔��3@5��G�!?*¥���@3-�O�ٿH��"��@�*�JY�3@wI'�!?�0W���@	9��ٿS��\�[�@�jI�3@����!?"7'B��@	9��ٿS��\�[�@�jI�3@����!?"7'B��@	9��ٿS��\�[�@�jI�3@����!?"7'B��@��!{�ٿ%��|!��@?�҆��3@� 3Jΐ!?�P�'Q�@��!{�ٿ%��|!��@?�҆��3@� 3Jΐ!?�P�'Q�@��!{�ٿ%��|!��@?�҆��3@� 3Jΐ!?�P�'Q�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@��o7�ٿa�O'n�@�U8؍�3@DO^ ɐ!?��.3^�@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@�u�vx�ٿ��eHa��@T�w���3@~Dbː!?i�o$��@ʾ�h��ٿ����@����3@K���!?�CΣ�#�@��Jݝٿ��s��@����3@I��[��!?p�'���@��Jݝٿ��s��@����3@I��[��!?p�'���@��Jݝٿ��s��@����3@I��[��!?p�'���@Ʒ�ɳ�ٿY�T��@66�;�3@�f&ܐ!?~�o��`�@��歟�ٿ�l�#��@Y����3@��/��!?�ыk�S�@��歟�ٿ�l�#��@Y����3@��/��!?�ыk�S�@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@Dz��ڥٿ�V/yε�@:._r�3@0-�A��!?q�q�M��@G*+�ٿ� �dOL�@:q����3@({�yk�!?�����@G*+�ٿ� �dOL�@:q����3@({�yk�!?�����@�7\�ٿ*�z�Q	�@�Gm���3@g�͐!?R�ء��@�7\�ٿ*�z�Q	�@�Gm���3@g�͐!?R�ء��@d����ٿ�?����@����3@`O�ب�!?�&�Fa,�@d����ٿ�?����@����3@`O�ب�!?�&�Fa,�@d����ٿ�?����@����3@`O�ب�!?�&�Fa,�@)��ٿ&w���@��h#V�3@��Đ!?(v֧��@)��ٿ&w���@��h#V�3@��Đ!?(v֧��@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@p�f�c�ٿ����,�@�&�w�3@-jK��!?؎�����@��>��ٿ7�^o6�@�:��|�3@v�ȅ	�!?sW.'"��@c�>�S�ٿ�;����@�����3@rzz'��!?>w�?
��@c�>�S�ٿ�;����@�����3@rzz'��!?>w�?
��@c�>�S�ٿ�;����@�����3@rzz'��!?>w�?
��@6�uۛٿŨ��ַ�@@p�i�3@�Y��!?G�b�O�@6�uۛٿŨ��ַ�@@p�i�3@�Y��!?G�b�O�@6�uۛٿŨ��ַ�@@p�i�3@�Y��!?G�b�O�@6�uۛٿŨ��ַ�@@p�i�3@�Y��!?G�b�O�@BK�ٿ^�Zx���@�먄��3@��o�y�!?/�Y�U�@xNcl�ٿp�N���@}T��3@"2٩o�!?"�ya��@xNcl�ٿp�N���@}T��3@"2٩o�!?"�ya��@���,�ٿ�Z4p�@�a����3@�DU���!?6.���@���,�ٿ�Z4p�@�a����3@�DU���!?6.���@���,�ٿ�Z4p�@�a����3@�DU���!?6.���@��l��ٿk�+~]�@�a1ɍ�3@bq	c�!?1Q�.-:�@��l��ٿk�+~]�@�a1ɍ�3@bq	c�!?1Q�.-:�@�<�X�ٿ�S-�Ɩ�@pS��.�3@wch�ݐ!?$)���@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�>�8ԥٿ!�؏���@h|�M&�3@A�Yް�!?cV쁿u�@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@�5i&�ٿ�N��L��@�t^X
�3@{[J�$�!?W-�Չ��@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@bj�֚ٿdkS_!�@@,Ub�3@i�9���!?U�6K!>�@��z�ٿi��� ��@mUYE��3@(T;`��!?�\�8��@��z�ٿi��� ��@mUYE��3@(T;`��!?�\�8��@��z�ٿi��� ��@mUYE��3@(T;`��!?�\�8��@��z�ٿi��� ��@mUYE��3@(T;`��!?�\�8��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@%ōa��ٿ��/%r�@�u��g�3@q�l'�!?�7ơ��@R�}�?�ٿz�\�R'�@~����3@�'lSÐ!?+�y)�@�S�ٿ���g��@]��)�3@ˍ��+�!?�Tڦ�@�S�ٿ���g��@]��)�3@ˍ��+�!?�Tڦ�@�S�ٿ���g��@]��)�3@ˍ��+�!?�Tڦ�@�S�ٿ���g��@]��)�3@ˍ��+�!?�Tڦ�@�S�ٿ���g��@]��)�3@ˍ��+�!?�Tڦ�@H@���ٿ�d�V��@�����3@�Z�j5�!?����}��@�A/�[�ٿ�f7kͧ�@��mD�3@ W+�!?��l�S�@�A/�[�ٿ�f7kͧ�@��mD�3@ W+�!?��l�S�@Lz�P��ٿt�S��C�@@E	�3@��#��!?�
���.�@���b��ٿ�v\�J��@�YƎ�3@�ܷR��!?a Q���@R�SP(�ٿ` \y�9�@zr�v!�3@��U�!?\x��n��@R�SP(�ٿ` \y�9�@zr�v!�3@��U�!?\x��n��@R�SP(�ٿ` \y�9�@zr�v!�3@��U�!?\x��n��@R�SP(�ٿ` \y�9�@zr�v!�3@��U�!?\x��n��@R�SP(�ٿ` \y�9�@zr�v!�3@��U�!?\x��n��@�w�ۂ�ٿ��eg!�@�3+`h�3@�_��s�!?���a�@�w�ۂ�ٿ��eg!�@�3+`h�3@�_��s�!?���a�@�w�ۂ�ٿ��eg!�@�3+`h�3@�_��s�!?���a�@�w�ۂ�ٿ��eg!�@�3+`h�3@�_��s�!?���a�@���<F�ٿ�sLY�D�@�-��N�3@��^Ɠ�!?���g*��@���<F�ٿ�sLY�D�@�-��N�3@��^Ɠ�!?���g*��@fk?�ٿ{$�d��@���2A�3@=c�!��!?���{���@fk?�ٿ{$�d��@���2A�3@=c�!��!?���{���@fk?�ٿ{$�d��@���2A�3@=c�!��!?���{���@fk?�ٿ{$�d��@���2A�3@=c�!��!?���{���@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@�ڏ�+�ٿ�|{��@!��l�3@�1��!?1��@��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@%py���ٿ^壟 ��@V�X?��3@��B��!?�_�.(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@
��l��ٿ�|�� ��@(ṏ��3@B�x��!?���(��@������ٿ���� ��@;Q����3@:�����!?��$4(��@������ٿ���� ��@;Q����3@:�����!?��$4(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@E!�f��ٿ��z� ��@��9%��3@�m��!?B"MN(��@<�SΩ�ٿ�C� ��@�+,i��3@w?��!?�3%@(��@<�SΩ�ٿ�C� ��@�+,i��3@w?��!?�3%@(��@V^Wo��ٿ�˙� ��@�Y����3@��u�!?�1Q(��@V^Wo��ٿ�˙� ��@�Y����3@��u�!?�1Q(��@V^Wo��ٿ�˙� ��@�Y����3@��u�!?�1Q(��@V^Wo��ٿ�˙� ��@�Y����3@��u�!?�1Q(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@�L��ٿ/R�� ��@��e��3@����!?�	�N(��@��p��ٿ⑅� ��@�0���3@���N�!?+�RM(��@��p��ٿ⑅� ��@�0���3@���N�!?+�RM(��@��p��ٿ⑅� ��@�0���3@���N�!?+�RM(��@'m��ٿw�i� ��@1�����3@�H��3�!?��@S(��@'m��ٿw�i� ��@1�����3@�H��3�!?��@S(��@	W8��ٿ�WU� ��@������3@v���!?�y�P(��@	W8��ٿ�WU� ��@������3@v���!?�y�P(��@�%<���ٿ��ً ��@���$��3@GW$(��!?���K(��@KY�5��ٿ"��� ��@Ȇ���3@�c:��!?��^(��@KY�5��ٿ"��� ��@Ȇ���3@�c:��!?��^(��@KY�5��ٿ"��� ��@Ȇ���3@�c:��!?��^(��@"�+��ٿ�@?� ��@IX-��3@�♧�!?��\(��@"�+��ٿ�@?� ��@IX-��3@�♧�!?��\(��@"�+��ٿ�@?� ��@IX-��3@�♧�!?��\(��@��˴�ٿ��.� ��@�����3@Nm�̕�!?;�Bb(��@��∬�ٿE�� ��@x�1��3@1�̐!? I�](��@dj�짚ٿ�l�� ��@����3@���!?�ga(��@dj�짚ٿ�l�� ��@����3@���!?�ga(��@u�}̪�ٿ�2�� ��@�����3@�d�ؐ!?B��`(��@u�}̪�ٿ�2�� ��@�����3@�d�ؐ!?B��`(��@q�x���ٿA"D� ��@Wm����3@R�!֐!?!��h(��@q�x���ٿA"D� ��@Wm����3@R�!֐!?!��h(��@q�x���ٿA"D� ��@Wm����3@R�!֐!?!��h(��@q�x���ٿA"D� ��@Wm����3@R�!֐!?!��h(��@P���ٿ�� ��@&��8��3@#�p��!?"+�`(��@���ٿ �d� ��@9�e��3@�
HS��!?�J[W(��@���ٿ �d� ��@9�e��3@�
HS��!?�J[W(��@���ٿ �d� ��@9�e��3@�
HS��!?�J[W(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@��9���ٿ�zS� ��@�� ���3@/��Ɛ!?��Y(��@�a����ٿ8�� ��@�uB��3@�uG��!?��`(��@w|�⩚ٿ�� ��@��=���3@izc��!?��i(��@w|�⩚ٿ�� ��@��=���3@izc��!?��i(��@��:��ٿt�� ��@.Z���3@�nID�!?��ho(��@RtzƢ�ٿf ��@�qФ��3@�\�L�!?=�r(��@RtzƢ�ٿf ��@�qФ��3@�\�L�!?=�r(��@RtzƢ�ٿf ��@�qФ��3@�\�L�!?=�r(��@RtzƢ�ٿf ��@�qФ��3@�\�L�!?=�r(��@���&��ٿ��� ��@��C���3@M6�]m�!?��Rs(��@���&��ٿ��� ��@��C���3@M6�]m�!?��Rs(��@>b=٤�ٿvM�� ��@/�N���3@�f�֢�!?�p�t(��@�#飚ٿ�@� ��@�S�T��3@�PՐ!?��{(��@�#飚ٿ�@� ��@�S�T��3@�PՐ!?��{(��@�#飚ٿ�@� ��@�S�T��3@�PՐ!?��{(��@�g�g��ٿ�� ��@Nh����3@�vN��!?�'Lu(��@�g�g��ٿ�� ��@Nh����3@�vN��!?�'Lu(��@���J��ٿ)R� ��@�p@��3@�Gg�!?=~v(��@���J��ٿ)R� ��@�p@��3@�Gg�!?=~v(��@���J��ٿ)R� ��@�p@��3@�Gg�!?=~v(��@1�0᠚ٿ��� ��@�W���3@-쨦��!?��z(��@1�0᠚ٿ��� ��@�W���3@-쨦��!?��z(��@��/��ٿ�d�� ��@�"����3@�JeX<�!?�C�|(��@���ٿ�?ė ��@�ޖG��3@2�|�-�!?��(��@���ٿ�?ė ��@�ޖG��3@2�|�-�!?��(��@���ٿ�?ė ��@�ޖG��3@2�|�-�!?��(��@���ٿ�?ė ��@�ޖG��3@2�|�-�!?��(��@�z\T��ٿ��m� ��@����3@R�z	1�!?����(��@���頚ٿT2�� ��@�0����3@�'��!?(��(��@���頚ٿT2�� ��@�0����3@�'��!?(��(��@L΅v��ٿ���� ��@������3@@�ʟ�!?�=�(��@V��7��ٿ�s%� ��@�j����3@��J@T�!?z>Έ(��@V��7��ٿ�s%� ��@�j����3@��J@T�!?z>Έ(��@���ٿ�៖ ��@�����3@/A�)�!?/�h�(��@��$���ٿ�VƓ ��@�����3@�pF�!?&!ۑ(��@��$���ٿ�VƓ ��@�����3@�pF�!?&!ۑ(��@�����ٿ�֏ ��@����3@b	�L0�!?wf�(��@��T��ٿ�
�� ��@�����3@�\O�8�!?�mɘ(��@?>I��ٿ��	� ��@IW���3@�'""��!?��N�(��@��᠚ٿŭ� ��@2M���3@O�����!?
�'�(��@��᠚ٿŭ� ��@2M���3@O�����!?
�'�(��@�W�Ȣ�ٿ�8� ��@swM��3@A��!?�VK�(��@�W�Ȣ�ٿ�8� ��@swM��3@A��!?�VK�(��@ޞ30��ٿ��� ��@N�5O��3@���ʫ�!?c1��(��@ޞ30��ٿ��� ��@N�5O��3@���ʫ�!?c1��(��@ޞ30��ٿ��� ��@N�5O��3@���ʫ�!?c1��(��@ޞ30��ٿ��� ��@N�5O��3@���ʫ�!?c1��(��@ޞ30��ٿ��� ��@N�5O��3@���ʫ�!?c1��(��@��U+��ٿ�{�� ��@ROi���3@D��͐!?_�]�(��@ȅbA��ٿG�U� ��@4t�;��3@s>if��!?'�(��@Lg�
��ٿx)�� ��@ؕ�G��3@�o��!?�f��(��@�%��ٿ�\ˎ ��@z=C��3@�`%�!?�X�(��@q�����ٿ�N� ��@�����3@4���!?�(��@q�����ٿ�N� ��@�����3@4���!?�(��@�H�a��ٿ�Zh� ��@�h��3@PY��!?�X]{(��@�H�a��ٿ�Zh� ��@�h��3@PY��!?�X]{(��@��n���ٿ�_� ��@�	iI��3@XI�!?Ղ��(��@m݂���ٿW�Đ ��@�dPi��3@1�oƸ�!?^�Ή(��@K�-�ٿ/@�� ��@��p���3@�BА!?��΃(��@�]���ٿo�h� ��@����3@�����!?����(��@=�B蔚ٿi0Q� ��@}�����3@���!?W/=�(��@,�c���ٿI�m� ��@9�.���3@��ͻ��!?�"��(��@vp�w��ٿ_��� ��@�y����3@�ԇǐ!?��Ն(��@vp�w��ٿ_��� ��@�y����3@�ԇǐ!?��Ն(��@R����ٿ�:�� ��@�����3@H��!?��H�(��@R����ٿ�:�� ��@�����3@H��!?��H�(��@�.�Ș�ٿ%�.� ��@B�Fj��3@?�����!?����(��@ao���ٿ��� ��@\�y���3@�(�Eʐ!?�f��(��@��L���ٿX�s� ��@��Md��3@��ΐ!?a��(��@�ٿ�2�� ��@��r��3@��i��!?H(k�(��@�
�d��ٿE��� ��@+ݞ���3@��O��!?!�Ē(��@!����ٿ�<� ��@�<���3@vX���!?�e�(��@�ځ<��ٿS�� ��@�jJ���3@>�ʣ �!?��}�(��@o�vq��ٿ���� ��@������3@����ݐ!?Ҕ��(��@��a���ٿ��X� ��@���3@�O��Ԑ!?!�k�(��@RqS���ٿ�Aȗ ��@a�����3@�ۗh��!?�B��(��@QX"���ٿ��� ��@�ip��3@��i���!?.��(��@QX"���ٿ��� ��@�ip��3@��i���!?.��(��@��rٿp֞� ��@Y�A��3@���梐!?�}�(��@�Z����ٿ�j� ��@<>���3@��]�ː!?ߣډ(��@Ku�b��ٿ�Ⲝ ��@�Tr|��3@�s0�!?��ّ(��@�+�7��ٿI� ��@_͛���3@�(�͐!?�Pڍ(��@W'��ٿc�0� ��@����3@����!?�W�(��@W'��ٿc�0� ��@����3@����!?�W�(��@�Iw���ٿr�ף ��@�˨`��3@�$��ʐ!?��p�(��@�����ٿy�� ��@`t�6��3@:5@�
�!?�d)�(��@�����ٿy�� ��@`t�6��3@:5@�
�!?�d)�(��@���
��ٿ�� ��@��}��3@~�94��!?u��(��@˂��ٿ��� ��@?EC���3@$!-���!?�A�(��@4{�y��ٿ�vy� ��@<.����3@�z
��!?�	�(��@7�D��ٿ���� ��@q���3@�+����!?/� �(��@�{���ٿ���� ��@��ԗ��3@��l�Ր!?�?ɞ(��@��E醚ٿ��q� ��@᧤���3@Kx∷�!?��(��@�����ٿImn� ��@������3@;����!?-���(��@t�����ٿ�"�� ��@Uc����3@2�R]��!? ��(��@t�����ٿ�"�� ��@Uc����3@2�R]��!? ��(��@t�����ٿ�"�� ��@Uc����3@2�R]��!? ��(��@t�����ٿ�"�� ��@Uc����3@2�R]��!? ��(��@��?��ٿ��_� ��@,�%���3@�X(Z��!?���(��@�����ٿ-χ� ��@�A�!��3@�o)�!?�o�(��@�����ٿ-χ� ��@�A�!��3@�o)�!?�o�(��@!��+��ٿք�� ��@I�!��3@�K3��!??�(��@!��+��ٿք�� ��@I�!��3@�K3��!??�(��@����ٿ��j� ��@+�(���3@�d����!?:{�(��@��,ږ�ٿU=�� ��@�-@���3@�z�ސ!?���(��@��,ږ�ٿU=�� ��@�-@���3@�z�ސ!?���(��@�*8Ӛ�ٿ�B� ��@`�M��3@/��ܐ!?�i�(��@�N���ٿ��� ��@��3���3@�m���!?�5��(��@��Dn��ٿle�� ��@�����3@�}����!?�F�(��@B��4��ٿ�t� ��@�����3@�VHݐ!?�l�(��@B��4��ٿ�t� ��@�����3@�VHݐ!?�l�(��@���Ꟛٿ��a� ��@�ھ���3@����!?
t�(��@���Ꟛٿ��a� ��@�ھ���3@����!?
t�(��@���Ꟛٿ��a� ��@�ھ���3@����!?
t�(��@���Ꟛٿ��a� ��@�ھ���3@����!?
t�(��@���Ꟛٿ��a� ��@�ھ���3@����!?
t�(��@�P�-��ٿ�8L� ��@J0<���3@����!?
W͝(��@�P�-��ٿ�8L� ��@J0<���3@����!?
W͝(��@��|��ٿc� ��@�z7���3@�V8iJ�!?�(Ϣ(��@�j��ٿ�)�� ��@OK���3@8J�.�!?��	�(��@� ���ٿ�m�� ��@�u���3@�k�]'�!?�#p�(��@�x� ��ٿD�Ԕ ��@%�t��3@���p�!?�k�(��@>�R��ٿ��� ��@�z3��3@j���v�!?�خ�(��@��G��ٿ�!�� ��@J�C���3@e*i�g�!?��(��@L�tY��ٿek� ��@��(���3@*��j)�!?S���(��@L�tY��ٿek� ��@��(���3@*��j)�!?S���(��@5�	���ٿ�,� ��@�F&��3@�HY�!?߲(��@�n�p��ٿ���� ��@��%��3@C�!ڐ!?���(��@��[���ٿ��� ��@EFY���3@����!?~�j�(��@�!蚚ٿ΍� ��@�d�I��3@�^t��!?k���(��@�!蚚ٿ΍� ��@�d�I��3@�^t��!?k���(��@�!蚚ٿ΍� ��@�d�I��3@�^t��!?k���(��@�!蚚ٿ΍� ��@�d�I��3@�^t��!?k���(��@��+&��ٿ�� ��@�i����3@��}��!?+4a�(��@��+&��ٿ�� ��@�i����3@��}��!?+4a�(��@GZ�>��ٿ�#� ��@�����3@��x�!?��E�(��@GZ�>��ٿ�#� ��@�����3@��x�!?��E�(��@GZ�>��ٿ�#� ��@�����3@��x�!?��E�(��@P�on��ٿ���� ��@]�O���3@z�=�Ɛ!?]��(��@��Ν�ٿ���� ��@�ׂ��3@?�縷!?�w�(��@lM䢚ٿ!�� ��@(�1f��3@@�0���!?u�s�(��@D��Ǧ�ٿwY� ��@�ҹ���3@�ؑ�͐!?���(��@�/u��ٿ�Dk� ��@t�����3@�OȐ!?L��(��@R����ٿ�Ր ��@Bn�r��3@7VJ��!?+k�(��@��^"��ٿx�� ��@�P���3@��2�ې!?bƃ�(��@@l��ٿ*�-� ��@��Y{��3@�>c*�!?4�#�(��@@l��ٿ*�-� ��@��Y{��3@�>c*�!?4�#�(��@Zm�K��ٿe�� ��@���U��3@��?��!?+���(��@�R=���ٿ�8 ��@�SA7��3@�5�Wʐ!?�
)��@�$9㭚ٿ]�^} ��@0a�%��3@� �_��!?��m�(��@��8��ٿ���� ��@�)<��3@��R��!?��d�(��@��V1��ٿO= � ��@�����3@u93xӐ!?V���(��@��V1��ٿO= � ��@�����3@u93xӐ!?V���(��@�z����ٿ��4� ��@��i���3@��&˷�!?(Ʋ(��@��H���ٿA��� ��@����3@e�%!?�B�(��@�l�n��ٿ�ʓ ��@>�{��3@���>��!?eKJ�(��@��՟�ٿ4F� ��@d�v���3@c*�S��!?N�(��@������ٿ��0� ��@���|��3@�?��!?�V�(��@c��Q��ٿ/�� ��@�|O��3@i�5 ː!?�٦�(��@�k� ��ٿ�9� ��@I�����3@��g&ɐ!?� :�(��@�k� ��ٿ�9� ��@I�����3@��g&ɐ!?� :�(��@�k� ��ٿ�9� ��@I�����3@��g&ɐ!?� :�(��@}'����ٿ3�� ��@����3@踣ؐ!?��v�(��@}'����ٿ3�� ��@����3@踣ؐ!?��v�(��@}'����ٿ3�� ��@����3@踣ؐ!?��v�(��@<
t��ٿ��� ��@,����3@܇:|ސ!?�Z*�(��@�ė���ٿ�O`z ��@G��
��3@�b�fڐ!?`$�(��@�;_��ٿ(�a| ��@N���3@�����!?���(��@3����ٿH�&� ��@\So���3@�]}P�!?���(��@Z��,��ٿ��o� ��@j�	��3@�]�%�!?%2b�(��@<Z$j��ٿF=� ��@�BA��3@l��0�!?; �(��@����ٿbs� ��@�r���3@7�:V�!?R�o�(��@����ٿbs� ��@�r���3@7�:V�!?R�o�(��@����ٿbs� ��@�r���3@7�:V�!?R�o�(��@f��c��ٿ6%� ��@�����3@Z�r*�!?� )�(��@s1ዝ�ٿ �� ��@���-��3@�W��!?�	��(��@1?���ٿd�� ��@�Ou��3@P�m���!?2*g�(��@�YJE��ٿ� � ��@1�`���3@Zc����!?�g)�(��@"F[���ٿ-�� ��@Ǟ����3@��4�k�!?d�&�(��@"F[���ٿ-�� ��@Ǟ����3@��4�k�!?d�&�(��@��8��ٿ�<�� ��@	S�Z��3@m%L�b�!?FK��(��@I�����ٿ��
� ��@�*6R��3@�#��!?ғ��(��@I�����ٿ��
� ��@�*6R��3@�#��!?ғ��(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@@��$��ٿQ�� ��@�+6���3@mh%��!?����(��@ч��ٿ�cq� ��@"��;��3@q��ˏ�!?��(��@D�����ٿ{�r ��@�n���3@G��u�!?�D��(��@t����ٿ/�'v ��@�>���3@���3�!?Y�e)��@t����ٿ/�'v ��@�>���3@���3�!?Y�e)��@*zr��ٿ�N�q ��@�L�Z��3@��*!,�!?���)��@*zr��ٿ�N�q ��@�L�Z��3@��*!,�!?���)��@r�׫�ٿ��i ��@�;���3@i��A�!?O6\:)��@/|��ٿ�hn~ ��@�����3@ W&H�!?	B�(��@/|��ٿ�hn~ ��@�����3@ W&H�!?	B�(��@/|��ٿ�hn~ ��@�����3@ W&H�!?	B�(��@/|��ٿ�hn~ ��@�����3@ W&H�!?	B�(��@d����ٿ��#� ��@�s���3@|�]L��!?���(��@p���ٿ�{�� ��@3Z4Z��3@�����!?�4�(��@��n��ٿ��� ��@W�ު��3@�C�W��!?/��(��@Q����ٿ��O� ��@�b^��3@A1Ypߐ!?���(��@$8�]��ٿ�� ��@�O���3@I��!?Ɋ��(��@f�����ٿ��B� ��@����3@�����!?�5}(��@gu���ٿ�̪ ��@F6d$��3@ay2Đ!?���Y(��@�����ٿ,,l� ��@ �d��3@,Hp�!?:F�[(��@�Nu��ٿ�C۬ ��@*����3@��~ ʐ!?4��g(��@�Nu��ٿ�C۬ ��@*����3@��~ ʐ!?4��g(��@�Nu��ٿ�C۬ ��@*����3@��~ ʐ!?4��g(��@g��2��ٿ샊� ��@N�=���3@'�_q�!?W��E(��@������ٿuk� ��@�+���3@�y��ې!?��:d(��@�2h��ٿШ� ��@:�J|��3@7vK��!?�K(��@�2h��ٿШ� ��@:�J|��3@7vK��!?�K(��@v����ٿ퀻� ��@�=���3@�,6ڞ�!?�=�](��@�C�[��ٿ�-&� ��@��c��3@
�9w��!?ª�](��@|A���ٿC�ڨ ��@;��*��3@��eO��!?>��}(��@ht�;��ٿ��� ��@���3@Mt�z�!?`��w(��@�=��}�ٿFRl� ��@�h(���3@!�Ƅ�!?։`(��@�>�
��ٿ�ꎮ ��@��j���3@�(]��!?DO�(��@�>�
��ٿ�ꎮ ��@��j���3@�(]��!?DO�(��@�m�8��ٿ;�5� ��@p�~��3@�a����!?ʀJ�(��@�m�8��ٿ;�5� ��@p�~��3@�a����!?ʀJ�(��@��À��ٿ���� ��@�3l��3@qƆ��!?��G�(��@��À��ٿ���� ��@�3l��3@qƆ��!?��G�(��@r?��Кٿ6G�; ��@�d(��3@N��9ϐ!?`��)��@���ǚٿ�5�Q ��@қ1y��3@���ɐ!?�{W6)��@���ǚٿ�5�Q ��@қ1y��3@���ɐ!?�{W6)��@a��|��ٿq|o ��@2/4S��3@�I2�!?sq��(��@.�Śٿ�c�X ��@�	�c��3@7n�p�!?c��")��@��Z֚ٿ�I�; ��@��4���3@�$��!?F�Zo)��@�R����ٿ��r. ��@8�Cg��3@�y��!?#�G�)��@�(���ٿ~�� ��@�}M� 4@�-G�ΐ!?ը*��@�(���ٿ~�� ��@�}M� 4@�-G�ΐ!?ը*��@�(���ٿ~�� ��@�}M� 4@�-G�ΐ!?ը*��@��ٿ�F3����@���< 4@��h]��!?�p*��@��ٿ�F3����@���< 4@��h]��!?�p*��@� ��
�ٿ�O�����@ +�, 4@\e�Ȏ�!?�:#!*��@���DI�ٿ�v�����@G��� 4@��v'Ґ!?Jk��*��@���DI�ٿ�v�����@G��� 4@��v'Ґ!?Jk��*��@�{�ٿT������@<� 4@7]�##�!?����)��@��X�ٿ���}���@6�hc 4@�����!?X�+��@�c��A�ٿ.6D����@��� 4@&�4K��!?��R�*��@�c��A�ٿ.6D����@��� 4@&�4K��!?��R�*��@�c��A�ٿ.6D����@��� 4@&�4K��!?��R�*��@�"\�a�ٿ��3`���@_Wg� 4@q�Q֐!?w:+��@�P��ٿ�������@{�{�8 4@����	�!?���Y,��@�P��ٿ�������@{�{�8 4@����	�!?���Y,��@W��X�ٿҧ|���@��Y` 4@o58z#�!?m�f+��@]��ԛٿ*f|����@��[> 4@�����!?���,��@�#�P��ٿb����@�MT6 4@�2��ې!?݇}F,��@�#�P��ٿb����@�MT6 4@�2��ې!?݇}F,��@�#�P��ٿb����@�MT6 4@�2��ې!?݇}F,��@WP��h�ٿ��Z���@j߷�  4@+����!?P�?{+��@�2��}�ٿ���?���@�(% 4@�J�T��!?��=�+��@�2��}�ٿ���?���@�(% 4@�J�T��!?��=�+��@ţ���ٿ�;X���@��* 4@@M�y�!?m�c�+��@ţ���ٿ�;X���@��* 4@@M�y�!?m�c�+��@$7�ؚٿ��- ��@�mu���3@#�Do�!?�雺)��@$7�ؚٿ��- ��@�mu���3@#�Do�!?�雺)��@߹C��ٿ~���@�f��3@�g'�!?I�"�%��@-���ٿ��*���@3�*J��3@G�ݵ'�!?�>=p&��@R7b5��ٿD�#^ ��@�/����3@$=�m�!?_u�-)��@R7b5��ٿD�#^ ��@�/����3@$=�m�!?_u�-)��@R7b5��ٿD�#^ ��@�/����3@$=�m�!?_u�-)��@��D�ٿw�����@Gu�< 4@�����!?��*��@��E��ٿ��a����@�[�> 4@W�r�!?���,��@�p[+�ٿ� �:���@`�oT 4@gpqAu�!?��-��@=��}�ٿ���J���@�[YR 4@_�i㦐!?���-��@=��}�ٿ���J���@�[YR 4@_�i㦐!?���-��@=��}�ٿ���J���@�[YR 4@_�i㦐!?���-��@=��}�ٿ���J���@�[YR 4@_�i㦐!?���-��@=��}�ٿ���J���@�[YR 4@_�i㦐!?���-��@mm���ٿ�$�����@j�;HF 4@�ǿ}�!? �-��@��{f�ٿ�5`���@���� 4@��י�!?���;+��@Q���[�ٿ��� ��@uf|o��3@�[��m�!?e��'��@ؓ ��ٿ��Ͷ��@B��׭�3@6�*)ɐ!?V-�T&��@��Ǣ��ٿ�����@ �ܸ�3@7�X��!?�&�&��@�̢1�ٿ9Mʹ��@d�����3@�A�Z��!?n�4$��@�̢1�ٿ9Mʹ��@d�����3@�A�Z��!?n�4$��@�sz���ٿ�Fx��@�%ӟ�3@��hSѐ!?P���%��@�sz���ٿ�Fx��@�%ӟ�3@��hSѐ!?P���%��@I�69��ٿP�<� ��@�G�]��3@��$r��!?����(��@I�69��ٿP�<� ��@�G�]��3@��$r��!?����(��@N�_��ٿ��Y����@�s�  4@1�m*��!?Z{/�)��@��	�M�ٿ�v�����@�I� 4@��`�!?��G�*��@��	�M�ٿ�v�����@�I� 4@��`�!?��G�*��@��	�M�ٿ�v�����@�I� 4@��`�!?��G�*��@gV[��ٿ&�W����@�7��C 4@��א!?�b�,��@x����ٿ�%9s���@�3��G 4@Z���o�!?�tq'-��@]��қٿ�������@�G��0 4@,�ņ�!?a��,��@]��қٿ�������@�G��0 4@,�ņ�!?a��,��@ܺ��ٿ� ����@��Gr��3@F�MБ�!?��~S&��@w}1��ٿ2��� ��@~�����3@K���ސ!?����'��@w}1��ٿ2��� ��@~�����3@K���ސ!?����'��@��<�ٿ�&� ��@E43S��3@i&�!?���0)��@)�^f��ٿ� ��@|m���3@�'��א!?�X�B'��@ꦷ��ٿg�� ��@\�~���3@*l��!?`���'��@P$�s�ٿxJ���@��B���3@JT4F��!?GZ���@P$�s�ٿxJ���@��B���3@JT4F��!?GZ���@P$�s�ٿxJ���@��B���3@JT4F��!?GZ���@Y��\�ٿ�3P��@Oz�49�3@�L�1Đ!?��� ��@�H�1�ٿà/����@��b��3@-C{8��!?4��)��@�H�1�ٿà/����@��b��3@-C{8��!?4��)��@%--�ٿ��{��@��Ҳ�3@��G ��!?�S�&��@:��#O�ٿ��/0���@����M 4@�~�K�!?�u��,��@��,dʜٿ1�����@�$��m 4@tϪ+�!?��L4.��@��,dʜٿ1�����@�$��m 4@tϪ+�!?��L4.��@^�|��ٿn`�����@��4@�JmRl�!?�N6��@ŔwT��ٿwC8w���@�{�f� 4@��6��!?����2��@ŔwT��ٿwC8w���@�{�f� 4@��6��!?����2��@I+�m��ٿ1�6)���@i��&4@������!?ⶺ;6��@��Fb��ٿKR�U���@�۹� 4@�ѣݐ!?nA�0��@4�>�4�ٿ���@D�E�/ 4@Yt���!?GR��*��@4�>�4�ٿ���@D�E�/ 4@Yt���!?GR��*��@�g���ٿ�b<j ��@�#q��3@Q�z��!?{J��&��@�����ٿת���@�RuJ�3@��홐!?�8��!��@[�j��ٿ�ǅ��@����3@��]��!?�̻b��@v�����ٿ��	��@+y7�3@�܎U��!?��K���@?"���ٿ$�����@%do��3@F���Y�!?6��P��@?"���ٿ$�����@%do��3@F���Y�!?6��P��@�y�'��ٿ|��V��@��Ki�3@˴`�!?m̙��@�y�'��ٿ|��V��@��Ki�3@˴`�!?m̙��@G�`�ەٿ��L��@�{�?^�3@౷TP�!?��g��@G�`�ەٿ��L��@�{�?^�3@౷TP�!?��g��@��P�p�ٿ2�*���@�t`���3@F�mL��!?�3���@#�Z0��ٿ�ȿ���@�G�,�3@�̜�!?FB�I ��@��:sΜٿ�X����@<2��M 4@y����!?�Ɵ)-��@��:sΜٿ�X����@<2��M 4@y����!?�Ɵ)-��@��:sΜٿ�X����@<2��M 4@y����!?�Ɵ)-��@O�鵛ٿ��	g���@�Ȁ���3@R�ғ�!?��M(��@O�鵛ٿ��	g���@�Ȁ���3@R�ғ�!?��M(��@O�鵛ٿ��	g���@�Ȁ���3@R�ғ�!?��M(��@l�
�c�ٿ������@t`�s 4@0B@�|�!?:�[/��@l�
�c�ٿ������@t`�s 4@0B@�|�!?:�[/��@l�
�c�ٿ������@t`�s 4@0B@�|�!?:�[/��@l�
�c�ٿ������@t`�s 4@0B@�|�!?:�[/��@b&{eu�ٿP��A���@|��ċ 4@UܦU��!?� 0��@b&{eu�ٿP��A���@|��ċ 4@UܦU��!?� 0��@b&{eu�ٿP��A���@|��ċ 4@UܦU��!?� 0��@b&{eu�ٿP��A���@|��ċ 4@UܦU��!?� 0��@1-i�m�ٿ8� ��@R����3@�DQg��!?M�s�'��@�Fεۡٿ�������@�6{�4@������!?�F�{<��@�[����ٿ𮢗���@Ƚ�x4@Z �䐐!?D�!/5��@W�l.��ٿ,��c���@�����3@�|lB��!?���X(��@W�l.��ٿ,��c���@�����3@�|lB��!?���X(��@�Dv�~�ٿU�����@O(*~� 4@*�.]�!?��.��@�E���ٿ��@���@1ze3�3@��er��!?%�D���@�E���ٿ��@���@1ze3�3@��er��!?%�D���@�7cޤ�ٿeax� ��@��M���3@gh��!?+=�N%��@�7cޤ�ٿeax� ��@��M���3@gh��!?+=�N%��@�7cޤ�ٿeax� ��@��M���3@gh��!?+=�N%��@�7cޤ�ٿeax� ��@��M���3@gh��!?+=�N%��@�s�,�ٿy%�!���@�#qJ4@Z�u�u�!?�V�:4��@�H"o�ٿJ�Φ ��@�I��< 4@����Ӑ!?���*��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Po����ٿ�I� ��@��� 4@s�JȐ!?�5��-��@Z����ٿ�j�����@�L�C4@P����!?6���7��@���i�ٿ��+���@�Y�=p 4@����א!?Ɖ��.��@�� ���ٿ�^�|���@6�?�4@FH;vϐ!?���;��@I���D�ٿ���x��@���C�3@/�u��!?��5r��@��9�ٿp�I����@�cU�� 4@�J���!?ݒ�.��@��9�ٿp�I����@�cU�� 4@�J���!?ݒ�.��@��9�ٿp�I����@�cU�� 4@�J���!?ݒ�.��@j�M�ٿe2�����@�s��4@Ga���!?�f�7��@�{G'd�ٿn֒����@��D5�4@2�s��!? Kd7?��@�{G'd�ٿn֒����@��D5�4@2�s��!? Kd7?��@�B���ٿ��X2���@;A�z�4@��#1ڐ!?i`N>8��@�B���ٿ��X2���@;A�z�4@��#1ڐ!?i`N>8��@a�j�P�ٿ.�d���@� ��4@w���!?�ZX4��@a�j�P�ٿ.�d���@� ��4@w���!?�ZX4��@�w1D��ٿ���u��@�O~!� 4@P]H���!?@��,��@�w1D��ٿ���u��@�O~!� 4@P]H���!?@��,��@�w1D��ٿ���u��@�O~!� 4@P]H���!?@��,��@�w1D��ٿ���u��@�O~!� 4@P]H���!?@��,��@�䌐�ٿ������@t0MrO4@}��]��!?�˷l@��@�䌐�ٿ������@t0MrO4@}��]��!?�˷l@��@�䌐�ٿ������@t0MrO4@}��]��!?�˷l@��@�䌐�ٿ������@t0MrO4@}��]��!?�˷l@��@�䌐�ٿ������@t0MrO4@}��]��!?�˷l@��@��}�|�ٿܽ�����@q��3�4@~�6E�!?��S4;��@���ҡٿk����@L\�C�4@��x��!?�jD=��@���ҡٿk����@L\�C�4@��x��!?�jD=��@���ҡٿk����@L\�C�4@��x��!?�jD=��@���ҡٿk����@L\�C�4@��x��!?�jD=��@���S�ٿ9u�k���@&�Fv/4@E��;��!?�O�2��@���S�ٿ9u�k���@&�Fv/4@E��;��!?�O�2��@���S�ٿ9u�k���@&�Fv/4@E��;��!?�O�2��@���S�ٿ9u�k���@&�Fv/4@E��;��!?�O�2��@���S�ٿ9u�k���@&�Fv/4@E��;��!?�O�2��@��*�(�ٿ��W	���@�i	XE4@��#�~�!?�uoM<��@��M�#�ٿ���o���@W���5 4@e ���!?ӸO/��@��M�#�ٿ���o���@W���5 4@e ���!?ӸO/��@��M�#�ٿ���o���@W���5 4@e ���!?ӸO/��@�c�[�ٿ{Y���@Z�EP�3@����!?�6�"��@q�AL��ٿ�'����@b�N���3@n��mΐ!?�Ue�!��@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@8X/b`�ٿ�E,���@G޿�3@Q%����!?�Y���@I�j�ٿm��Z��@��$0��3@z��;�!?��n���@I�j�ٿm��Z��@��$0��3@z��;�!?��n���@I�j�ٿm��Z��@��$0��3@z��;�!?��n���@I�j�ٿm��Z��@��$0��3@z��;�!?��n���@	�fšٿ�)!����@�L�:4@��̐!?�#?��@	�fšٿ�)!����@�L�:4@��̐!?�#?��@	�fšٿ�)!����@�L�:4@��̐!?�#?��@	�fšٿ�)!����@�L�:4@��̐!?�#?��@	�fšٿ�)!����@�L�:4@��̐!?�#?��@	�fšٿ�)!����@�L�:4@��̐!?�#?��@!8?[�ٿt����@yN[-�4@l�#���!?
+��C��@!8?[�ٿt����@yN[-�4@l�#���!?
+��C��@!8?[�ٿt����@yN[-�4@l�#���!?
+��C��@!8?[�ٿt����@yN[-�4@l�#���!?
+��C��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@�wB)
�ٿk#X���@���R�4@<h�ǐ!?j݅�=��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@w��E1�ٿG},���@�U�3@������!?��?#��@���0�ٿ�_����@|��8�3@>4 �!?*�d�$��@���0�ٿ�_����@|��8�3@>4 �!?*�d�$��@���0�ٿ�_����@|��8�3@>4 �!?*�d�$��@�~��~�ٿ�4�m���@v��I 4@m���!?q]5K3��@�~��~�ٿ�4�m���@v��I 4@m���!?q]5K3��@�~��~�ٿ�4�m���@v��I 4@m���!?q]5K3��@�~��~�ٿ�4�m���@v��I 4@m���!?q]5K3��@�9�'��ٿõe���@�7jA�3@ѷ�b�!?pA� ��@�9�'��ٿõe���@�7jA�3@ѷ�b�!?pA� ��@�9�'��ٿõe���@�7jA�3@ѷ�b�!?pA� ��@�ch�ٿ���f��@�!�K��3@Ş�)А!?[;m�	��@�ch�ٿ���f��@�!�K��3@Ş�)А!?[;m�	��@�ch�ٿ���f��@�!�K��3@Ş�)А!?[;m�	��@L��
�ٿ.U�����@�K�d��3@��~��!?�vWJ)��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@ꊢ�V�ٿ��x���@؜�)C�3@�5��!?�I`Z��@�U�ٿ@IH��@����3@��}S��!?��h����@�U�ٿ@IH��@����3@��}S��!?��h����@�U�ٿ@IH��@����3@��}S��!?��h����@�U�ٿ@IH��@����3@��}S��!?��h����@�U�ٿ@IH��@����3@��}S��!?��h����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@�Բ
�ٿ՟�2���@<֋���3@�>�E��!?_0����@��a�Öٿ.��3��@sz?���3@�6��!?f�K����@��a�Öٿ.��3��@sz?���3@�6��!?f�K����@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@��K�7�ٿ7�p���@�-��3@����!?U�I���@�;gI}�ٿ��UD���@ PtZ��3@xSِ!?�y����@�;gI}�ٿ��UD���@ PtZ��3@xSِ!?�y����@�;gI}�ٿ��UD���@ PtZ��3@xSِ!?�y����@#*�W�ٿxt	����@�S�e��3@;�צ��!?���J���@#*�W�ٿxt	����@�S�e��3@;�צ��!?���J���@#*�W�ٿxt	����@�S�e��3@;�צ��!?���J���@#*�W�ٿxt	����@�S�e��3@;�צ��!?���J���@#*�W�ٿxt	����@�S�e��3@;�צ��!?���J���@i�C��ٿ��F� ��@��!d�3@dk*b��!?�7�a���@�y6�іٿ�;x	��@s5�9��3@o�V��!?�	Y���@�y6�іٿ�;x	��@s5�9��3@o�V��!?�	Y���@�y6�іٿ�;x	��@s5�9��3@o�V��!?�	Y���@�g�-�ٿ����@����3@��zݐ!?������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@�V��ٿa���@��j���3@%z(Ր!?�������@+�֣��ٿө~`��@�	G1�3@��ؐ!?�~@`���@+�֣��ٿө~`��@�	G1�3@��ؐ!?�~@`���@+�֣��ٿө~`��@�	G1�3@��ؐ!?�~@`���@�gr�ٿ? ����@+ϲI��3@�xL�!?������@�gr�ٿ? ����@+ϲI��3@�xL�!?������@0F�g��ٿl@���@�����3@dnp��!?pIW����@0F�g��ٿl@���@�����3@dnp��!?pIW����@0F�g��ٿl@���@�����3@dnp��!?pIW����@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@���k3�ٿR�x���@����Q�3@�K��!?���J���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@	���ٿ�C�-���@U��(�3@�}���!?�װA���@DO�Ǡٿ��r����@3��<��3@_ٻx�!?�{t���@DO�Ǡٿ��r����@3��<��3@_ٻx�!?�{t���@DO�Ǡٿ��r����@3��<��3@_ٻx�!?�{t���@DO�Ǡٿ��r����@3��<��3@_ٻx�!?�{t���@��_��ٿ�J�����@�����3@� NW��!?5GX���@��_��ٿ�J�����@�����3@� NW��!?5GX���@����֞ٿn�Z~ ��@?W����3@�	m��!?�Y�l���@����֞ٿn�Z~ ��@?W����3@�	m��!?�Y�l���@����֞ٿn�Z~ ��@?W����3@�	m��!?�Y�l���@����֞ٿn�Z~ ��@?W����3@�	m��!?�Y�l���@[v 6�ٿ_�.� ��@�rV+y�3@'�^���!?���Y���@[v 6�ٿ_�.� ��@�rV+y�3@'�^���!?���Y���@�oS��ٿ�=L��@������3@G戏�!?�7�o���@�oS��ٿ�=L��@������3@G戏�!?�7�o���@�oS��ٿ�=L��@������3@G戏�!?�7�o���@�oS��ٿ�=L��@������3@G戏�!?�7�o���@�oS��ٿ�=L��@������3@G戏�!?�7�o���@Ŧ��M�ٿ�e�S���@����3@��!?������@ON����ٿ�]FC���@<�����3@�Ĩݳ�!?N�����@ON����ٿ�]FC���@<�����3@�Ĩݳ�!?N�����@��[���ٿ9� ����@�\���3@"1!���!?���	���@��[���ٿ9� ����@�\���3@"1!���!?���	���@��[���ٿ9� ����@�\���3@"1!���!?���	���@ùFl�ٿ�� ����@Ϧ^��3@|a!��!?Ԯ����@ùFl�ٿ�� ����@Ϧ^��3@|a!��!?Ԯ����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@�m_*�ٿ�p�����@�Ҥ[G�3@�ˣ~�!?�1F����@;v�KD�ٿ�����@5�9��3@`���!?Ud�D��@FfОٿc*����@7:�Ě�3@1G+��!?D����@FfОٿc*����@7:�Ě�3@1G+��!?D����@FfОٿc*����@7:�Ě�3@1G+��!?D����@FfОٿc*����@7:�Ě�3@1G+��!?D����@FfОٿc*����@7:�Ě�3@1G+��!?D����@s�B2��ٿ�8���@~��c�3@�{�A��!?sA�l���@>MO�
�ٿp�.���@�����3@暸�!?�	xq���@c��ٿ\%&����@���3@���Y��!?������@ҭ�P@�ٿ~�j����@�wO!x�3@DZ5��!?	������@ҭ�P@�ٿ~�j����@�wO!x�3@DZ5��!?	������@sWl��ٿ"���@�'���3@:G�jv�!?B������@sWl��ٿ"���@�'���3@:G�jv�!?B������@sWl��ٿ"���@�'���3@:G�jv�!?B������@S�M�ٿ��@r ��@�P�kF�3@ǰ��!?�>�&���@S�M�ٿ��@r ��@�P�kF�3@ǰ��!?�>�&���@S�M�ٿ��@r ��@�P�kF�3@ǰ��!?�>�&���@S�M�ٿ��@r ��@�P�kF�3@ǰ��!?�>�&���@S�M�ٿ��@r ��@�P�kF�3@ǰ��!?�>�&���@��ٿ�.�n���@�����3@��+�!?]����@��ٿ�.�n���@�����3@��+�!?]����@��ٿ�.�n���@�����3@��+�!?]����@�=���ٿ��S��@g�	o��3@,��k�!?X��@�=���ٿ��S��@g�	o��3@,��k�!?X��@�=���ٿ��S��@g�	o��3@,��k�!?X��@�=���ٿ��S��@g�	o��3@,��k�!?X��@�=���ٿ��S��@g�	o��3@,��k�!?X��@*�I�ٿJ3;n���@�=�Y��3@��zߐ!?��Y/��@*�I�ٿJ3;n���@�=�Y��3@��zߐ!?��Y/��@*�I�ٿJ3;n���@�=�Y��3@��zߐ!?��Y/��@*�I�ٿJ3;n���@�=�Y��3@��zߐ!?��Y/��@*�I�ٿJ3;n���@�=�Y��3@��zߐ!?��Y/��@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@R؀��ٿ������@�7����3@�C��!?4��^���@���i1�ٿ�@U����@���M\�3@Ú��!??����@���i1�ٿ�@U����@���M\�3@Ú��!??����@���i1�ٿ�@U����@���M\�3@Ú��!??����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@�0m�t�ٿ-:e���@u���3@ẇdr�!?�8�����@.�U<�ٿ;�׌���@C���I�3@�h����!?�gر;��@.�U<�ٿ;�׌���@C���I�3@�h����!?�gر;��@.�U<�ٿ;�׌���@C���I�3@�h����!?�gر;��@.�U<�ٿ;�׌���@C���I�3@�h����!?�gر;��@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@��V>Υٿ�3 "��@�Gzb�3@�9N��!?j�M���@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@MB��y�ٿ'�! ��@�J�R��3@ܽ9��!?������@i�C{d�ٿ�����@��'���3@o�\)�!?��+���@i�C{d�ٿ�����@��'���3@o�\)�!?��+���@i�C{d�ٿ�����@��'���3@o�\)�!?��+���@�]Յ��ٿ7.���@�o?��3@��!�ѐ!?�z�L���@�]Յ��ٿ7.���@�o?��3@��!�ѐ!?�z�L���@Uw��ٿ]z���@_rk��3@��݈��!?8�F�q��@Uw��ٿ]z���@_rk��3@��݈��!?8�F�q��@Uw��ٿ]z���@_rk��3@��݈��!?8�F�q��@Uw��ٿ]z���@_rk��3@��݈��!?8�F�q��@=���0�ٿs�]����@
=���3@l)�M�!?S�����@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@r}�[L�ٿ�Y5N���@!��i��3@k<��Ő!?��m ���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@��W=�ٿ �����@���E�3@D�h�!?�0>���@�~̘�ٿRq�5��@�?�D�3@}��X��!?�K}�L��@�~̘�ٿRq�5��@�?�D�3@}��X��!?�K}�L��@�~̘�ٿRq�5��@�?�D�3@}��X��!?�K}�L��@�~̘�ٿRq�5��@�?�D�3@}��X��!?�K}�L��@H�%�ͥٿ�p����@��d���3@�QBh��!?�|�r��@H�%�ͥٿ�p����@��d���3@�QBh��!?�|�r��@H�%�ͥٿ�p����@��d���3@�QBh��!?�|�r��@H�%�ͥٿ�p����@��d���3@�QBh��!?�|�r��@H�%�ͥٿ�p����@��d���3@�QBh��!?�|�r��@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@�&iN��ٿ�O�6���@�+R���3@v9����!?!����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@s�k��ٿ�����@���1p�3@�ɠ���!?O�5����@|�!h�ٿ��bG���@��l��3@�����!?N�"����@|�!h�ٿ��bG���@��l��3@�����!?N�"����@0Js��ٿ�����@j?e���3@�H��!?�XH����@0Js��ٿ�����@j?e���3@�H��!?�XH����@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@�4w���ٿ��ܿ��@�΄�I�3@|X�N��!?�j�f��@��>�ٿ�99��@��G`]�3@&�!?أ'����@��>�ٿ�99��@��G`]�3@&�!?أ'����@R�{"J�ٿr�S���@Uʞ+��3@����!?z�����@R�{"J�ٿr�S���@Uʞ+��3@����!?z�����@~F#A�ٿ�d!����@�'����3@U2��!?9���@~F#A�ٿ�d!����@�'����3@U2��!?9���@�I��ؠٿY��� ��@w��*�3@��!�Ɛ!?U�L�q��@�I��ؠٿY��� ��@w��*�3@��!�Ɛ!?U�L�q��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@��/~�ٿ �~���@��~�c�3@t�7}��!?δ�K��@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@>r�m�ٿW�Ȥ��@�����3@
d����!?\@W���@����ٿp�����@�>7�3@�Γ��!?w*.���@����ٿp�����@�>7�3@�Γ��!?w*.���@����ٿp�����@�>7�3@�Γ��!?w*.���@\�>Ϙ�ٿ�hn�.��@��|i�3@��.���!?�Ɍ��@\�>Ϙ�ٿ�hn�.��@��|i�3@��.���!?�Ɍ��@\�>Ϙ�ٿ�hn�.��@��|i�3@��.���!?�Ɍ��@\�>Ϙ�ٿ�hn�.��@��|i�3@��.���!?�Ɍ��@=��힘ٿz�
T��@��
���3@�3F_��!?�|K����@=��힘ٿz�
T��@��
���3@�3F_��!?�|K����@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@���?��ٿ;W1�B��@��}*�3@ t��_�!?���H*��@�A#%�ٿN���$��@X�q=��3@�ºY��!?H޹;��@�A#%�ٿN���$��@X�q=��3@�ºY��!?H޹;��@�A#%�ٿN���$��@X�q=��3@�ºY��!?H޹;��@�A#%�ٿN���$��@X�q=��3@�ºY��!?H޹;��@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@zZ���ٿ�ąX*��@r�5��3@��5��!?�����@ \���ٿC�ʵF��@4d��3@9sJː!?Z�uܧ��@ \���ٿC�ʵF��@4d��3@9sJː!?Z�uܧ��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�"��V�ٿ y�g��@Lvo���3@��RU��!?F�4NT��@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�{�M��ٿy{����@ca����3@բ�Ƿ�!?y,T2���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@�H�5�ٿJ�J��@�6��3@�&.�!?�	dL���@��J.�ٿm�����@΢����3@l�ɕ�!?������@��J.�ٿm�����@΢����3@l�ɕ�!?������@��J.�ٿm�����@΢����3@l�ɕ�!?������@��J.�ٿm�����@΢����3@l�ɕ�!?������@��LN�ٿ��m��@�(�a�3@i� 5��!?eҔ�s��@��LN�ٿ��m��@�(�a�3@i� 5��!?eҔ�s��@��LN�ٿ��m��@�(�a�3@i� 5��!?eҔ�s��@��LN�ٿ��m��@�(�a�3@i� 5��!?eҔ�s��@�m����ٿ鮄pB��@�F�G�3@&���!?E�����@�m����ٿ鮄pB��@�F�G�3@&���!?E�����@�m����ٿ鮄pB��@�F�G�3@&���!?E�����@�m����ٿ鮄pB��@�F�G�3@&���!?E�����@�����ٿ��x�O��@��ӟz�3@3��!?؂m��@�����ٿ��x�O��@��ӟz�3@3��!?؂m��@�����ٿ��x�O��@��ӟz�3@3��!?؂m��@�����ٿ��x�O��@��ӟz�3@3��!?؂m��@/�yKQ�ٿ��W��@�3���3@�W�ې!?=��K��@/�yKQ�ٿ��W��@�3���3@�W�ې!?=��K��@/�yKQ�ٿ��W��@�3���3@�W�ې!?=��K��@�RW��ٿ�?�m��@����3@]���i�!?���c���@�RW��ٿ�?�m��@����3@]���i�!?���c���@�RW��ٿ�?�m��@����3@]���i�!?���c���@�RW��ٿ�?�m��@����3@]���i�!?���c���@�RW��ٿ�?�m��@����3@]���i�!?���c���@�RW��ٿ�?�m��@����3@]���i�!?���c���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@j�&K�ٿ���(��@��w�}�3@��-���!?�6B^���@6���D�ٿ�����@N�o@�3@��:7��!?г8/���@6���D�ٿ�����@N�o@�3@��:7��!?г8/���@�Yޱf�ٿi��S���@�iJ���3@#�F��!?�X��a��@�Yޱf�ٿi��S���@�iJ���3@#�F��!?�X��a��@�Yޱf�ٿi��S���@�iJ���3@#�F��!?�X��a��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@��-�ٿ��u�և�@���>�3@6G��!?���E��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@ﯗ�Ҟٿ~7�*��@5�<1��3@܂>ߐ!?��LG��@+�|�G�ٿ2����@���R�3@��4̐!?!Oڗ���@+�|�G�ٿ2����@���R�3@��4̐!?!Oڗ���@+�|�G�ٿ2����@���R�3@��4̐!?!Oڗ���@+�|�G�ٿ2����@���R�3@��4̐!?!Oڗ���@+�|�G�ٿ2����@���R�3@��4̐!?!Oڗ���@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@ʴ*��ٿ������@h+���3@N�(�ؐ!?y�6�|��@�!�n�ٿd�v·�@[Kʘ�3@���Ս�!?���U��@o��'��ٿ�a���@�C���3@ߠ!q��!?Ȳ�w>��@o��'��ٿ�a���@�C���3@ߠ!q��!?Ȳ�w>��@o��'��ٿ�a���@�C���3@ߠ!q��!?Ȳ�w>��@o��'��ٿ�a���@�C���3@ߠ!q��!?Ȳ�w>��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@� �PU�ٿ�>����@����#�3@��%4��!?,�HE��@0�NH�ٿ���$&��@�p6��3@������!?�.Db���@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�8'��ٿ�l�N4��@1;&�3�3@�Ő!?��}��@�y�ڗٿJ����@��ux�3@�W=��!?H������@�y�ڗٿJ����@��ux�3@�W=��!?H������@�M7ّ�ٿ꫙���@v�K�5�3@C�y-ې!?Z�
"��@uMu�ٿ`i��ć�@RW�ye�3@O�ʐ!?��T^��@uMu�ٿ`i��ć�@RW�ye�3@O�ʐ!?��T^��@uMu�ٿ`i��ć�@RW�ye�3@O�ʐ!?��T^��@1	���ٿn�K·�@{t� �3@�zH���!?O����@1	���ٿn�K·�@{t� �3@�zH���!?O����@iǽ�-�ٿ��
3��@��*��3@}�|"�!?.�zM��@�m�G�ٿ�h���@�!��3@9��Tc�!?�l���@�m�G�ٿ�h���@�!��3@9��Tc�!?�l���@�m�G�ٿ�h���@�!��3@9��Tc�!?�l���@���2p�ٿ�B.A���@�W�{�3@Φ��Ő!?}f�r ��@���2p�ٿ�B.A���@�W�{�3@Φ��Ő!?}f�r ��@���2p�ٿ�B.A���@�W�{�3@Φ��Ő!?}f�r ��@�U���ٿV|I&V��@� A�)�3@����!?6z?�y��@�y�\7�ٿh3��·�@����y�3@נϐ!?���p��@�y�\7�ٿh3��·�@����y�3@נϐ!?���p��@%;��.�ٿ�@�['��@G8����3@'��ڐ!??�*ӣ��@�4��ٿ
�c��@��2p�3@IH@s�!?l�bx��@�e���ٿ���w��@0����3@���Ð!?��W���@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@ �@���ٿ[��L��@�h�*��3@k
�ϐ!?ˍ$����@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@��N��ٿ�*´���@Q�*��3@�X뮐!?�k�ey�@WG���ٿ֫uwx��@��Y��3@����!? ���� �@������ٿ��6u��@W���P�3@r~� �!?>%�{F��@������ٿ��6u��@W���P�3@r~� �!?>%�{F��@������ٿ��6u��@W���P�3@r~� �!?>%�{F��@������ٿ��6u��@W���P�3@r~� �!?>%�{F��@������ٿ��6u��@W���P�3@r~� �!?>%�{F��@ު�ؒ�ٿ��R7(��@)��M��3@�})㮐!?������@ު�ؒ�ٿ��R7(��@)��M��3@�})㮐!?������@��{�ٿ�bZ߆�@�c��O�3@48擐!?��hy���@��{�ٿ�bZ߆�@�c��O�3@48擐!?��hy���@��{�ٿ�bZ߆�@�c��O�3@48擐!?��hy���@��{�ٿ�bZ߆�@�c��O�3@48擐!?��hy���@+�w���ٿ@ޑ{��@��dw�3@'�q�!?�iL���@+�w���ٿ@ޑ{��@��dw�3@'�q�!?�iL���@���1�ٿ���kh��@���e��3@f+��!?2f_��@���1�ٿ���kh��@���e��3@f+��!?2f_��@���1�ٿ���kh��@���e��3@f+��!?2f_��@���1�ٿ���kh��@���e��3@f+��!?2f_��@�7�k
�ٿ� °��@(����3@���!?��Qw��@�7�k
�ٿ� °��@(����3@���!?��Qw��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@�w�<�ٿ������@�|�d�3@�|�!?-eA��@���/��ٿ�y��G��@.�J���3@޷��|�!?�����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@��k�ٿʐ�Z���@�����3@<�oː!?��h����@�b\uڜٿl�D���@ل;���3@U�	�Ɛ!?6��r���@�	�-F�ٿJ6_����@;�K�&�3@�[����!?����@�	�-F�ٿJ6_����@;�K�&�3@�[����!?����@�	�-F�ٿJ6_����@;�K�&�3@�[����!?����@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�蹰]�ٿs��lQ��@2�M�3�3@<��R�!?_u���@�t�ϡٿ�2HՂ��@ĕ.���3@f"���!?��)�l��@�t�ϡٿ�2HՂ��@ĕ.���3@f"���!?��)�l��@�t�ϡٿ�2HՂ��@ĕ.���3@f"���!?��)�l��@�t�ϡٿ�2HՂ��@ĕ.���3@f"���!?��)�l��@�t�ϡٿ�2HՂ��@ĕ.���3@f"���!?��)�l��@�Gk��ٿ��pp��@�J���3@�1+��!?J@��̣�@�Gk��ٿ��pp��@�J���3@�1+��!?J@��̣�@$�#���ٿ|���n��@�''�3@F�����!?�Jo ��@$�#���ٿ|���n��@�''�3@F�����!?�Jo ��@$�#���ٿ|���n��@�''�3@F�����!?�Jo ��@$�#���ٿ|���n��@�''�3@F�����!?�Jo ��@$�#���ٿ|���n��@�''�3@F�����!?�Jo ��@a�t,�ٿ{��S�@nޣR��3@�MА!?��sM�s�@a�t,�ٿ{��S�@nޣR��3@�MА!?��sM�s�@a�t,�ٿ{��S�@nޣR��3@�MА!?��sM�s�@a�t,�ٿ{��S�@nޣR��3@�MА!?��sM�s�@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@ Oꥸ�ٿ@X�ǀ�@�A/�F�3@�R�n��!?��7rP��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@2�^��ٿ�)|?dt�@&g��3@a=�ߐ!?��w ��@�S%l��ٿ<O���s�@d��!��3@G����!?Fc��@�S%l��ٿ<O���s�@d��!��3@G����!?Fc��@o�lm�ٿ�?P�Xh�@y�u��3@�Ԧ���!?9ݵa�@o�lm�ٿ�?P�Xh�@y�u��3@�Ԧ���!?9ݵa�@o�lm�ٿ�?P�Xh�@y�u��3@�Ԧ���!?9ݵa�@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@�x)�ٿ8�A�Cu�@t'c���3@5�򺷐!?�9����@G�t啨ٿRI�@o�@9��>�3@)�!?V����@G�t啨ٿRI�@o�@9��>�3@)�!?V����@G�t啨ٿRI�@o�@9��>�3@)�!?V����@G�t啨ٿRI�@o�@9��>�3@)�!?V����@G�t啨ٿRI�@o�@9��>�3@)�!?V����@�)m�ԡٿ��٩Es�@�|���3@�S,�!?=1ܸ�@�)m�ԡٿ��٩Es�@�|���3@�S,�!?=1ܸ�@�)m�ԡٿ��٩Es�@�|���3@�S,�!?=1ܸ�@�)m�ԡٿ��٩Es�@�|���3@�S,�!?=1ܸ�@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@
�&�k�ٿM�3?r�@�}�(�3@x�u�ܐ!?r�^���@�<����ٿ��cdg�@N�-(�3@����֐!?����@�<����ٿ��cdg�@N�-(�3@����֐!?����@�<����ٿ��cdg�@N�-(�3@����֐!?����@�<����ٿ��cdg�@N�-(�3@����֐!?����@�<����ٿ��cdg�@N�-(�3@����֐!?����@�<����ٿ��cdg�@N�-(�3@����֐!?����@�'���ٿ��X�s�@5�P�j�3@���Ɛ!?��X_��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@9�W�ٿ�X�ka�@���3@�-���!?��	��@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@~^R}Оٿ�Q`g�@=�[��3@�ͥlא!?�L���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@�fv��ٿ;P �`�@��%�J�3@�w� Ð!?Jm.3���@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@���:ȣٿf�f_�@��oļ�3@Қ�)ݐ!?0���2}�@�	�
��ٿ�ꦜ�d�@�U��3@�
���!?�K� ���@�-Ʌ�ٿ�5�zxu�@��v�3@��ͼ��!?�6>���@�-Ʌ�ٿ�5�zxu�@��v�3@��ͼ��!?�6>���@�-Ʌ�ٿ�5�zxu�@��v�3@��ͼ��!?�6>���@�-Ʌ�ٿ�5�zxu�@��v�3@��ͼ��!?�6>���@Y���ٿ��Fn�@�VP	�3@z(	G��!?׌Yc�@Y���ٿ��Fn�@�VP	�3@z(	G��!?׌Yc�@Y���ٿ��Fn�@�VP	�3@z(	G��!?׌Yc�@Y���ٿ��Fn�@�VP	�3@z(	G��!?׌Yc�@���AP�ٿ0�\?n�@��� '�3@dO����!?S���8j�@���AP�ٿ0�\?n�@��� '�3@dO����!?S���8j�@���AP�ٿ0�\?n�@��� '�3@dO����!?S���8j�@���AP�ٿ0�\?n�@��� '�3@dO����!?S���8j�@���AP�ٿ0�\?n�@��� '�3@dO����!?S���8j�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@!v��؜ٿ��;�Dl�@z��Rl�3@*�K�Đ!?���_F�@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@���qo�ٿ�s{�a�@ۧ�1�3@��!?�������@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@<qR�Ʀٿe�B�p�@���Ӯ�3@����!?Q4��@\_rA�ٿ(|�:�_�@PM����3@E��!?C6	G��@\_rA�ٿ(|�:�_�@PM����3@E��!?C6	G��@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@����ٿ�\U6k�@���b��3@s��)��!?�i��8�@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�T���ٿ���f�@yƙ��3@ELIT��!?��1��@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@�Ca�ٿ߾sT�g�@��;��3@q\����!?�����@q:�N�ٿ�m�Wim�@�h�+��3@�4orȐ!?�$"]?�@q:�N�ٿ�m�Wim�@�h�+��3@�4orȐ!?�$"]?�@q:�N�ٿ�m�Wim�@�h�+��3@�4orȐ!?�$"]?�@q:�N�ٿ�m�Wim�@�h�+��3@�4orȐ!?�$"]?�@q:�N�ٿ�m�Wim�@�h�+��3@�4orȐ!?�$"]?�@��q�ܝٿ�� eg�@~��2�3@�W�K��!?�/�L��@��q�ܝٿ�� eg�@~��2�3@�W�K��!?�/�L��@��q�ܝٿ�� eg�@~��2�3@�W�K��!?�/�L��@��q�ܝٿ�� eg�@~��2�3@�W�K��!?�/�L��@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@\1����ٿ]=��p�@�o�7�3@\B�5��!?jٳ��j�@3%�y�ٿ� Q�e�@1�*K��3@�e����!?C�F�ݱ�@3%�y�ٿ� Q�e�@1�*K��3@�e����!?C�F�ݱ�@3%�y�ٿ� Q�e�@1�*K��3@�e����!?C�F�ݱ�@�����ٿ��/h�@uZZ"�3@�C��!?��%���@�����ٿ��/h�@uZZ"�3@�C��!?��%���@�����ٿ��/h�@uZZ"�3@�C��!?��%���@�����ٿ��/h�@uZZ"�3@�C��!?��%���@�����ٿ��/h�@uZZ"�3@�C��!?��%���@�����ٿ��/h�@uZZ"�3@�C��!?��%���@_�H爝ٿ��ՄJd�@�n>�3@::���!?�Do\���@�j叡�ٿ3��sa�@ö}���3@�Vڈ�!?^��`�@�j叡�ٿ3��sa�@ö}���3@�Vڈ�!?^��`�@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@ի_՜ٿg�-�j�@���\��3@��!?e��|��@����ٿ��3��b�@A��3��3@��B���!?�� �w��@����ٿ��3��b�@A��3��3@��B���!?�� �w��@� ��d�ٿ�O�{�l�@a���3@`IR��!?|א��1�@� ��d�ٿ�O�{�l�@a���3@`IR��!?|א��1�@� ��d�ٿ�O�{�l�@a���3@`IR��!?|א��1�@� ��d�ٿ�O�{�l�@a���3@`IR��!?|א��1�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@@~���ٿ*���[�@��%�3@�N<!?ƒ{��V�@8�9#��ٿ�y���o�@瀼���3@��0��!?X�^pT��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@6�܌�ٿ�Ƽ�q�@b%��Y�3@��p�!?qCcv��@ӻϽM�ٿD�f�@eT�m�3@�i�6��!?~��v7�@C}A���ٿ͝��c�@Q�fB�3@I�����!?�i��M�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@f�W���ٿ�p��v�@�K!�3@�����!?��1�O�@nL�٦ٿ7ɇ�Ko�@%-�3@=�ѱ�!?&��Z���@<g2<«ٿa���t�@5�_��3@3F�ސ!?h�����@<g2<«ٿa���t�@5�_��3@3F�ސ!?h�����@<g2<«ٿa���t�@5�_��3@3F�ސ!?h�����@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@��&��ٿDq�Y-o�@���B8�3@OlӐ!?���x;��@�R�7�ٿR:g�t�@�Mb}��3@Ui�M��!?�	����@�R�7�ٿR:g�t�@�Mb}��3@Ui�M��!?�	����@�R�7�ٿR:g�t�@�Mb}��3@Ui�M��!?�	����@�R�7�ٿR:g�t�@�Mb}��3@Ui�M��!?�	����@��P���ٿ��6g�@hQx5�3@q���!?$�h�y�@���r��ٿP�U�n�@��_�N�3@A��!?x���@���r��ٿP�U�n�@��_�N�3@A��!?x���@���t�ٿ3�e�m�@+$Z̫�3@|�mԐ!?�������@����ѥٿ��;�qo�@��B0�3@8`�|��!?2lV����@����ѥٿ��;�qo�@��B0�3@8`�|��!?2lV����@����ѥٿ��;�qo�@��B0�3@8`�|��!?2lV����@����ѥٿ��;�qo�@��B0�3@8`�|��!?2lV����@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@I,���ٿ����s�@,���3@�-�!?KU7G��@uŽ�D�ٿQ���m�@�Zy��3@��ʥ�!? �3�@uŽ�D�ٿQ���m�@�Zy��3@��ʥ�!? �3�@uŽ�D�ٿQ���m�@�Zy��3@��ʥ�!? �3�@��&H��ٿ�Cг(l�@U���i�3@O���ܐ!?�L崏�@��&H��ٿ�Cг(l�@U���i�3@O���ܐ!?�L崏�@��&H��ٿ�Cг(l�@U���i�3@O���ܐ!?�L崏�@��&H��ٿ�Cг(l�@U���i�3@O���ܐ!?�L崏�@��&H��ٿ�Cг(l�@U���i�3@O���ܐ!?�L崏�@���֞ٿ�>Z�zn�@{1��3@���Ő!?�P(�u�@���֞ٿ�>Z�zn�@{1��3@���Ő!?�P(�u�@�t���ٿ�
n�@ 5�Ԑ�3@�g;/��!??�����@�t���ٿ�
n�@ 5�Ԑ�3@�g;/��!??�����@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@'oӆ��ٿ7Vh,�l�@6m/�3@'���!?�TY�+��@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@ j�}��ٿHU\L�u�@�����3@��͒̐!?V��&`k�@���6��ٿ��rg�r�@�����3@|0�!?%��*��@���6��ٿ��rg�r�@�����3@|0�!?%��*��@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@k9��#�ٿ1��y�@?O�9o�3@垁j��!?���E�@�!؈u�ٿ��{b�@)�P"�3@𥨗��!?=�����@�!؈u�ٿ��{b�@)�P"�3@𥨗��!?=�����@�!؈u�ٿ��{b�@)�P"�3@𥨗��!?=�����@�!؈u�ٿ��{b�@)�P"�3@𥨗��!?=�����@�,�.��ٿ.��\�@��#��3@\��B��!?�^�Z{ �@g���~�ٿl��bq�@:l���3@����!?���%<�@���˕ٿ���Lr�@=i<R|�3@�i�5��!?C�����@���˕ٿ���Lr�@=i<R|�3@�i�5��!?C�����@���˕ٿ���Lr�@=i<R|�3@�i�5��!?C�����@���˕ٿ���Lr�@=i<R|�3@�i�5��!?C�����@���˕ٿ���Lr�@=i<R|�3@�i�5��!?C�����@=��qL�ٿ�����s�@����3@[�߅��!?�5	�|n�@=��qL�ٿ�����s�@����3@[�߅��!?�5	�|n�@�i�a�ٿh����v�@�f����3@���8i�!?�6����@�i�a�ٿh����v�@�f����3@���8i�!?�6����@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@���Ȧٿ��υ���@Y���3@�|�O|�!?KZ���@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@f�m�<�ٿW��@��@ ��ِ�3@{kS�{�!?��)IJ��@�_��V�ٿ���<�~�@���4�3@�'�o��!?�Ai���@�_��V�ٿ���<�~�@���4�3@�'�o��!?�Ai���@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@E��B�ٿlm���]�@Y���3@t�&8ː!?[Bn��L�@�j��Q�ٿ8��>Nz�@X� c�3@��6�ΐ!?8� �L`�@2B��ٿ)�Ǎ�@�t�Ub�3@X�=l�!?��1*wj�@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@&��8�ٿ-hѳ��@�����3@Y�thې!?t��/*��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@�m���ٿ���1p�@=^V��3@V��^��!?K�+١��@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@���+"�ٿ��l�@O����3@#1�7ڐ!?:R3PK�@��-��ٿK^�Rx�@�b#��3@̛�P�!?��.�-O�@�UB�
�ٿ pD�܌�@�Aڗ��3@+���!?8j���@~���ٿk�����@|>�8��3@3]�»�!?�%_ʔ��@~���ٿk�����@|>�8��3@3]�»�!?�%_ʔ��@~���ٿk�����@|>�8��3@3]�»�!?�%_ʔ��@~���ٿk�����@|>�8��3@3]�»�!?�%_ʔ��@t_A�Кٿ���x!��@�b�h�3@��ܐ!?w��q���@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@�Dx���ٿ�*����@���й�3@�S��!?�}v/��@���T-�ٿ`�0�/��@2��F �3@�R�=�!?�\���$�@���T-�ٿ`�0�/��@2��F �3@�R�=�!?�\���$�@���T-�ٿ`�0�/��@2��F �3@�R�=�!?�\���$�@���T-�ٿ`�0�/��@2��F �3@�R�=�!?�\���$�@���T-�ٿ`�0�/��@2��F �3@�R�=�!?�\���$�@�mp���ٿ��6�o}�@�yMI��3@��Ҿ�!?8�i-"�@�mp���ٿ��6�o}�@�yMI��3@��Ҿ�!?8�i-"�@�mp���ٿ��6�o}�@�yMI��3@��Ҿ�!?8�i-"�@���J��ٿ��VC>u�@v���3@Á����!?C�#�G�@���J��ٿ��VC>u�@v���3@Á����!?C�#�G�@���J��ٿ��VC>u�@v���3@Á����!?C�#�G�@���J��ٿ��VC>u�@v���3@Á����!?C�#�G�@�F�ɤٿ�1Ⅶ�@x��UR�3@��A�!?�y�!:e�@�F�ɤٿ�1Ⅶ�@x��UR�3@��A�!?�y�!:e�@�F�ɤٿ�1Ⅶ�@x��UR�3@��A�!?�y�!:e�@�F�ɤٿ�1Ⅶ�@x��UR�3@��A�!?�y�!:e�@���,Q�ٿQ�VP��@p�3���3@�*��͐!?2�B�x��@���,Q�ٿQ�VP��@p�3���3@�*��͐!?2�B�x��@���,Q�ٿQ�VP��@p�3���3@�*��͐!?2�B�x��@���,Q�ٿQ�VP��@p�3���3@�*��͐!?2�B�x��@���,Q�ٿQ�VP��@p�3���3@�*��͐!?2�B�x��@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@�4>��ٿ٫�����@0 f�;�3@���!?��Yk�@;WI�ߟٿo�L@�@�����3@��-�!?C���@;WI�ߟٿo�L@�@�����3@��-�!?C���@;WI�ߟٿo�L@�@�����3@��-�!?C���@;WI�ߟٿo�L@�@�����3@��-�!?C���@@��ٿq۰d �@���d�3@paT�!? �KG�>�@@��ٿq۰d �@���d�3@paT�!? �KG�>�@@��ٿq۰d �@���d�3@paT�!? �KG�>�@@��ٿq۰d �@���d�3@paT�!? �KG�>�@@��ٿq۰d �@���d�3@paT�!? �KG�>�@��6�#�ٿ��3��@/���3@��1��!?�HtT>,�@��6�#�ٿ��3��@/���3@��1��!?�HtT>,�@%T����ٿ�ԇ����@ |��3@r����!?)�m��@%T����ٿ�ԇ����@ |��3@r����!?)�m��@%T����ٿ�ԇ����@ |��3@r����!?)�m��@R�dA�ٿo\ϼ��@<���I�3@>Q�!?�䒞d�@R�dA�ٿo\ϼ��@<���I�3@>Q�!?�䒞d�@R�dA�ٿo\ϼ��@<���I�3@>Q�!?�䒞d�@Z�{��ٿ ��4��@�|����3@�:9�!?}�(>��@Z�{��ٿ ��4��@�|����3@�:9�!?}�(>��@Z�{��ٿ ��4��@�|����3@�:9�!?}�(>��@Z�{��ٿ ��4��@�|����3@�:9�!?}�(>��@Z�{��ٿ ��4��@�|����3@�:9�!?}�(>��@�摳s�ٿ�*m�<A�@�h����3@ڹ��ѐ!?q*�"�@*��K�ٿ�"��mR�@�_]�d�3@뭻��!?f������@*��K�ٿ�"��mR�@�_]�d�3@뭻��!?f������@*��K�ٿ�"��mR�@�_]�d�3@뭻��!?f������@*��K�ٿ�"��mR�@�_]�d�3@뭻��!?f������@�ilu�ٿ
��_��@[��Y��3@]���א!?�-���d�@�ilu�ٿ
��_��@[��Y��3@]���א!?�-���d�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@�<g�t�ٿ\��:I�@��"��3@��Dؐ!?b��^Ҹ�@����ٿ��%*
��@ʋ��q�3@(M��r�!?Qku~8�@����ٿ��%*
��@ʋ��q�3@(M��r�!?Qku~8�@����ٿ��%*
��@ʋ��q�3@(M��r�!?Qku~8�@#*W ��ٿ��|�C�@����3@pk�!?��Y;��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@��6�ٿ)m�=��@Υg��3@%��!?kF]��@ˡ���ٿ������@�Z����3@@JV*�!?�3��.�@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@t��G�ٿ;Y"�@�ϛ�W�3@��`� �!?r�M(��@�!;��ٿH���J��@o�B��3@4�f!?B!е��@�!;��ٿH���J��@o�B��3@4�f!?B!е��@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@2m⠚ٿ�u��)�@��.��3@�v2&�!?�m����@��-ʹ�ٿ&2�|��@�{U���3@čDw3�!?�6� ��@��-ʹ�ٿ&2�|��@�{U���3@čDw3�!?�6� ��@��-ʹ�ٿ&2�|��@�{U���3@čDw3�!?�6� ��@��-ʹ�ٿ&2�|��@�{U���3@čDw3�!?�6� ��@aV&n�ٿ6Y澁��@1DPi��3@ǦN��!?4��Bpo�@aV&n�ٿ6Y澁��@1DPi��3@ǦN��!?4��Bpo�@��O`�ٿ^y���#�@��e�+�3@�^���!?4���-�@��O`�ٿ^y���#�@��e�+�3@�^���!?4���-�@��O`�ٿ^y���#�@��e�+�3@�^���!?4���-�@$S�S_�ٿ�8�����@^�G��3@ �����!?ҙ��M��@$S�S_�ٿ�8�����@^�G��3@ �����!?ҙ��M��@$S�S_�ٿ�8�����@^�G��3@ �����!?ҙ��M��@�z_u��ٿ��aqȬ�@(�D$v�3@*H����!?���Kl��@�z_u��ٿ��aqȬ�@(�D$v�3@*H����!?���Kl��@�z_u��ٿ��aqȬ�@(�D$v�3@*H����!?���Kl��@�z_u��ٿ��aqȬ�@(�D$v�3@*H����!?���Kl��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@���ٿ=-U��@,�.��3@�Mg�!?�HZ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@����~�ٿ�=��}��@q���:�3@��8Ӑ!?y��ͧ��@�N]m�ٿ�ǂ��@x���L�3@w82��!?��qi�@�N]m�ٿ�ǂ��@x���L�3@w82��!?��qi�@�N]m�ٿ�ǂ��@x���L�3@w82��!?��qi�@�*Ԡٿ�Js���@�
l\>�3@^���ݐ!?���%��@�*Ԡٿ�Js���@�
l\>�3@^���ݐ!?���%��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@�aah�ٿ���h�@�'G�s�3@����!?�h�s|��@9�S�ٿ��$ݾ��@�I�/��3@�#�h��!?�J����@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@��N���ٿj	��nA�@1F��3@��̼�!?㢀k�Y�@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@�iA
:�ٿЩp����@]�Ҹ<�3@�ɸr�!?I$N)���@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@����ڦٿڛ�QL^�@��C��3@��3,�!?P}>�'�@�
���ٿ�[�* 8�@m�T3��3@��(��!?�7��Q�@�
���ٿ�[�* 8�@m�T3��3@��(��!?�7��Q�@�
���ٿ�[�* 8�@m�T3��3@��(��!?�7��Q�@�����ٿ�tl���@�[c���3@m����!?QH���@�����ٿ�tl���@�[c���3@m����!?QH���@]�\�ٿ�N��y?�@��v=�3@���͉�!?�	��|��@]�\�ٿ�N��y?�@��v=�3@���͉�!?�	��|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@:�E��ٿ)�|D�@��$o�3@�����!?C���|��@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�J,��ٿ>�W�
	�@a+�&�3@����!?0=�a���@�ٱcg�ٿ�����@���dX�3@�A<���!?��Sq�)�@�ٱcg�ٿ�����@���dX�3@�A<���!?��Sq�)�@�ٱcg�ٿ�����@���dX�3@�A<���!?��Sq�)�@�ٱcg�ٿ�����@���dX�3@�A<���!?��Sq�)�@�ٱcg�ٿ�����@���dX�3@�A<���!?��Sq�)�@?T� e�ٿ��T�i�@�zC��3@�+��!?�a�tKy�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@;4����ٿ
�/��0�@��w9[�3@n*�ͼ�!?t�|3W�@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@��7��ٿ��'(4��@}Zr���3@l�i*��!?d����@l�$6�ٿ�������@�pLYS�3@�6�2��!?_Ld��@l�$6�ٿ�������@�pLYS�3@�6�2��!?_Ld��@l�$6�ٿ�������@�pLYS�3@�6�2��!?_Ld��@l�$6�ٿ�������@�pLYS�3@�6�2��!?_Ld��@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�J��ٿ��Q�2�@��ZF�3@�A���!?�J��R�@�z��@�ٿ������@k���E�3@8����!?F �9^:�@J�{�Қٿfs���@Q�#��3@�x$��!?���I��@_-#QR�ٿ̿��@�ȋ�3@���!?P�=�rn�@_-#QR�ٿ̿��@�ȋ�3@���!?P�=�rn�@_-#QR�ٿ̿��@�ȋ�3@���!?P�=�rn�@_-#QR�ٿ̿��@�ȋ�3@���!?P�=�rn�@_-#QR�ٿ̿��@�ȋ�3@���!?P�=�rn�@��+�ѣٿ��q*��@)��!�3@B�$Nt�!?j���i7�@��+�ѣٿ��q*��@)��!�3@B�$Nt�!?j���i7�@�.~�4�ٿ�
<*�R�@(S���3@o��#��!?���jt!�@��tŨٿJ$�}��@�d���3@�~	k��!?�Bd��@��tŨٿJ$�}��@�d���3@�~	k��!?�Bd��@>2W�ٿ�@�F��@�+|G��3@C��@�!?��N-p��@>2W�ٿ�@�F��@�+|G��3@C��@�!?��N-p��@O��7>�ٿ�S�Ц�@�ɹ��3@_��4�!?,�[����@O��7>�ٿ�S�Ц�@�ɹ��3@_��4�!?,�[����@O��7>�ٿ�S�Ц�@�ɹ��3@_��4�!?,�[����@q��T{�ٿ��ИK�@Ǜ����3@Mӡ]N�!?9ҚI��@,dG��ٿ�ϵ�X�@U�R<�3@�:l�e�!?�j�[?�@,dG��ٿ�ϵ�X�@U�R<�3@�:l�e�!?�j�[?�@,dG��ٿ�ϵ�X�@U�R<�3@�:l�e�!?�j�[?�@,dG��ٿ�ϵ�X�@U�R<�3@�:l�e�!?�j�[?�@���T�ٿ�I=����@W�����3@޲#o�!?Y�L�d��@e� ��ٿ<�*k8��@<��n�3@I��1�!?�5���'�@e� ��ٿ<�*k8��@<��n�3@I��1�!?�5���'�@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@P����ٿ o	��@h~2�p�3@��s'
�!?[���{��@l����ٿ�QI�o�@W��V��3@�B���!?S��/u�@l����ٿ�QI�o�@W��V��3@�B���!?S��/u�@�x�ٿ�6
�{�@���3�3@V��j�!?�"�P/�@�x�ٿ�6
�{�@���3�3@V��j�!?�"�P/�@�A/�~�ٿ�׎g~��@�9��+�3@M	��>�!?6n����@�A/�~�ٿ�׎g~��@�9��+�3@M	��>�!?6n����@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@w[��_�ٿ�+�"�,�@H�>��3@�]�2�!?g�L��+�@�:E�a�ٿ�K2vD��@Mc{�R�3@����А!?�V]F���@�:E�a�ٿ�K2vD��@Mc{�R�3@����А!?�V]F���@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@i��8�ٿ�i��V��@3è�~�3@z���!?#!v8r��@�NЄ��ٿ��1�C�@{}����3@©��ϐ!?���N�@�NЄ��ٿ��1�C�@{}����3@©��ϐ!?���N�@�NЄ��ٿ��1�C�@{}����3@©��ϐ!?���N�@�NЄ��ٿ��1�C�@{}����3@©��ϐ!?���N�@8\�z�ٿ&�r����@���!�3@	>	�!?��	��@8\�z�ٿ&�r����@���!�3@	>	�!?��	��@ա���ٿj�'-�@)���3@�0���!?�j^��@ա���ٿj�'-�@)���3@�0���!?�j^��@ա���ٿj�'-�@)���3@�0���!?�j^��@ա���ٿj�'-�@)���3@�0���!?�j^��@ա���ٿj�'-�@)���3@�0���!?�j^��@ա���ٿj�'-�@)���3@�0���!?�j^��@�_#gj�ٿdD�D���@���H�3@~��+��!?�6���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@��m��ٿ���M�@d���-�3@k`W��!?~*8���@�4l�ٿ���'9E�@f�T+�3@PV���!?�9����@�4l�ٿ���'9E�@f�T+�3@PV���!?�9����@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@�n��ٿ��}�S�@(jaF�3@Bɋmڐ!?�K�,t��@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@S`{��ٿ4�����@�NV�J�3@�p3?��!?�x�|���@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@��R�5�ٿ�}GԱ��@���++�3@��Kz�!?S���$�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�E$�B�ٿ<���C��@�R)��3@7}��ϐ!?�4�ca�@�i����ٿ��I�a��@6�,��3@W����!?u�&�͇�@�i����ٿ��I�a��@6�,��3@W����!?u�&�͇�@�i����ٿ��I�a��@6�,��3@W����!?u�&�͇�@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�Dݳ�ٿ|�b���@*o���3@�;�e��!?�lX.���@�62짢ٿ�h�b�@=��3@����!?��p!���@I�9�ٿ��L�s��@�S� �3@h��g��!?�i��a�@I�9�ٿ��L�s��@�S� �3@h��g��!?�i��a�@I�9�ٿ��L�s��@�S� �3@h��g��!?�i��a�@I�9�ٿ��L�s��@�S� �3@h��g��!?�i��a�@iSh��ٿ��܉u.�@QzZf�3@�lÐ!?re(9�@iSh��ٿ��܉u.�@QzZf�3@�lÐ!?re(9�@iSh��ٿ��܉u.�@QzZf�3@�lÐ!?re(9�@h��q�ٿQ	��3?�@A�~ZW�3@��~��!?9 ��p�@h��q�ٿQ	��3?�@A�~ZW�3@��~��!?9 ��p�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@LǸtr�ٿ�V�~�@�Yf��3@��.���!?h���*�@j�]z�ٿ�6u�~��@Ss��K�3@$�ߖ�!?��otu'�@�#�J �ٿC��PZt�@<T���3@�p�:6�!?o�.����@�#�J �ٿC��PZt�@<T���3@�p�:6�!?o�.����@$Z��$�ٿN?��/�@>E��3@�W1���!?ꜘ Y��@$Z��$�ٿN?��/�@>E��3@�W1���!?ꜘ Y��@$Z��$�ٿN?��/�@>E��3@�W1���!?ꜘ Y��@
<#���ٿ�?�S���@t��Q��3@a��e%�!?�+����@3�D�ٿ���@��@�ʌ�H�3@�Ш�+�!?�-o�w��@3�D�ٿ���@��@�ʌ�H�3@�Ш�+�!?�-o�w��@3�D�ٿ���@��@�ʌ�H�3@�Ш�+�!?�-o�w��@3�D�ٿ���@��@�ʌ�H�3@�Ш�+�!?�-o�w��@3�D�ٿ���@��@�ʌ�H�3@�Ш�+�!?�-o�w��@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@p�v��ٿXs����@*�&'��3@/L�2�!?�f95�-�@O�~+�ٿ��2�i��@�vU���3@�E���!?ı�o��@O�~+�ٿ��2�i��@�vU���3@�E���!?ı�o��@O�~+�ٿ��2�i��@�vU���3@�E���!?ı�o��@O�~+�ٿ��2�i��@�vU���3@�E���!?ı�o��@O�~+�ٿ��2�i��@�vU���3@�E���!?ı�o��@7C����ٿK;n7o�@)��(�3@�>�ֵ�!?O�����@7C����ٿK;n7o�@)��(�3@�>�ֵ�!?O�����@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@���ٿ{2xȡ�@����3@#�ε��!?HJ7�J��@0�V�/�ٿN�d���@W����3@���m�!?��e��@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@�z{ʄ�ٿLn&�B�@o��#]�3@4�W��!?{T��:�@`t�Μٿ��`�'��@��h��3@��JԐ!?2�^����@`t�Μٿ��`�'��@��h��3@��JԐ!?2�^����@`t�Μٿ��`�'��@��h��3@��JԐ!?2�^����@`t�Μٿ��`�'��@��h��3@��JԐ!?2�^����@`t�Μٿ��`�'��@��h��3@��JԐ!?2�^����@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@a&�_�ٿv�i��=�@9T�4>�3@�酽�!?���K�x�@*�̙ �ٿ{6����@PC=�W�3@ۤ�힐!?9�[�@*�̙ �ٿ{6����@PC=�W�3@ۤ�힐!?9�[�@*�̙ �ٿ{6����@PC=�W�3@ۤ�힐!?9�[�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@r�u��ٿ���}vN�@5�vD��3@|�E��!?��~]�&�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@����0�ٿ��a�R�@�X<(_�3@�᯳��!?�h|�@R��E��ٿDt�j��@��	���3@<K��!?���/��@R��E��ٿDt�j��@��	���3@<K��!?���/��@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@b��:�ٿ���R���@�^��>�3@hb˃ِ!?�,�����@�հ:��ٿ)�����@)�$���3@����ِ!?��s�!��@�հ:��ٿ)�����@)�$���3@����ِ!?��s�!��@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�!��բٿ�&����@f���3@"�_�!?I*���@�0:Z�ٿ@&�
%��@ ����3@B��ؐ!?3ng�p�@��Sz�ٿ G�ȕ�@�.N��3@���U��!?��&���@��Sz�ٿ G�ȕ�@�.N��3@���U��!?��&���@��Sz�ٿ G�ȕ�@�.N��3@���U��!?��&���@��Sz�ٿ G�ȕ�@�.N��3@���U��!?��&���@�P��r�ٿ>N�l�7�@������3@�c*���!?�+��Ӱ�@�P��r�ٿ>N�l�7�@������3@�c*���!?�+��Ӱ�@�P��r�ٿ>N�l�7�@������3@�c*���!?�+��Ӱ�@�P��r�ٿ>N�l�7�@������3@�c*���!?�+��Ӱ�@ɼ'8��ٿ�%�$�@	_��z 4@;(��!?�oNЬ��@ɼ'8��ٿ�%�$�@	_��z 4@;(��!?�oNЬ��@ɼ'8��ٿ�%�$�@	_��z 4@;(��!?�oNЬ��@ɼ'8��ٿ�%�$�@	_��z 4@;(��!?�oNЬ��@ɼ'8��ٿ�%�$�@	_��z 4@;(��!?�oNЬ��@���N��ٿU���@�?�3@�`�[�!?��\7i�@���N��ٿU���@�?�3@�`�[�!?��\7i�@��K��ٿ4"L#���@�T$��3@�[���!? ���e��@��K��ٿ4"L#���@�T$��3@�[���!? ���e��@C7�ɣٿ�����@kQ�'��3@�����!?�#3��q�@C7�ɣٿ�����@kQ�'��3@�����!?�#3��q�@C7�ɣٿ�����@kQ�'��3@�����!?�#3��q�@OB)��ٿ��T�?��@D�N�S�3@s�x���!?!���l��@����ٿ��<+j-�@'���>�3@�s�W��!?��:��@����ٿ��<+j-�@'���>�3@�s�W��!?��:��@����ٿ��<+j-�@'���>�3@�s�W��!?��:��@����ٿ��<+j-�@'���>�3@�s�W��!?��:��@�C����ٿ��\E��@B��ۃ�3@�&�B��!?>�ь���@�C����ٿ��\E��@B��ۃ�3@�&�B��!?>�ь���@�C����ٿ��\E��@B��ۃ�3@�&�B��!?>�ь���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@���z�ٿ����m�@���3��3@�CX��!?=�8���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@"L��Ρٿ���m���@?H���3@��@ǐ!?m���@GOH�Y�ٿ �t��@'�k�Y�3@@���!?��.�)q�@GOH�Y�ٿ �t��@'�k�Y�3@@���!?��.�)q�@GOH�Y�ٿ �t��@'�k�Y�3@@���!?��.�)q�@GOH�Y�ٿ �t��@'�k�Y�3@@���!?��.�)q�@�����ٿ�q�נ��@�.;��3@4�D���!?����d�@�����ٿ�q�נ��@�.;��3@4�D���!?����d�@����ٿ��H
Hi�@~����3@��⭲�!?�c�����@����ٿ��H
Hi�@~����3@��⭲�!?�c�����@����ٿ��H
Hi�@~����3@��⭲�!?�c�����@}���ٿ�+"���@��J�3�3@�HJ�!?'p(ݟ�@}���ٿ�+"���@��J�3�3@�HJ�!?'p(ݟ�@}���ٿ�+"���@��J�3�3@�HJ�!?'p(ݟ�@}���ٿ�+"���@��J�3�3@�HJ�!?'p(ݟ�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@���ٿ6�'���@8���H�3@��y��!?HX�oj�@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@��QK�ٿ�s��a��@��_��3@-�	wӐ!?6t�`��@ih�|��ٿ�b ���@��y�o�3@�f���!?䚎�Z�@ih�|��ٿ�b ���@��y�o�3@�f���!?䚎�Z�@ih�|��ٿ�b ���@��y�o�3@�f���!?䚎�Z�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@J(S/�ٿ�Dw�
5�@׉ر5�3@5�\!?�zd�k�@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@3�?u�ٿ�=�g��@��pЖ�3@���ʐ!?�b�N���@�7�[�ٿ!P�ܽ9�@�4���3@4�s�!?Zl9���@�7�[�ٿ!P�ܽ9�@�4���3@4�s�!?Zl9���@�7�[�ٿ!P�ܽ9�@�4���3@4�s�!?Zl9���@�x6�I�ٿC��s���@>�����3@_����!?�æ����@�x6�I�ٿC��s���@>�����3@_����!?�æ����@�x6�I�ٿC��s���@>�����3@_����!?�æ����@�x6�I�ٿC��s���@>�����3@_����!?�æ����@�p���ٿ���(��@��E���3@n|,�!?�X蝵��@�p���ٿ���(��@��E���3@n|,�!?�X蝵��@�p���ٿ���(��@��E���3@n|,�!?�X蝵��@�5A�ٿO�p$�@�%����3@@K"�Ґ!?��c��@�5A�ٿO�p$�@�%����3@@K"�Ґ!?��c��@0��5��ٿ�A�b��@�rL�C�3@��!?G��I��@�01�ٿ>&<yq'�@#�����3@�>J+�!?��P����@�01�ٿ>&<yq'�@#�����3@�>J+�!?��P����@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@� �T$�ٿ&3��ן�@��#��3@���l��!?������@��KՠٿS�����@W��w-�3@���Y��!?�k�$�[�@�-D�ٿњK/���@`��g��3@�%����!?`�Y���@�-D�ٿњK/���@`��g��3@�%����!?`�Y���@�-D�ٿњK/���@`��g��3@�%����!?`�Y���@�-D�ٿњK/���@`��g��3@�%����!?`�Y���@֓𳸠ٿ����?G�@p�
�3@`�TC�!?��H	$�@֓𳸠ٿ����?G�@p�
�3@`�TC�!?��H	$�@֓𳸠ٿ����?G�@p�
�3@`�TC�!?��H	$�@��j.a�ٿp-�����@bOJ�t�3@h:V�ސ!?�����@��j.a�ٿp-�����@bOJ�t�3@h:V�ސ!?�����@��j.a�ٿp-�����@bOJ�t�3@h:V�ސ!?�����@��j.a�ٿp-�����@bOJ�t�3@h:V�ސ!?�����@)��1��ٿq�F��
�@��^��3@�^ ��!?��=�v�@7�C�^�ٿ���Y�@4����3@��0��!?�\';%�@����ٿ��^�XI�@��ך;�3@���dM�!?=���U��@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��L��ٿ�F{��n�@z���<�3@�V���!?�Ih�e�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@��]P��ٿ�[A���@u�94�3@M�7���!?C%:�$f�@�D[���ٿM�ia��@�G���3@��M�V�!?Mh�mɠ�@�D[���ٿM�ia��@�G���3@��M�V�!?Mh�mɠ�@�D[���ٿM�ia��@�G���3@��M�V�!?Mh�mɠ�@B��K�ٿ���N3D�@�-�aV�3@K�́��!?�X>�Cw�@B��K�ٿ���N3D�@�-�aV�3@K�́��!?�X>�Cw�@�I���ٿ��4���@� �k�3@���C�!?&��Y���@�I���ٿ��4���@� �k�3@���C�!?&��Y���@�I���ٿ��4���@� �k�3@���C�!?&��Y���@�I���ٿ��4���@� �k�3@���C�!?&��Y���@�I���ٿ��4���@� �k�3@���C�!?&��Y���@�I���ٿ��4���@� �k�3@���C�!?&��Y���@v�s�٘ٿ��J��@k��Ng�3@�6���!?F�L�!��@�D��ٿ��TL�)�@5X�X�3@��λ�!?> Nke*�@�D��ٿ��TL�)�@5X�X�3@��λ�!?> Nke*�@�D��ٿ��TL�)�@5X�X�3@��λ�!?> Nke*�@��It�ٿ�`����@�x	ʚ�3@�J�ڐ!?$;U���@��It�ٿ�`����@�x	ʚ�3@�J�ڐ!?$;U���@��It�ٿ�`����@�x	ʚ�3@�J�ڐ!?$;U���@��It�ٿ�`����@�x	ʚ�3@�J�ڐ!?$;U���@̑w���ٿ�)�+#�@��ϛ%�3@{�H���!?8��S���@̑w���ٿ�)�+#�@��ϛ%�3@{�H���!?8��S���@s�R��ٿ)�����@��A�3@Y͘��!?�B�z�%�@s�R��ٿ)�����@��A�3@Y͘��!?�B�z�%�@s�R��ٿ)�����@��A�3@Y͘��!?�B�z�%�@��c��ٿ�	lδ�@~�*y�3@2��-�!?�Y���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@X	���ٿ���-Z��@��6�3@���Ɨ�!? oY���@��>�ٿ1�?�(/�@�V.9�3@�Y}��!?�wI�A�@�K�3�ٿb�u2��@�&�8�3@��Ő!?G�e�'��@�K�3�ٿb�u2��@�&�8�3@��Ő!?G�e�'��@�K�3�ٿb�u2��@�&�8�3@��Ő!?G�e�'��@�K�3�ٿb�u2��@�&�8�3@��Ő!?G�e�'��@O��{�ٿ�@��H��@�\����3@Y+X:�!?5,H���@�O��ٿV�RQ�@Ȁ� 0�3@�;��!?��y]&�@�O��ٿV�RQ�@Ȁ� 0�3@�;��!?��y]&�@�O��ٿV�RQ�@Ȁ� 0�3@�;��!?��y]&�@%E^�ٿ��[���@Ƅk*�3@�1Xm��!?CD��c�@%E^�ٿ��[���@Ƅk*�3@�1Xm��!?CD��c�@%E^�ٿ��[���@Ƅk*�3@�1Xm��!?CD��c�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@~!�0ܤٿAᗮcL�@�T�G�3@'K�Ӑ!?s��e�@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�"f[��ٿ��
�R/�@c���3@�}���!?;��_r��@�0_�ٿ�p�&�4�@�����3@�B�Ӑ!?�n�.���@�0_�ٿ�p�&�4�@�����3@�B�Ӑ!?�n�.���@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@%,��ٿ�8���@/i	��3@�ׂ��!?j�;YV�@N,���ٿ�9]�7��@C����3@��ؿ�!?P3�O�L�@b?���ٿ������@R7���3@������!?�fS�@b?���ٿ������@R7���3@������!?�fS�@b?���ٿ������@R7���3@������!?�fS�@N�A�ٿ��#)W�@�D��3@G��)��!?�K�yLJ�@��=,�ٿd�(�n�@��~�3@���ؐ!?#��+ �@Q?֝C�ٿ���)��@ҜK�L�3@Meg��!?�:5�4d�@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@�f{�ٿp�0s�@�:��s�3@S݃��!?��{"��@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@`/�6!�ٿ�t��<Z�@����3@��M���!?�;��y�@�n�?�ٿ����vM�@�t�3@HZܐ!?�|�B�@�n�?�ٿ����vM�@�t�3@HZܐ!?�|�B�@�6��ٿxN�G�R�@��߾b�3@�����!?�!6�+�@k��詞ٿ�>��@Q�@��
��3@1�x��!?���a��@k��詞ٿ�>��@Q�@��
��3@1�x��!?���a��@k��詞ٿ�>��@Q�@��
��3@1�x��!?���a��@k��詞ٿ�>��@Q�@��
��3@1�x��!?���a��@��"�?�ٿ7�����@�K'q��3@��$���!?���ı��@��"�?�ٿ7�����@�K'q��3@��$���!?���ı��@��"�?�ٿ7�����@�K'q��3@��$���!?���ı��@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�M{�ٿq�x�$�@+$����3@�G�ڌ�!?s�8P���@�Ǚ��ٿo�t*��@c���3@N	B{�!?��ONG�@�Ǚ��ٿo�t*��@c���3@N	B{�!?��ONG�@�Ǚ��ٿo�t*��@c���3@N	B{�!?��ONG�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@[�����ٿw�SǓ�@iT�>��3@6�
si�!?��c�F�@�I5��ٿ	�Ӣݗ�@>�ּ&�3@&v�L��!?$Y�[��@�I5��ٿ	�Ӣݗ�@>�ּ&�3@&v�L��!?$Y�[��@�I5��ٿ	�Ӣݗ�@>�ּ&�3@&v�L��!?$Y�[��@�I5��ٿ	�Ӣݗ�@>�ּ&�3@&v�L��!?$Y�[��@�;���ٿ�o`h�7�@�����3@��'��!?����l��@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@�pcK��ٿb�6w�@E'�R��3@|��h�!?z֔�n�@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@����&�ٿ: �@�L�e�3@���#��!?�:5~@��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@;�3�^�ٿ��!|���@�w!�>�3@`?j'��!?����L��@\����ٿ�&�\��@)�	l�3@\ZKq�!?}1͛�@b�O1�ٿR���o�@ ��t�3@l޿룐!?��k��Y�@b�O1�ٿR���o�@ ��t�3@l޿룐!?��k��Y�@b�O1�ٿR���o�@ ��t�3@l޿룐!?��k��Y�@b�O1�ٿR���o�@ ��t�3@l޿룐!?��k��Y�@b�O1�ٿR���o�@ ��t�3@l޿룐!?��k��Y�@�^���ٿ�I�E:�@P����3@w4GI��!?�n"� �@����#�ٿ�����@���x�3@	W�8n�!?e�2\2B�@����#�ٿ�����@���x�3@	W�8n�!?e�2\2B�@����#�ٿ�����@���x�3@	W�8n�!?e�2\2B�@����#�ٿ�����@���x�3@	W�8n�!?e�2\2B�@x�V�ٿ�,]S��@�'��3@�9�Pɐ!?̀,�"��@x�V�ٿ�,]S��@�'��3@�9�Pɐ!?̀,�"��@x�V�ٿ�,]S��@�'��3@�9�Pɐ!?̀,�"��@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@����a�ٿU�%l<�@EK ��3@^����!?}=�2���@?1c�)�ٿ$yKm��@�QK[��3@}��ܿ�!?�fo�C�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��z�ٿ�V-�H�@���Tc�3@P�$��!?����ơ�@��7'�ٿ�@�Y-N�@�=@��3@��Rl�!?�����@��7'�ٿ�@�Y-N�@�=@��3@��Rl�!?�����@��7'�ٿ�@�Y-N�@�=@��3@��Rl�!?�����@��7'�ٿ�@�Y-N�@�=@��3@��Rl�!?�����@𣬷Q�ٿ������@�̎���3@4Q��q�!?}�a��@𣬷Q�ٿ������@�̎���3@4Q��q�!?}�a��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@&�}�ٿ��-j�$�@���u�3@�?�m��!?P��@��@\����ٿ�w$�n�@ "~A�3@=�����!?�(C�Q�@\����ٿ�w$�n�@ "~A�3@=�����!?�(C�Q�@\����ٿ�w$�n�@ "~A�3@=�����!?�(C�Q�@\����ٿ�w$�n�@ "~A�3@=�����!?�(C�Q�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@�|��6�ٿ��D���@G3����3@��!�Ґ!?����La�@.I,�A�ٿ�a�+yg�@�j���3@[Z�Ɛ!?��DW�@.I,�A�ٿ�a�+yg�@�j���3@[Z�Ɛ!?��DW�@.I,�A�ٿ�a�+yg�@�j���3@[Z�Ɛ!?��DW�@.I,�A�ٿ�a�+yg�@�j���3@[Z�Ɛ!?��DW�@.I,�A�ٿ�a�+yg�@�j���3@[Z�Ɛ!?��DW�@�=�0�ٿbgw���@��#��3@V�MΔ�!?�@�\߰�@�=�0�ٿbgw���@��#��3@V�MΔ�!?�@�\߰�@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@G�x��ٿ��(4��@ʨ���3@I��ې!?�H $��@��&��ٿS����?�@�%���3@1C@�ѐ!?p��#X�@��&��ٿS����?�@�%���3@1C@�ѐ!?p��#X�@��&��ٿS����?�@�%���3@1C@�ѐ!?p��#X�@�O����ٿ�'����@�j��W�3@lh��!?�*�~wS�@�O����ٿ�'����@�j��W�3@lh��!?�*�~wS�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@V����ٿdT��'�@�ܜ�3@%���̐!?�ڢ@D�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@J��J�ٿ�W����@���S�3@�Ns�!?���MI�@�����ٿ"�d�@R�b&��3@��
�ސ!?m��G{O�@�����ٿ"�d�@R�b&��3@��
�ސ!?m��G{O�@1��6X�ٿ��yHc��@�%}��3@Cd=}��!?���|�@��_l��ٿ6L�c�@"/\d��3@�%
�!?/:8���@��_l��ٿ6L�c�@"/\d��3@�%
�!?/:8���@W�a�6�ٿ�zm��@�"n��3@ta�ǐ!?0�6��,�@�Z7��ٿ6	�T�@�" U��3@��Ͼ�!?-�����@�Z7��ٿ6	�T�@�" U��3@��Ͼ�!?-�����@M"!� �ٿ��ZԤ`�@�1/��3@�,�Kː!?æ�3ݷ�@�w�*�ٿ�jC�_Q�@�P���3@�u�㾐!?��%Eo�@�D�n(�ٿ@�����@2�U�W�3@�T��ʐ!?��s��{�@�D�n(�ٿ@�����@2�U�W�3@�T��ʐ!?��s��{�@�D�n(�ٿ@�����@2�U�W�3@�T��ʐ!?��s��{�@�D�n(�ٿ@�����@2�U�W�3@�T��ʐ!?��s��{�@�D�n(�ٿ@�����@2�U�W�3@�T��ʐ!?��s��{�@i]�(�ٿ������@b'���3@�c���!?g�����@i]�(�ٿ������@b'���3@�c���!?g�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@ͣc==�ٿ���e�@��&f�3@`Ȑ!?�#�����@�T�
D�ٿ��ul�7�@x���u�3@�p���!?�14��&�@4�=H��ٿ�J���@ �mt)�3@��t�!?�5nP51�@4�=H��ٿ�J���@ �mt)�3@��t�!?�5nP51�@�\3�ٿ �8��@�S�$Y�3@�a�i�!?�:�`��@�n���ٿ�E�Ml�@}�v4�3@n�|�>�!?ᴚqo~�@�x�̾�ٿ��k��@��`���3@I��r�!?�J���@�x�̾�ٿ��k��@��`���3@I��r�!?�J���@�x�̾�ٿ��k��@��`���3@I��r�!?�J���@����/�ٿoT*ن��@�߲���3@�UAu�!?r$;����@����/�ٿoT*ن��@�߲���3@�UAu�!?r$;����@����/�ٿoT*ن��@�߲���3@�UAu�!?r$;����@��uX��ٿ��=l��@"}:���3@" ���!?�j_��@��uX��ٿ��=l��@"}:���3@" ���!?�j_��@�bw/ܦٿ�@����@,��.�3@���Jy�!?K�y���@�bw/ܦٿ�@����@,��.�3@���Jy�!?K�y���@�bw/ܦٿ�@����@,��.�3@���Jy�!?K�y���@��� �ٿR胝��@�q�y�3@-ZDm��!?	&ͩ��@��� �ٿR胝��@�q�y�3@-ZDm��!?	&ͩ��@��� �ٿR胝��@�q�y�3@-ZDm��!?	&ͩ��@��� �ٿR胝��@�q�y�3@-ZDm��!?	&ͩ��@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@�$Qs�ٿ���sh�@Z�(_�3@�3S��!?Z��H���@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@���P�ٿ5�=Ԙ��@�נ}��3@2L;�֐!?Q���8��@0jz���ٿF��z�@̀�('�3@�v�Ɛ!?DEtC�:�@0jz���ٿF��z�@̀�('�3@�v�Ɛ!?DEtC�:�@	���ٿ7���3�@S8(�3@	oא!?��xn*�@	���ٿ7���3�@S8(�3@	oא!?��xn*�@	���ٿ7���3�@S8(�3@	oא!?��xn*�@	���ٿ7���3�@S8(�3@	oא!?��xn*�@͓��̢ٿ�g���{�@]�b��3@�����!?� ���@͓��̢ٿ�g���{�@]�b��3@�����!?� ���@͓��̢ٿ�g���{�@]�b��3@�����!?� ���@͓��̢ٿ�g���{�@]�b��3@�����!?� ���@��#�ɢٿ�+���@H;Ei�3@P�+S�!?�����@��#�ɢٿ�+���@H;Ei�3@P�+S�!?�����@��#�ɢٿ�+���@H;Ei�3@P�+S�!?�����@��#�ɢٿ�+���@H;Ei�3@P�+S�!?�����@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@�Z��ٿ&*��s`�@f�ԕ��3@�ۗᑐ!?A&z]	��@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@k��l�ٿFp��/@�@�� JH�3@}.��!?zj�����@��I��ٿ^7ٸ��@��Z��3@�d�GŐ!?^�X�;�@~\I}�ٿ�Ⱥ��5�@O�4��3@�H�!?�g]	i��@~\I}�ٿ�Ⱥ��5�@O�4��3@�H�!?�g]	i��@!#R
��ٿ�"�<f��@�$�e��3@�vʪ�!?�V�n I�@����ٿ#t��:��@�{�
��3@�����!?�A{�@����ٿ#t��:��@�{�
��3@�����!?�A{�@����ٿ#t��:��@�{�
��3@�����!?�A{�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@;tl&�ٿMЁ/�`�@����3@q�]͐!?H�1sj�@sT���ٿ�ɮ����@��}w��3@�K߀��!?�?)��`�@sT���ٿ�ɮ����@��}w��3@�K߀��!?�?)��`�@>M��ٿgi�����@�Ҧ�_�3@C�]���!? �e4$<�@>M��ٿgi�����@�Ҧ�_�3@C�]���!? �e4$<�@>M��ٿgi�����@�Ҧ�_�3@C�]���!? �e4$<�@>M��ٿgi�����@�Ҧ�_�3@C�]���!? �e4$<�@>M��ٿgi�����@�Ҧ�_�3@C�]���!? �e4$<�@C��U�ٿ�)�D�"�@5�\���3@�,?��!?��ގ~�@7�	��ٿ���"���@KLܾ�3@o����!?������@���I��ٿՃWH.y�@ɗ��3@&*kw��!?������@���I��ٿՃWH.y�@ɗ��3@&*kw��!?������@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@�7�!�ٿ5Z���@�+0f�3@��iʐ!?2L�r�}�@QQ�9�ٿ���t0�@ +Hh�3@�C��$�!?�����@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@C3_���ٿ)?�[�@N����3@���X�!?6t;?��@���O�ٿ���c��@�o˺�3@-fiA��!?F>qA��@Ke�Y�ٿ[������@��@�,�3@Gs��U�!?�K��@�@Ke�Y�ٿ[������@��@�,�3@Gs��U�!?�K��@�@Ke�Y�ٿ[������@��@�,�3@Gs��U�!?�K��@�@Ke�Y�ٿ[������@��@�,�3@Gs��U�!?�K��@�@����ٿ�,e�t�@�u����3@�/�姐!?q���;Y�@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@cd~�ԟٿ>����!�@�A�Ѡ�3@�g�2��!?L\T���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�)�r�ٿ�k����@�!]R�3@� ��֐!?XXu[���@�j�	?�ٿ�V��J�@X5����3@�\vϳ�!?C�:.\6�@�j�	?�ٿ�V��J�@X5����3@�\vϳ�!?C�:.\6�@�j�	?�ٿ�V��J�@X5����3@�\vϳ�!?C�:.\6�@�j�	?�ٿ�V��J�@X5����3@�\vϳ�!?C�:.\6�@�[VԤٿ~]"���@Ĵ*�3@��2��!?T/�����@�[VԤٿ~]"���@Ĵ*�3@��2��!?T/�����@�[VԤٿ~]"���@Ĵ*�3@��2��!?T/�����@�[VԤٿ~]"���@Ĵ*�3@��2��!?T/�����@g��z�ٿ��2�I�@�aD}�3@HG�p��!?S��Ve�@g��z�ٿ��2�I�@�aD}�3@HG�p��!?S��Ve�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@�#�}�ٿF,+[t9�@���c��3@�	���!?	�ҷ<r�@GB�)��ٿaF�eҌ�@�/�hy�3@ݦ1���!?B#�9��@��!uq�ٿ����S��@:�}i��3@��8���!?��i?��@#�
S�ٿ~���D�@4��W�3@��Ẑ!?�!�>[�@fd�aA�ٿM���݉�@�④��3@	D�8̐!?r肨���@ԋ]b��ٿ�i��p��@r�ts��3@\E��c�!?Wm��'��@ԋ]b��ٿ�i��p��@r�ts��3@\E��c�!?Wm��'��@ԋ]b��ٿ�i��p��@r�ts��3@\E��c�!?Wm��'��@ԋ]b��ٿ�i��p��@r�ts��3@\E��c�!?Wm��'��@ԋ]b��ٿ�i��p��@r�ts��3@\E��c�!?Wm��'��@\��;�ٿϩC�z�@��#�L�3@�I�[�!?@h&���@1r�Z�ٿ��|WG�@k{� �3@�r���!?��v�E�@1r�Z�ٿ��|WG�@k{� �3@�r���!?��v�E�@1r�Z�ٿ��|WG�@k{� �3@�r���!?��v�E�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@��V�o�ٿ˚!O��@/���3@S0
���!?#[�J�|�@ۆ-��ٿ�6�o���@�}���3@�&���!?E8�	�@ۆ-��ٿ�6�o���@�}���3@�&���!?E8�	�@ۆ-��ٿ�6�o���@�}���3@�&���!?E8�	�@ۆ-��ٿ�6�o���@�}���3@�&���!?E8�	�@ۆ-��ٿ�6�o���@�}���3@�&���!?E8�	�@�c~�ٿ�Kf>�g�@+_����3@�����!?�3����@��d��ٿ>;�\�@㹔�B�3@t_���!?Q�̆��@��d��ٿ>;�\�@㹔�B�3@t_���!?Q�̆��@��d��ٿ>;�\�@㹔�B�3@t_���!?Q�̆��@��d��ٿ>;�\�@㹔�B�3@t_���!?Q�̆��@�3�ٿ-�%o[�@U�
�N�3@c�����!?z��	�@�3�ٿ-�%o[�@U�
�N�3@c�����!?z��	�@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@�����ٿ�����B�@Ò�7��3@�˱��!?e=���@��[��ٿ	���H�@���V-�3@��f���!?xb&
o��@��[��ٿ	���H�@���V-�3@��f���!?xb&
o��@��[��ٿ	���H�@���V-�3@��f���!?xb&
o��@y�xಥٿ7�H["c�@r"���3@��2zА!?������@y�xಥٿ7�H["c�@r"���3@��2zА!?������@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@㼘���ٿى/m��@�`�S��3@�9T�!?zn�%��@�@S��ٿz���U�@-r���3@�&xʐ!?�l�:���@�@S��ٿz���U�@-r���3@�&xʐ!?�l�:���@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@Vw�,t�ٿ�GA�a@�@m�`o�3@؀ިߐ!?"�I��@�$�雥ٿ�fH���@,����3@�I���!?? �!�n�@�$�雥ٿ�fH���@,����3@�I���!?? �!�n�@�u-L��ٿ�0�Ե��@�����3@��^��!?^G��"~�@�u-L��ٿ�0�Ե��@�����3@��^��!?^G��"~�@�u-L��ٿ�0�Ե��@�����3@��^��!?^G��"~�@�u-L��ٿ�0�Ե��@�����3@��^��!?^G��"~�@���hi�ٿ�If}K�@�֟��3@o��!?{����@���hi�ٿ�If}K�@�֟��3@o��!?{����@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@A�]J��ٿZ��1��@��R#	�3@S���!?a�.�G�@��,��ٿb�x�y��@=ZzP�3@33�!?#�����@��,��ٿb�x�y��@=ZzP�3@33�!?#�����@��,��ٿb�x�y��@=ZzP�3@33�!?#�����@!��h�ٿ�ϗ��I�@���e�3@y�� ��!?4	|(`��@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@
J�[��ٿ�w��f��@�Cg���3@��x��!?�O�Y���@Tj�U2�ٿ|J���@h�����3@�e�}�!?��u��@n��ٿ!�!�W�@�gN&��3@a�#��!?R��_r��@n��ٿ!�!�W�@�gN&��3@a�#��!?R��_r��@n��ٿ!�!�W�@�gN&��3@a�#��!?R��_r��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@�6@�w�ٿ(���9��@����9�3@kVS͐!?��l"��@g1qح�ٿJrM��@�L�&�3@14���!?n���@g1qح�ٿJrM��@�L�&�3@14���!?n���@g1qح�ٿJrM��@�L�&�3@14���!?n���@g1qح�ٿJrM��@�L�&�3@14���!?n���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@i�����ٿ=�����@\|��3@�
�=��!?�C*/���@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@B8��ٿ��Sޜ��@P��Pw�3@al�w�!?�����@`�B$��ٿF��պ�@�j��w�3@���Dʐ!?Dh���@`�B$��ٿF��պ�@�j��w�3@���Dʐ!?Dh���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@*���ٿ}#K4�@��	?l�3@�~���!?"��w���@m!��}�ٿf��.-�@=����3@Z>f���!?�j+-��@m!��}�ٿf��.-�@=����3@Z>f���!?�j+-��@m!��}�ٿf��.-�@=����3@Z>f���!?�j+-��@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@�8�F2�ٿ=�@�@��,Hn�3@}6 ?��!?K�#�@\�ŧٿ����@ay��3@�
'O��!?��*�@\�ŧٿ����@ay��3@�
'O��!?��*�@\�ŧٿ����@ay��3@�
'O��!?��*�@\�ŧٿ����@ay��3@�
'O��!?��*�@d�����ٿ;1%D�8�@c�%��3@��X��!?�M���*�@�}rM��ٿ��FD��@K:5R�3@�>�w֐!?)#*h�@�}rM��ٿ��FD��@K:5R�3@�>�w֐!?)#*h�@����,�ٿ=% ���@��h6�3@�{�mȐ!?��	�r�@�����ٿVM�q�@���Y�3@����x�!?F�����@�����ٿVM�q�@���Y�3@����x�!?F�����@�����ٿVM�q�@���Y�3@����x�!?F�����@�����ٿVM�q�@���Y�3@����x�!?F�����@�����ٿVM�q�@���Y�3@����x�!?F�����@N�P��ٿH�<�@a�Y;$�3@�/o_�!?k����^�@'zyL�ٿy��X��@ o{��3@��;n�!?}��ˌ�@'zyL�ٿy��X��@ o{��3@��;n�!?}��ˌ�@'zyL�ٿy��X��@ o{��3@��;n�!?}��ˌ�@'zyL�ٿy��X��@ o{��3@��;n�!?}��ˌ�@'zyL�ٿy��X��@ o{��3@��;n�!?}��ˌ�@
�#�+�ٿ������@F�k���3@O[,{f�!?����@
�#�+�ٿ������@F�k���3@O[,{f�!?����@
�#�+�ٿ������@F�k���3@O[,{f�!?����@
�#�+�ٿ������@F�k���3@O[,{f�!?����@��]�ٿ������@?���T�3@�y�[��!?��u��@��]�ٿ������@?���T�3@�y�[��!?��u��@��]�ٿ������@?���T�3@�y�[��!?��u��@��]�ٿ������@?���T�3@�y�[��!?��u��@��n�ٿgF3q���@����3@k��d��!?���4ʌ�@��n�ٿgF3q���@����3@k��d��!?���4ʌ�@���1��ٿ��~)w/�@�
����3@��̝Ր!?= ��V��@���1��ٿ��~)w/�@�
����3@��̝Ր!?= ��V��@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@��ٿu��(�@wok��3@����!?��U���@�Ft��ٿ�9��@��4��3@fG�W$�!?�����=�@�Ft��ٿ�9��@��4��3@fG�W$�!?�����=�@�Ft��ٿ�9��@��4��3@fG�W$�!?�����=�@%u;m��ٿ����@�ӟ/��3@Roy���!?����J�@%u;m��ٿ����@�ӟ/��3@Roy���!?����J�@c�3R�ٿ���1�@Ԇ��)�3@��oe��!?�*���@c�3R�ٿ���1�@Ԇ��)�3@��oe��!?�*���@c�3R�ٿ���1�@Ԇ��)�3@��oe��!?�*���@c�3R�ٿ���1�@Ԇ��)�3@��oe��!?�*���@��B���ٿ]�����@m����3@�@�k��!?L�J��@��B���ٿ]�����@m����3@�@�k��!?L�J��@��B���ٿ]�����@m����3@�@�k��!?L�J��@P���ٿ�>�@k�m�3@��E~v�!?���)�@P���ٿ�>�@k�m�3@��E~v�!?���)�@P���ٿ�>�@k�m�3@��E~v�!?���)�@�kt��ٿu�O�B�@�=X��3@4�Lx��!?ʲ����@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@��o��ٿ1-��|��@ǒh��3@K~���!?We�h���@���ٿ�������@0hf��3@�\'@�!?���.��@жn�ٿ<���A��@��3@�@k��!?��(�D�@жn�ٿ<���A��@��3@�@k��!?��(�D�@�b͝ٿ��0��@�6K��3@wXo5 �!?��O�6�@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@���E��ٿH���r�@=1���3@�d�ѐ!?�Z�y��@eE��˝ٿ����� �@����3@J��!?�y%)�@eE��˝ٿ����� �@����3@J��!?�y%)�@eE��˝ٿ����� �@����3@J��!?�y%)�@eE��˝ٿ����� �@����3@J��!?�y%)�@eE��˝ٿ����� �@����3@J��!?�y%)�@;y��ٿq���h�@����3@�Q*�!?��҉���@;y��ٿq���h�@����3@�Q*�!?��҉���@ٮ��ġٿ~�|��@�d:E�3@Yg����!?j;����@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@^=x�J�ٿ����S�@�?��a�3@��:�!?v~�TmH�@�3�iK�ٿ ���4�@�r���3@չ�[��!?�Ki2���@�3�iK�ٿ ���4�@�r���3@չ�[��!?�Ki2���@�3�iK�ٿ ���4�@�r���3@չ�[��!?�Ki2���@�3�iK�ٿ ���4�@�r���3@չ�[��!?�Ki2���@�3�iK�ٿ ���4�@�r���3@չ�[��!?�Ki2���@^��R�ٿ��I�T�@�8���3@XnN*��!?H�4�;�@^��R�ٿ��I�T�@�8���3@XnN*��!?H�4�;�@��U��ٿrH�Q���@��s���3@_�!?1�E8�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@�(m��ٿ��a��@��bq�3@�kU�u�!?9���ٚ�@W�	��ٿ͎��8��@&/i{�3@��8vt�!?@�aJ�6�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@��y�8�ٿvu��@�^Z��3@��c���!?��ks'�@�M�u�ٿ�Y�%?�@�����3@wH'y��!?��h�p�@�M�u�ٿ�Y�%?�@�����3@wH'y��!?��h�p�@�M�u�ٿ�Y�%?�@�����3@wH'y��!?��h�p�@���⒣ٿں0#1d�@a��H.�3@?i��!?��O��"�@Q�#
�ٿ+���3�@��\S�3@�?t_��!?����@Q�#
�ٿ+���3�@��\S�3@�?t_��!?����@Q�#
�ٿ+���3�@��\S�3@�?t_��!?����@Q�#
�ٿ+���3�@��\S�3@�?t_��!?����@Q�#
�ٿ+���3�@��\S�3@�?t_��!?����@��h�ٿaq����@�@��`�3@r�AO��!?u� V�-�@1�^%��ٿN탪�	�@H���3@8�i�!?�'�j�!�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@͐5�ğٿ��)�4��@�mk��3@j囏�!?��Ԗ;�@f�uo��ٿ�`�e�@Z����3@��!?��U{�@f�uo��ٿ�`�e�@Z����3@��!?��U{�@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@Go"�2�ٿ]lC��@e*�V�3@�	S��!?K�"�Z��@+$�r�ٿ)�P%�@���:�3@����ߐ!?͊Qn<��@+$�r�ٿ)�P%�@���:�3@����ߐ!?͊Qn<��@+$�r�ٿ)�P%�@���:�3@����ߐ!?͊Qn<��@+$�r�ٿ)�P%�@���:�3@����ߐ!?͊Qn<��@+$�r�ٿ)�P%�@���:�3@����ߐ!?͊Qn<��@'s|��ٿ4�q٫��@����3@�Pխ��!?o�r����@�&�_�ٿ_'A��@���3@ezO��!?Y˵`-��@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@���J�ٿ�GG��@��Qۯ�3@D剂ѐ!?b�L+�@�z�-�ٿ�������@������3@=���֐!?G�!Xz��@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@O��/�ٿ�z\
�~�@y�����3@��+��!?�(�+�@sER�ٿ���F�@Z�Xg�3@!s*��!?�F���@��S���ٿO��P��@�����3@e���!?���x���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@�lѣ�ٿ��(eY��@k�I�K�3@rH��!?K�g���@m�1��ٿTb�U�o�@�-(e�3@}����!?Pr���	�@���tf�ٿAa!���@��?� �3@����Ő!?Bv��&��@���tf�ٿAa!���@��?� �3@����Ő!?Bv��&��@�,/e9�ٿn(�ժ��@=�&��3@3�2���!?�KuTo6�@�����ٿ�k����@D�֮��3@�0��!?B&]����@�����ٿ�k����@D�֮��3@�0��!?B&]����@ly??A�ٿl�\ک�@��=8�3@�����!? �ڨ���@ly??A�ٿl�\ک�@��=8�3@�����!? �ڨ���@ly??A�ٿl�\ک�@��=8�3@�����!? �ڨ���@ly??A�ٿl�\ک�@��=8�3@�����!? �ڨ���@��u��ٿ�S\Z���@��7��3@$c%�!?%��[���@ʰ�ꂝٿ���-��@�|E��3@n>�� �!?�d%���@ʰ�ꂝٿ���-��@�|E��3@n>�� �!?�d%���@ʰ�ꂝٿ���-��@�|E��3@n>�� �!?�d%���@ʰ�ꂝٿ���-��@�|E��3@n>�� �!?�d%���@ʰ�ꂝٿ���-��@�|E��3@n>�� �!?�d%���@��1H�ٿQ�ţ�C�@��"��3@��'�!?F��\���@��1H�ٿQ�ţ�C�@��"��3@��'�!?F��\���@��1H�ٿQ�ţ�C�@��"��3@��'�!?F��\���@��1H�ٿQ�ţ�C�@��"��3@��'�!?F��\���@&�~��ٿ�}�����@K�3�>�3@�3�A��!?Τ�O1T�@&�~��ٿ�}�����@K�3�>�3@�3�A��!?Τ�O1T�@&�~��ٿ�}�����@K�3�>�3@�3�A��!?Τ�O1T�@&�~��ٿ�}�����@K�3�>�3@�3�A��!?Τ�O1T�@d�T��ٿ�����@�KQ��3@s �w��!?L�3��N�@d�T��ٿ�����@�KQ��3@s �w��!?L�3��N�@d�T��ٿ�����@�KQ��3@s �w��!?L�3��N�@d�T��ٿ�����@�KQ��3@s �w��!?L�3��N�@]w�ٿ�hu����@`��&��3@K���!?�r����@]w�ٿ�hu����@`��&��3@K���!?�r����@]w�ٿ�hu����@`��&��3@K���!?�r����@Ϣ,n�ٿ6����@��_��3@NI��Ɛ!?��K�,�@Ϣ,n�ٿ6����@��_��3@NI��Ɛ!?��K�,�@Ϣ,n�ٿ6����@��_��3@NI��Ɛ!?��K�,�@Ϣ,n�ٿ6����@��_��3@NI��Ɛ!?��K�,�@Ϣ,n�ٿ6����@��_��3@NI��Ɛ!?��K�,�@9<�u�ٿ;E�iA�@<C܅��3@j� ��!?�l���@9<�u�ٿ;E�iA�@<C܅��3@j� ��!?�l���@9<�u�ٿ;E�iA�@<C܅��3@j� ��!?�l���@9<�u�ٿ;E�iA�@<C܅��3@j� ��!?�l���@9<�u�ٿ;E�iA�@<C܅��3@j� ��!?�l���@��d�ٿ��_K�@��JE��3@�bF��!?vS�s��@��d�ٿ��_K�@��JE��3@�bF��!?vS�s��@���F>�ٿS>@J��@�[g��3@��蚦�!?s ��S��@���F>�ٿS>@J��@�[g��3@��蚦�!?s ��S��@���F>�ٿS>@J��@�[g��3@��蚦�!?s ��S��@���F>�ٿS>@J��@�[g��3@��蚦�!?s ��S��@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@d��7ǘٿ��S�ʮ�@aڥ�3@QE1ې!?^ZYtW�@&����ٿjm3�QZ�@5Ap�M�3@�XL��!?���:��@�}�GI�ٿ뇙�E��@��Rʿ�3@`ۖ�!?h�����@�}�GI�ٿ뇙�E��@��Rʿ�3@`ۖ�!?h�����@v:|��ٿ��n���@��׫�3@L�����!?9u`!���@v:|��ٿ��n���@��׫�3@L�����!?9u`!���@v:|��ٿ��n���@��׫�3@L�����!?9u`!���@O��@�ٿa�]���@Ԋ�7H�3@��%B�!?gc	�
m�@O��@�ٿa�]���@Ԋ�7H�3@��%B�!?gc	�
m�@O��@�ٿa�]���@Ԋ�7H�3@��%B�!?gc	�
m�@�'W���ٿu��-��@[gP��3@ �x�
�!?F�5!�@ja�B�ٿc�x��]�@;���3@n��֐!?����$2�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@J$//�ٿE�p����@]�C���3@���	�!?���.?P�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@�A�m�ٿ��6[z��@��9�<�3@����!?��m�@ �-"��ٿ�c�q.�@'���3@.c�Ð!?��߲�	�@ �-"��ٿ�c�q.�@'���3@.c�Ð!?��߲�	�@E�`@�ٿd�Ù��@T��?��3@�2ǧ�!?)�n9E�@E�`@�ٿd�Ù��@T��?��3@�2ǧ�!?)�n9E�@E�`@�ٿd�Ù��@T��?��3@�2ǧ�!?)�n9E�@�q�ٿ�ڙz���@[��Ji�3@�Sᬐ!?l4�W��@�q�ٿ�ڙz���@[��Ji�3@�Sᬐ!?l4�W��@�q�ٿ�ڙz���@[��Ji�3@�Sᬐ!?l4�W��@��h��ٿ�n��J:�@7�[3\�3@�ʟ�Đ!?AI���@��h��ٿ�n��J:�@7�[3\�3@�ʟ�Đ!?AI���@��h��ٿ�n��J:�@7�[3\�3@�ʟ�Đ!?AI���@��h��ٿ�n��J:�@7�[3\�3@�ʟ�Đ!?AI���@_�)�!�ٿyg�+���@�����3@������!?�~��'��@_�)�!�ٿyg�+���@�����3@������!?�~��'��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@��։Ρٿv76���@���u�3@�:���!?�JB/|��@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�Oq��ٿ�Q9��@T*����3@�(W�!?��5Gv�@�RĔ��ٿ�U$�r=�@^u@��3@᩽��!?mG���@�RĔ��ٿ�U$�r=�@^u@��3@᩽��!?mG���@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@�k�4�ٿ��Y0���@lp-�3@�&��!?+�6�
o�@PC��ٿ<.�!��@~�U:��3@�*d�!?kcKU�O�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@�}�_m�ٿZL@��@�ѣ��3@��D2	�!?��:�Hg�@����æٿ:!�m8�@�_��F�3@Zus���!? �Щ^W�@z�#�S�ٿ���v	9�@�hr���3@���A��!?W�n�n�@z�#�S�ٿ���v	9�@�hr���3@���A��!?W�n�n�@z�#�S�ٿ���v	9�@�hr���3@���A��!?W�n�n�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@Z?��E�ٿ/Y:���@Ưdʎ�3@�z�oϐ!?�[��u�@���e��ٿw�p�i��@��ۤ�3@�R݂��!?2����@���e��ٿw�p�i��@��ۤ�3@�R݂��!?2����@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@f�)��ٿ����@�F���3@������!?Ѡ}���@������ٿ|������@�-k�\�3@*����!?ŗ�W���@������ٿ|������@�-k�\�3@*����!?ŗ�W���@��3R�ٿ�٪K�@:���1�3@y'��!?
�TD��@��3R�ٿ�٪K�@:���1�3@y'��!?
�TD��@r�$�ٿ\Qd��@�Z���3@Ͱ���!?�ǡ��L�@r�$�ٿ\Qd��@�Z���3@Ͱ���!?�ǡ��L�@i�0���ٿ�����	�@��j���3@?El5�!?0���@�y?�`�ٿ���4��@�0���3@�a��!?äO̵��@�y?�`�ٿ���4��@�0���3@�a��!?äO̵��@�y?�`�ٿ���4��@�0���3@�a��!?äO̵��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@-O
���ٿ������@&�|Y��3@����!?Sz�e��@|�b�ٿniR����@�5��3@����!?k�a0i��@|�b�ٿniR����@�5��3@����!?k�a0i��@|�b�ٿniR����@�5��3@����!?k�a0i��@|�b�ٿniR����@�5��3@����!?k�a0i��@0F���ٿ�*��ԅ�@�'�0�3@L2�ސ!?���C�:�@�ُz'�ٿ�H���@��I�y�3@��� �!?���B�@�ُz'�ٿ�H���@��I�y�3@��� �!?���B�@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@7�|�ٿ�+T�9�@o�Ɨm�3@o?����!? �����@��"s-�ٿ�GE%�@l�,j�3@�$?N��!?�ƎM]��@��"s-�ٿ�GE%�@l�,j�3@�$?N��!?�ƎM]��@��"s-�ٿ�GE%�@l�,j�3@�$?N��!?�ƎM]��@�W8/�ٿ
F c��@�;2��3@wE+�!?��q���@.�X��ٿ���M�@6d��3@��mC�!?��+��D�@.�X��ٿ���M�@6d��3@��mC�!?��+��D�@.�X��ٿ���M�@6d��3@��mC�!?��+��D�@.�X��ٿ���M�@6d��3@��mC�!?��+��D�@��E�ٿ7FF���@�H���3@	�r'�!?�����T�@��E�ٿ7FF���@�H���3@	�r'�!?�����T�@��E�ٿ7FF���@�H���3@	�r'�!?�����T�@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@�s�_��ٿZ�@�)��3@��>4�!?I-����@��v�ٿ^	a&H��@�Ƣ�3@Z�(g(�!?Z�+�g�@��v�ٿ^	a&H��@�Ƣ�3@Z�(g(�!?Z�+�g�@ ��f�ٿ�/��3��@Q�^M}�3@�/�5
�!?��>�$�@6|F��ٿ��C����@^���w�3@%���!?�*���@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@px��ٿ
*Z� �@e4����3@ܾ�㥐!?������@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@��եٿ�~W��@�è��3@6�M6��!?/1J�C�@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@?1�D�ٿF=�@W�@H�>L��3@t��)��!?1yݵ���@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�K�:��ٿ��jlߥ�@�Zt�D�3@^*�Bv�!?��'	d�@�#W��ٿJu�|g�@�Ɛ���3@<L�K�!?Ek�e��@�#W��ٿJu�|g�@�Ɛ���3@<L�K�!?Ek�e��@�#W��ٿJu�|g�@�Ɛ���3@<L�K�!?Ek�e��@�@��/�ٿ��[4��@����3@Q�[=�!?ܯ.L�y�@�AUp�ٿanB粢�@��$9�3@n���!?��ч.�@�AUp�ٿanB粢�@��$9�3@n���!?��ч.�@�H��ݢٿ��Р��@�"ǔ�3@[��ː!?���!�3�@�H��ݢٿ��Р��@�"ǔ�3@[��ː!?���!�3�@�H��ݢٿ��Р��@�"ǔ�3@[��ː!?���!�3�@�H��ݢٿ��Р��@�"ǔ�3@[��ː!?���!�3�@�H��ݢٿ��Р��@�"ǔ�3@[��ː!?���!�3�@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@D[}�h�ٿ�!�$ ��@��ɖ��3@\�cn�!?đk����@^�=��ٿ�;�ι��@o�)��3@�0A�֐!?�tp~�J�@^�=��ٿ�;�ι��@o�)��3@�0A�֐!?�tp~�J�@^�=��ٿ�;�ι��@o�)��3@�0A�֐!?�tp~�J�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@�̔��ٿ�-�6���@�-����3@��h���!?=o��Y�@Nu�-��ٿ ���M�@�j�q�3@��L��!?����/��@Nu�-��ٿ ���M�@�j�q�3@��L��!?����/��@Nu�-��ٿ ���M�@�j�q�3@��L��!?����/��@Nu�-��ٿ ���M�@�j�q�3@��L��!?����/��@�+����ٿ�P�Ť��@L9����3@�qB<Ő!?*T���@ Q��ߥٿ=�Wp�@�)���3@h��è�!?�HY�Y��@ Q��ߥٿ=�Wp�@�)���3@h��è�!?�HY�Y��@ Q��ߥٿ=�Wp�@�)���3@h��è�!?�HY�Y��@ Q��ߥٿ=�Wp�@�)���3@h��è�!?�HY�Y��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�)����ٿ*C���@ٯn|�3@�/Ʉ�!?��k��@�É=��ٿۿ��(�@�J�$�3@O*ʌ�!?��*�v��@�É=��ٿۿ��(�@�J�$�3@O*ʌ�!?��*�v��@�É=��ٿۿ��(�@�J�$�3@O*ʌ�!?��*�v��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@R����ٿ�QQT��@�\���3@t�T�!?���.��@w��K�ٿߝ��W3�@����2�3@��'��!?H�	�l�@w��K�ٿߝ��W3�@����2�3@��'��!?H�	�l�@w��K�ٿߝ��W3�@����2�3@��'��!?H�	�l�@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@��$��ٿO�ǅZ�@�y6���3@H�}埐!?vddC���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@x���	�ٿ2�i5�@A���
�3@�M�Đ!?�kH���@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@9�YΡٿi�f)��@�(���3@�P�+ΐ!?��W����@�}����ٿ�	b���@�"V��3@T�ʐ!?����@�}����ٿ�	b���@�"V��3@T�ʐ!?����@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@�c|��ٿ���K|��@:��'��3@�����!?�x��/�@~�hS�ٿ�9����@�$C7�3@}5b�Ӑ!?µ,!3,�@,�n�9�ٿ������@qbU���3@|Ϸ*��!?�f�Uz�@,�n�9�ٿ������@qbU���3@|Ϸ*��!?�f�Uz�@�ͅ
�ٿ|��k ��@<cFȬ�3@wzH�z�!?	���)��@{|F�Τٿ�"���@�Q?؊�3@�q1a��!?y�k�ˁ�@c�;<ŠٿD!�f2w�@�%��p�3@*�?�Ɛ!?��@�~A�@c�;<ŠٿD!�f2w�@�%��p�3@*�?�Ɛ!?��@�~A�@<+�ɣٿx� �~�@d���4�3@�fX�Ð!?�-����@<+�ɣٿx� �~�@d���4�3@�fX�Ð!?�-����@)�k��ٿ�
�Y�s�@����3@��~�Z�!?@�F�j��@)�k��ٿ�
�Y�s�@����3@��~�Z�!?@�F�j��@;��b�ٿM����@��~�^�3@0��%�!?q��q{�@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@�n4�ٿʄN��@��듎�3@ ��!?7�
G��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@6<�֞ٿ��T����@� ��3@��!�!?��ϡ]��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��(h=�ٿ���gY|�@r`a8��3@���"��!?rE�@��@��B�ٿ�"0
��@��,w��3@�c)��!?��aK��@��B�ٿ�"0
��@��,w��3@�c)��!?��aK��@��B�ٿ�"0
��@��,w��3@�c)��!?��aK��@��B�ٿ�"0
��@��,w��3@�c)��!?��aK��@0�};�ٿSSuW��@���9��3@�a���!?V�d���@0�};�ٿSSuW��@���9��3@�a���!?V�d���@0�};�ٿSSuW��@���9��3@�a���!?V�d���@0�};�ٿSSuW��@���9��3@�a���!?V�d���@0�};�ٿSSuW��@���9��3@�a���!?V�d���@0�};�ٿSSuW��@���9��3@�a���!?V�d���@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@�C��K�ٿZ������@�U���3@�-���!?�"Eǀ�@ʑ�7�ٿ����>�@~Wk8�3@�-�u�!?04���T�@���cٜٿ�^�O�@)?s�3@I�2h��!? S-}F��@���cٜٿ�^�O�@)?s�3@I�2h��!? S-}F��@���cٜٿ�^�O�@)?s�3@I�2h��!? S-}F��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@�H��!�ٿ��EU�@W�Н�3@བ�!?���u��@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@;o9�w�ٿ�I�����@d,N�3�3@:�bƔ�!?���_g@�@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@9�bڰ�ٿz����@�e����3@��*��!?��L ���@!�HŢٿs��~��@ A����3@9��!?:5��CM�@!�HŢٿs��~��@ A����3@9��!?:5��CM�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@�]Kjڠٿ���ĺ�@�d��3@��Q��!?��Z�l�@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@څI��ٿ��^m��@L�`>B�3@��>|�!?�����@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@���A�ٿ�9/<��@�`B���3@_ه6��!?p+��_��@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@9\�J�ٿ�x���@N����3@j2��̐!?>� �t �@�B<���ٿo��=��@�Gw�M�3@9�Q��!?	Șd@|�@�B<���ٿo��=��@�Gw�M�3@9�Q��!?	Șd@|�@uieXS�ٿ���E��@��"�^�3@:;k��!?XJ�&%�@uieXS�ٿ���E��@��"�^�3@:;k��!?XJ�&%�@����ٝٿ#Ρ�*��@ex��3@8���ɐ!?��X�@�@����ٝٿ#Ρ�*��@ex��3@8���ɐ!?��X�@�@����ٝٿ#Ρ�*��@ex��3@8���ɐ!?��X�@�@\��A�ٿ?B�N2��@�"֌6�3@�O�)!?��TR��@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@�{Ɏ��ٿH���$��@�v�	�3@����u�!?%s�����@l�tW��ٿ�_,\�`�@D���3@�_���!?�����@O�)�r�ٿ�Z*�2�@��c��3@Rҗ ��!?(��?�@O�)�r�ٿ�Z*�2�@��c��3@Rҗ ��!?(��?�@O�)�r�ٿ�Z*�2�@��c��3@Rҗ ��!?(��?�@O�)�r�ٿ�Z*�2�@��c��3@Rҗ ��!?(��?�@O�)�r�ٿ�Z*�2�@��c��3@Rҗ ��!?(��?�@է +��ٿo�2�,�@,��3@�����!?崤�.y�@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�k���ٿ�j*u{�@Q+�ƿ�3@�^"v��!?$i=U���@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@�L#��ٿ�{� ]�@ؑaM��3@�ñ>��!?�P�&�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@>d=ѠٿA�An�N�@����3@�~v�0�!?�����W�@��J�.�ٿR��ù�@�B���3@�g�x�!?ʿ��8��@���)�ٿ�8�39��@�pp��3@E���֐!?I��4��@���)�ٿ�8�39��@�pp��3@E���֐!?I��4��@���-�ٿ�2��jA�@��g��3@�͝ǐ!?�Ѵ�_E�@���-�ٿ�2��jA�@��g��3@�͝ǐ!?�Ѵ�_E�@w�� �ٿJ�A��^�@j31�R�3@�@���!?�K�TV�@w�� �ٿJ�A��^�@j31�R�3@�@���!?�K�TV�@w�� �ٿJ�A��^�@j31�R�3@�@���!?�K�TV�@w�� �ٿJ�A��^�@j31�R�3@�@���!?�K�TV�@%;׶��ٿG����@�?�f��3@_��K��!?e�M��@%;׶��ٿG����@�?�f��3@_��K��!?e�M��@%;׶��ٿG����@�?�f��3@_��K��!?e�M��@%;׶��ٿG����@�?�f��3@_��K��!?e�M��@%;׶��ٿG����@�?�f��3@_��K��!?e�M��@-!m���ٿ�T�?�=�@�' fa�3@x�Ѹ�!?�|��L�@-!m���ٿ�T�?�=�@�' fa�3@x�Ѹ�!?�|��L�@-!m���ٿ�T�?�=�@�' fa�3@x�Ѹ�!?�|��L�@$����ٿ��g��@>h�3@0��� �!?X�"fD�@���O�ٿT��y��@�����3@�
���!?���a��@��O�ߜٿ�e�Տ�@�l���3@�%,�!?�7\�΢�@��O�ߜٿ�e�Տ�@�l���3@�%,�!?�7\�΢�@��O�ߜٿ�e�Տ�@�l���3@�%,�!?�7\�΢�@��O�ߜٿ�e�Տ�@�l���3@�%,�!?�7\�΢�@��O�ߜٿ�e�Տ�@�l���3@�%,�!?�7\�΢�@]�e�@�ٿ��QX�3�@�h�o�3@20���!?�u����@]�e�@�ٿ��QX�3�@�h�o�3@20���!?�u����@]�e�@�ٿ��QX�3�@�h�o�3@20���!?�u����@}cF��ٿ�W	����@�����3@�\F��!?����<�@}cF��ٿ�W	����@�����3@�\F��!?����<�@}cF��ٿ�W	����@�����3@�\F��!?����<�@}cF��ٿ�W	����@�����3@�\F��!?����<�@}cF��ٿ�W	����@�����3@�\F��!?����<�@���ٿy]����@G��*�3@�:�ֹ�!?�.�x��@���{��ٿK��j��@zJ���3@F�&2Ɛ!?�����@�=1ɚٿ�4�ً��@&{%D�3@���!?�=���n�@�=1ɚٿ�4�ً��@&{%D�3@���!?�=���n�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@2���o�ٿr��#���@.�5�3@H�Bi!?�_.R	�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@B��[��ٿO��nM$�@F����3@��qu�!?e.bt�@�HK�ٿ���.A�@��F���3@�3:�!?L	ߥ��@">̖q�ٿm2V\N�@�B����3@P�թ�!?1�v��>�@">̖q�ٿm2V\N�@�B����3@P�թ�!?1�v��>�@">̖q�ٿm2V\N�@�B����3@P�թ�!?1�v��>�@">̖q�ٿm2V\N�@�B����3@P�թ�!?1�v��>�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@�M����ٿ��N���@�"RJ�3@-/�{�!?� �$�@#yw���ٿ��}0���@��|��3@���\�!?�
p� ��@#yw���ٿ��}0���@��|��3@���\�!?�
p� ��@��~���ٿ�,e3n�@�n����3@KlQא!?�����Q�@��~���ٿ�,e3n�@�n����3@KlQא!?�����Q�@��~���ٿ�,e3n�@�n����3@KlQא!?�����Q�@Y2�$�ٿ*\g�m�@��:D�3@�>����!?i�Y��@Y2�$�ٿ*\g�m�@��:D�3@�>����!?i�Y��@Y2�$�ٿ*\g�m�@��:D�3@�>����!?i�Y��@Y2�$�ٿ*\g�m�@��:D�3@�>����!?i�Y��@Y2�$�ٿ*\g�m�@��:D�3@�>����!?i�Y��@�� �ٿD*��v�@A�!��3@�N���!?<��'V��@�� �ٿD*��v�@A�!��3@�N���!?<��'V��@�� �ٿD*��v�@A�!��3@�N���!?<��'V��@��@�ٿST�t��@��+6�3@�`���!?s@�6F�@��@�ٿST�t��@��+6�3@�`���!?s@�6F�@���3L�ٿK��g�]�@��1�r�3@�+�9��!?%b�*X�@���3L�ٿK��g�]�@��1�r�3@�+�9��!?%b�*X�@���3L�ٿK��g�]�@��1�r�3@�+�9��!?%b�*X�@���3L�ٿK��g�]�@��1�r�3@�+�9��!?%b�*X�@��򠪜ٿ-M���@ 4�B�3@��p�!?��\�@��򠪜ٿ-M���@ 4�B�3@��p�!?��\�@��򠪜ٿ-M���@ 4�B�3@��p�!?��\�@��򠪜ٿ-M���@ 4�B�3@��p�!?��\�@��򠪜ٿ-M���@ 4�B�3@��p�!?��\�@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@ۛ�I�ٿ\�,�K��@� ��,�3@�6�W��!?�o�j���@K�����ٿ��F��@��)�h�3@瓇ڐ!?d˅H/�@K�����ٿ��F��@��)�h�3@瓇ڐ!?d˅H/�@K�����ٿ��F��@��)�h�3@瓇ڐ!?d˅H/�@K�����ٿ��F��@��)�h�3@瓇ڐ!?d˅H/�@K�����ٿ��F��@��)�h�3@瓇ڐ!?d˅H/�@(b��ţٿ��^���@:ֆ�3@��N&;�!?��)]i��@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@m}��m�ٿv��`��@�c��H�3@8y�&;�!?${�\i�@ DUX�ٿu�X1�@�f�*��3@?�켻�!?�{�/�@ DUX�ٿu�X1�@�f�*��3@?�켻�!?�{�/�@ DUX�ٿu�X1�@�f�*��3@?�켻�!?�{�/�@ DUX�ٿu�X1�@�f�*��3@?�켻�!?�{�/�@Х揜ٿ��K��o�@`�"�I�3@Rc�P��!?��7����@I9C?�ٿ-�X9�i�@�����3@l�t�!?2:�[���@�ޚ�_�ٿ1�d��(�@��O��3@e��ͽ�!?�Ot���@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@�A%��ٿ��:��<�@���3@@C��!?�!f ˄�@��Q�ٿ�W�f0%�@�Y��3@���8͐!?�m�P�&�@��Q�ٿ�W�f0%�@�Y��3@���8͐!?�m�P�&�@���ٿ��LW��@��d�3@��i���!?g����W�@���ٿ��LW��@��d�3@��i���!?g����W�@���ٿ��LW��@��d�3@��i���!?g����W�@���ٿ��LW��@��d�3@��i���!?g����W�@���ٿ��LW��@��d�3@��i���!?g����W�@���
x�ٿ�/7h,�@�S�3@\����!?����@�ou�|�ٿd�b#s�@cOO��3@����!?z��yC�@CO>��ٿX��@�F-��3@:��_��!?�����^�@CO>��ٿX��@�F-��3@:��_��!?�����^�@CO>��ٿX��@�F-��3@:��_��!?�����^�@CO>��ٿX��@�F-��3@:��_��!?�����^�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@�J1X�ٿƷ�,�@�@"�3@��pт�!?�z��.]�@������ٿɆz�P�@�cٶ��3@?#hƐ!?)�\
[�@<��ٿyȇ�T�@Tv{^��3@4�e��!?O�S"!x�@<��ٿyȇ�T�@Tv{^��3@4�e��!?O�S"!x�@��/��ٿ�i��q��@U�3��3@=�!?�uB�@��/��ٿ�i��q��@U�3��3@=�!?�uB�@��/��ٿ�i��q��@U�3��3@=�!?�uB�@��/��ٿ�i��q��@U�3��3@=�!?�uB�@Ֆ]P�ٿ��?� ��@��P9��3@��}�!?��ZKư�@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@ �o�ٿ��3$�@�+��3@�v׽f�!?�=`�(��@}�"�w�ٿ�,�Z��@c����3@���ꡐ!?"L���S�@�o���ٿ�4����@����3@u���!?�M�=uI�@�o���ٿ�4����@����3@u���!?�M�=uI�@�o���ٿ�4����@����3@u���!?�M�=uI�@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@Z��e�ٿm{�k��@m�f<�3@Q=2�!?m5�̧��@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@�[�R�ٿ���X�q�@�2h�v�3@���>��!?<ܷY[�@���ٿ�0����@�l5v}�3@+v&��!?dq���[�@eZ�ti�ٿ�
��R��@8d�۟�3@KY��!?sc����@eZ�ti�ٿ�
��R��@8d�۟�3@KY��!?sc����@eZ�ti�ٿ�
��R��@8d�۟�3@KY��!?sc����@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@�'��ٿ}���P��@		��3@�x��!?�* >��@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@� �ߞٿkÉ��@{Y^��3@`ea4�!?ڒW��z�@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@�bs;�ٿ2��"��@ ����3@-�؉�!?; ���@���]��ٿV��IU��@�L-�=�3@գ[���!?��P��@���]��ٿV��IU��@�L-�=�3@գ[���!?��P��@���]��ٿV��IU��@�L-�=�3@գ[���!?��P��@���]��ٿV��IU��@�L-�=�3@գ[���!?��P��@$��2�ٿ�B��p�@ʼ���3@4��ʲ�!?��SU��@$��2�ٿ�B��p�@ʼ���3@4��ʲ�!?��SU��@߿�5�ٿ4����@&�����3@�K���!?�2;~��@߿�5�ٿ4����@&�����3@�K���!?�2;~��@e'���ٿ��t��M�@�0E���3@'�n5�!?��G����@e'���ٿ��t��M�@�0E���3@'�n5�!?��G����@e'���ٿ��t��M�@�0E���3@'�n5�!?��G����@e'���ٿ��t��M�@�0E���3@'�n5�!?��G����@e'���ٿ��t��M�@�0E���3@'�n5�!?��G����@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@ꅱAٿ"�@�'�%��3@�V���!?6;:�
�@=E�#��ٿO����@3<"~�3@�$��!?)����@=E�#��ٿO����@3<"~�3@�$��!?)����@*Y�Sw�ٿ ����}�@��Q���3@�J��!?���WJ�@*Y�Sw�ٿ ����}�@��Q���3@�J��!?���WJ�@*Y�Sw�ٿ ����}�@��Q���3@�J��!?���WJ�@*Y�Sw�ٿ ����}�@��Q���3@�J��!?���WJ�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@N�m�f�ٿv��u��@ �n{��3@׷rؐ!?��P_?>�@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@üa���ٿQƷY
��@xKx���3@}%ݐ!?��`���@�ק�7�ٿ�B�3�@�)�3@j^�Ő!?a��#Q�@�ק�7�ٿ�B�3�@�)�3@j^�Ő!?a��#Q�@�ק�7�ٿ�B�3�@�)�3@j^�Ő!?a��#Q�@�ק�7�ٿ�B�3�@�)�3@j^�Ő!?a��#Q�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@�c���ٿ"��v�@�:�Y�3@P!��w�!?i�)�e�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@_I>�k�ٿ|02�P�@Hw*��3@$ܫ8��!?6��Z�0�@�J-��ٿ���Oq�@_��x��3@�f�ϋ�!?E:E�Z�@�J-��ٿ���Oq�@_��x��3@�f�ϋ�!?E:E�Z�@�J-��ٿ���Oq�@_��x��3@�f�ϋ�!?E:E�Z�@���(��ٿ}FK���@w��I	�3@_����!?��D�J��@{���ٿ�c����@dO\[�3@�+ER֐!?PQ��g�@{���ٿ�c����@dO\[�3@�+ER֐!?PQ��g�@�И,�ٿ��,	&�@?�?���3@�����!?6�K�q�@�И,�ٿ��,	&�@?�?���3@�����!?6�K�q�@�И,�ٿ��,	&�@?�?���3@�����!?6�K�q�@��Ϛٿ=*� ��@j\Tn��3@��Fʐ!?���w�@"�(h��ٿ�a���@l��|d�3@u6�)c�!?ɪ�':�@"�(h��ٿ�a���@l��|d�3@u6�)c�!?ɪ�':�@!�&��ٿ7���F�@b�C�3@��P��!?J�{�jL�@b\@y��ٿ<�����@n���Y�3@�l�!?="a{��@b\@y��ٿ<�����@n���Y�3@�l�!?="a{��@b\@y��ٿ<�����@n���Y�3@�l�!?="a{��@b\@y��ٿ<�����@n���Y�3@�l�!?="a{��@��
l��ٿ,�lb�@�����3@�,Z�!?�R�`���@�ī$�ٿ��&6��@$�����3@��ΐ!?���#�@�ī$�ٿ��&6��@$�����3@��ΐ!?���#�@�E"}�ٿ�Gw]���@�0}>��3@��v?%�!?L��X���@f�`	�ٿؼjۭ�@<^���3@~���!?]1��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@��x�~�ٿ��P�d��@y��*��3@��⺐!?U�e��@"�)c��ٿ~
w�f�@�jb6�3@''�ې!?s�MYI��@"�)c��ٿ~
w�f�@�jb6�3@''�ې!?s�MYI��@����ٿ䲴�K�@��<�3@c���ِ!?�;��o}�@GQ@�ٿ��i��@Z���o�3@��;���!?�uv5v�@GQ@�ٿ��i��@Z���o�3@��;���!?�uv5v�@GQ@�ٿ��i��@Z���o�3@��;���!?�uv5v�@GQ@�ٿ��i��@Z���o�3@��;���!?�uv5v�@�����ٿm�_�6�@V-�B�3@�����!?9w�;Zm�@���ٿh�5>��@��.���3@-��K͐!?TgS�q��@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@�4�[�ٿ���;K�@�b��3�3@�謐!?�]?CI�@����E�ٿ��<���@'�<��3@�O���!?b��n�@����E�ٿ��<���@'�<��3@�O���!?b��n�@����E�ٿ��<���@'�<��3@�O���!?b��n�@����E�ٿ��<���@'�<��3@�O���!?b��n�@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@B�?Md�ٿK�%2��@�u���3@E9�#�!?��^���@P�r���ٿQ��t��@�imE��3@σc�'�!?��35�Z�@P�r���ٿQ��t��@�imE��3@σc�'�!?��35�Z�@��A֡�ٿ;��6��@ތ���3@Ҹ�⹐!?�Sr��B�@��A֡�ٿ;��6��@ތ���3@Ҹ�⹐!?�Sr��B�@��A֡�ٿ;��6��@ތ���3@Ҹ�⹐!?�Sr��B�@��A֡�ٿ;��6��@ތ���3@Ҹ�⹐!?�Sr��B�@�|'x�ٿk����O�@A<�2�3@����!?�8����@�|'x�ٿk����O�@A<�2�3@����!?�8����@�|'x�ٿk����O�@A<�2�3@����!?�8����@�|'x�ٿk����O�@A<�2�3@����!?�8����@H�p�ٿ.tO/�@���*:�3@o�u!R�!?�h����@H�p�ٿ.tO/�@���*:�3@o�u!R�!?�h����@��l��ٿ�>���@�П���3@�ӣw^�!?}��~,�@��l��ٿ�>���@�П���3@�ӣw^�!?}��~,�@��l��ٿ�>���@�П���3@�ӣw^�!?}��~,�@��b.�ٿ��#���@��q;��3@�J�p�!?d�3aL��@��b.�ٿ��#���@��q;��3@�J�p�!?d�3aL��@��b.�ٿ��#���@��q;��3@�J�p�!?d�3aL��@��b.�ٿ��#���@��q;��3@�J�p�!?d�3aL��@��b.�ٿ��#���@��q;��3@�J�p�!?d�3aL��@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��Sc�ٿz9'���@�D>�i�3@�@=���!?�XH�@��,ҵ�ٿ���ƭ=�@�%[5��3@�FSC�!?���Q��@��,ҵ�ٿ���ƭ=�@�%[5��3@�FSC�!?���Q��@�n�m^�ٿv��l�@���bm�3@J���ǐ!?I����@�n�m^�ٿv��l�@���bm�3@J���ǐ!?I����@�n�m^�ٿv��l�@���bm�3@J���ǐ!?I����@�n�m^�ٿv��l�@���bm�3@J���ǐ!?I����@�4C���ٿPPo=]��@ż 5��3@���4֐!?�@)2��@4)�{�ٿ�1�:O��@��{�r�3@��Qoʐ!?���?F�@4)�{�ٿ�1�:O��@��{�r�3@��Qoʐ!?���?F�@4)�{�ٿ�1�:O��@��{�r�3@��Qoʐ!?���?F�@4)�{�ٿ�1�:O��@��{�r�3@��Qoʐ!?���?F�@4)�{�ٿ�1�:O��@��{�r�3@��Qoʐ!?���?F�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@��F��ٿ!O�_rE�@eՊ���3@�N�)�!?8�se�@}�-L�ٿ~x�
�@@�˷�3@3}ah��!?�r���@}�-L�ٿ~x�
�@@�˷�3@3}ah��!?�r���@}�-L�ٿ~x�
�@@�˷�3@3}ah��!?�r���@�����ٿ����@MG*x��3@�̀���!?���f�0�@�����ٿ����@MG*x��3@�̀���!?���f�0�@�����ٿ����@MG*x��3@�̀���!?���f�0�@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@�e� �ٿ��_�Ϟ�@uG<��3@k~�e��!?����@|��&�ٿ���	U�@����3@���!?I,����@|��&�ٿ���	U�@����3@���!?I,����@|��&�ٿ���	U�@����3@���!?I,����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@ ��¡ٿ<<����@*<�!��3@pi-噐!?�+|����@0�r�ٿ2i�x��@�M�:�3@i����!?[���0��@>��+٠ٿp�~�/�@A�L/J�3@SP�7��!?���̱��@>��+٠ٿp�~�/�@A�L/J�3@SP�7��!?���̱��@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@�7(��ٿ]|
��@6��3�3@�/�+Ő!?F6����@{?�_��ٿ)f.!��@J���5�3@�m	�ǐ!?�.]y6��@{?�_��ٿ)f.!��@J���5�3@�m	�ǐ!?�.]y6��@{?�_��ٿ)f.!��@J���5�3@�m	�ǐ!?�.]y6��@{?�_��ٿ)f.!��@J���5�3@�m	�ǐ!?�.]y6��@\x�OУٿ'�;���@Z��+��3@��&k��!?����	��@\x�OУٿ'�;���@Z��+��3@��&k��!?����	��@\x�OУٿ'�;���@Z��+��3@��&k��!?����	��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@���ܣٿu5�ԅ�@D��>�3@O5e��!?�%�t��@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@�P)m|�ٿ6i��w�@�v-?�3@-�����!?��pdXV�@te��Ѣٿ���ո?�@��Tć�3@{nZf��!?v�Â��@te��Ѣٿ���ո?�@��Tć�3@{nZf��!?v�Â��@�B��ٿ�O�,1�@RPGK��3@�7`V�!?
�(e��@�B��ٿ�O�,1�@RPGK��3@�7`V�!?
�(e��@�B��ٿ�O�,1�@RPGK��3@�7`V�!?
�(e��@�B��ٿ�O�,1�@RPGK��3@�7`V�!?
�(e��@�B��ٿ�O�,1�@RPGK��3@�7`V�!?
�(e��@H�ʧٿF�{g_�@'!S3��3@�_
���!?��Ԙh��@H�ʧٿF�{g_�@'!S3��3@�_
���!?��Ԙh��@{`����ٿ�.>-���@���3@���!?�8ί�@{`����ٿ�.>-���@���3@���!?�8ί�@{`����ٿ�.>-���@���3@���!?�8ί�@{`����ٿ�.>-���@���3@���!?�8ί�@��'�ٿtF��;.�@��O��3@B�&@��!?G�j^�@��'�ٿtF��;.�@��O��3@B�&@��!?G�j^�@��'�ٿtF��;.�@��O��3@B�&@��!?G�j^�@LH���ٿ.�0�@b��@�3@e
Y4Ȑ!?X<Z_��@LH���ٿ.�0�@b��@�3@e
Y4Ȑ!?X<Z_��@�'�&0�ٿӉy���@�P���3@$��G�!?�Z�Y�A�@[d-��ٿR��*��@~cj��3@� ܆��!?lof�Nc�@[d-��ٿR��*��@~cj��3@� ܆��!?lof�Nc�@[d-��ٿR��*��@~cj��3@� ܆��!?lof�Nc�@[d-��ٿR��*��@~cj��3@� ܆��!?lof�Nc�@[d-��ٿR��*��@~cj��3@� ܆��!?lof�Nc�@��o�ٿ�ݭ�9�@�Ķ�3@^��ɐ!?MG?'.��@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@�!��ٿN��h��@'Ή���3@���ؐ�!?B}E>l�@����ٿ����@p�#M�3@�9��n�!?��:�,J�@����ٿ����@p�#M�3@�9��n�!?��:�,J�@����ٿ����@p�#M�3@�9��n�!?��:�,J�@6���A�ٿ]�#�0�@Dk���3@���w��!?zq�o�@�Ώ�x�ٿ�H�r��@��]�3@i��n�!?1M��@�Ώ�x�ٿ�H�r��@��]�3@i��n�!?1M��@{T��G�ٿ�����@��)�3@������!?�m-��@{T��G�ٿ�����@��)�3@������!?�m-��@�Ϧ��ٿj�*g�F�@��E���3@�PU46�!?�;�g5�@�Ϧ��ٿj�*g�F�@��E���3@�PU46�!?�;�g5�@�Ϧ��ٿj�*g�F�@��E���3@�PU46�!?�;�g5�@�圙I�ٿ0�
ש�@�tF{��3@����!?�&s��<�@�圙I�ٿ0�
ש�@�tF{��3@����!?�&s��<�@�圙I�ٿ0�
ש�@�tF{��3@����!?�&s��<�@��d��ٿο���@`����3@`TzNݐ!?tB��uZ�@��d��ٿο���@`����3@`TzNݐ!?tB��uZ�@��d��ٿο���@`����3@`TzNݐ!?tB��uZ�@��d��ٿο���@`����3@`TzNݐ!?tB��uZ�@��d��ٿο���@`����3@`TzNݐ!?tB��uZ�@Mq���ٿ�.�g�@"-����3@A����!?x��a]�@Mq���ٿ�.�g�@"-����3@A����!?x��a]�@Mq���ٿ�.�g�@"-����3@A����!?x��a]�@UrV`��ٿz���.�@NȁQ��3@<���+�!?����tW�@UrV`��ٿz���.�@NȁQ��3@<���+�!?����tW�@UrV`��ٿz���.�@NȁQ��3@<���+�!?����tW�@UrV`��ٿz���.�@NȁQ��3@<���+�!?����tW�@UrV`��ٿz���.�@NȁQ��3@<���+�!?����tW�@_���Y�ٿ�P�+R��@b�'�k�3@�Kl���!?�e��@�@_���Y�ٿ�P�+R��@b�'�k�3@�Kl���!?�e��@�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�%yϝٿ`�`�{�@ϋUi�3@i�t��!?(pLŽ�@�6�:^�ٿTӷ��@�[
H��3@%�ߐ!?�N`��
�@������ٿ�1���@�ذF��3@����!?6Xғ��@���ٿ�+��@�!c��3@�o?��!?Y'߅)��@���ٿ�+��@�!c��3@�o?��!?Y'߅)��@���ٿ�+��@�!c��3@�o?��!?Y'߅)��@���ٿ�+��@�!c��3@�o?��!?Y'߅)��@Q}�RM�ٿ>~<]�@�t�c��3@	�!�!?Ӛ�q$��@Q}�RM�ٿ>~<]�@�t�c��3@	�!�!?Ӛ�q$��@g�<��ٿ�ƍZ*��@J�#��3@w��~�!?]�m&Ah�@U_V�ٿ���_D�@h�G�q�3@��Uܐ!?�`YA��@�g�R�ٿO�).*[�@^�#��3@X���!?��ןJ�@�g�R�ٿO�).*[�@^�#��3@X���!?��ןJ�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@��K��ٿmNk��@;M�ϑ�3@�I�cА!?A��r]8�@L�0ǡٿ��b�|b�@+<�z�3@�^%��!?|i��o�@��у�ٿ�KL����@��O�E�3@�bZ=��!?;�ߛ�u�@*U��9�ٿ�+̆�n�@�Y�k��3@���C��!?=2�Th��@*U��9�ٿ�+̆�n�@�Y�k��3@���C��!?=2�Th��@*U��9�ٿ�+̆�n�@�Y�k��3@���C��!?=2�Th��@*U��9�ٿ�+̆�n�@�Y�k��3@���C��!?=2�Th��@: ��ϥٿ��Ө��@�* #w�3@`|#��!?{o0u��@: ��ϥٿ��Ө��@�* #w�3@`|#��!?{o0u��@: ��ϥٿ��Ө��@�* #w�3@`|#��!?{o0u��@: ��ϥٿ��Ө��@�* #w�3@`|#��!?{o0u��@�;���ٿ��ͱ���@��J�B�3@�2�oʐ!?Z�HB%V�@�;���ٿ��ͱ���@��J�B�3@�2�oʐ!?Z�HB%V�@�;���ٿ��ͱ���@��J�B�3@�2�oʐ!?Z�HB%V�@�;���ٿ��ͱ���@��J�B�3@�2�oʐ!?Z�HB%V�@Q(�3�ٿN����@Q{�" �3@D{_!?Г��mP�@Q(�3�ٿN����@Q{�" �3@D{_!?Г��mP�@WY��ٿL1�����@�k�2�3@�7XY�!?U,s=�@UW��ٿ�J�=���@Y`1"��3@y�P˕�!?·	��d�@eڂ˞�ٿ+�ɱ(Q�@t��f�3@�'��[�!?��V)�@eڂ˞�ٿ+�ɱ(Q�@t��f�3@�'��[�!?��V)�@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@{~�ġٿ+$E���@MJ2�S�3@�@9���!?������@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�fU0�ٿV_�]��@�ѽ$��3@ds��!?�U���@�ԩ�ٿ��Wxq�@��n�3@��-���!?N~!m ��@�ԩ�ٿ��Wxq�@��n�3@��-���!?N~!m ��@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@u��LۣٿE���&I�@X^-H��3@JJj��!?]�=���@�B���ٿ�-��T��@K�����3@W,G��!?�vn���@�B���ٿ�-��T��@K�����3@W,G��!?�vn���@�B���ٿ�-��T��@K�����3@W,G��!?�vn���@�B���ٿ�-��T��@K�����3@W,G��!?�vn���@�B���ٿ�-��T��@K�����3@W,G��!?�vn���@/-V~��ٿ���[8��@]����3@�H�/��!?$Ä�e�@/-V~��ٿ���[8��@]����3@�H�/��!?$Ä�e�@/-V~��ٿ���[8��@]����3@�H�/��!?$Ä�e�@/-V~��ٿ���[8��@]����3@�H�/��!?$Ä�e�@�Vw]�ٿ��/B�P�@�,���3@�F�-��!?0!7��@�Vw]�ٿ��/B�P�@�,���3@�F�-��!?0!7��@�Vw]�ٿ��/B�P�@�,���3@�F�-��!?0!7��@�Vw]�ٿ��/B�P�@�,���3@�F�-��!?0!7��@��%�ٿΒu����@�F��3@��Ր!?Ԭ<tI�@��%�ٿΒu����@�F��3@��Ր!?Ԭ<tI�@�%�$��ٿ7/	��,�@4��� 4@KG�*��!?I�R����@�%�$��ٿ7/	��,�@4��� 4@KG�*��!?I�R����@�%�$��ٿ7/	��,�@4��� 4@KG�*��!?I�R����@=O�0h�ٿ�-����@�>/��3@d�����!?�o:fT�@=O�0h�ٿ�-����@�>/��3@d�����!?�o:fT�@{����ٿ�׳�3�@U�=��3@Mx��!?��H�u1�@{����ٿ�׳�3�@U�=��3@Mx��!?��H�u1�@h8�͠ٿ���i�@1!���3@Ȅ��֐!?V�4h�I�@h@I�ٿ%:w�IM�@~9S��3@�+F[��!?�r�S�@h@I�ٿ%:w�IM�@~9S��3@�+F[��!?�r�S�@h@I�ٿ%:w�IM�@~9S��3@�+F[��!?�r�S�@&�Ľ�ٿ]b�ц�@=��� �3@l�ށ}�!?jt��_�@�v�a6�ٿ���K��@s���h�3@�h��!? :���T�@fҵ��ٿ��dsǊ�@S'���3@c��&�!?�*ƣ��@fҵ��ٿ��dsǊ�@S'���3@c��&�!?�*ƣ��@fҵ��ٿ��dsǊ�@S'���3@c��&�!?�*ƣ��@fҵ��ٿ��dsǊ�@S'���3@c��&�!?�*ƣ��@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@�AH�'�ٿ��NEc�@��p���3@��X4��!?�*�A���@M�#��ٿ�cQؤ��@�8�J�3@v����!?`��� ��@M�#��ٿ�cQؤ��@�8�J�3@v����!?`��� ��@M�#��ٿ�cQؤ��@�8�J�3@v����!?`��� ��@M�#��ٿ�cQؤ��@�8�J�3@v����!?`��� ��@M�#��ٿ�cQؤ��@�8�J�3@v����!?`��� ��@�� ��ٿ�L9��e�@C�i��3@�Zۘ�!?�`�D��@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Ϳo�Ϝٿ��W��@�~�S��3@b^nX��!?a�Z�$�@Y%���ٿ4�ǜ`��@y潯o�3@V�6��!?-� ���@Y%���ٿ4�ǜ`��@y潯o�3@V�6��!?-� ���@Y%���ٿ4�ǜ`��@y潯o�3@V�6��!?-� ���@ަO�ٿ�E����@ �*���3@���ϐ!?����@ަO�ٿ�E����@ �*���3@���ϐ!?����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�WR��ٿ�~Ah���@f�{���3@�Ȼ�!?�[����@�龀,�ٿ�Tԏ
�@��I��3@��㝙�!?����y�@eє�A�ٿғ��8�@%*��3@�#�!��!?'������@�2ނD�ٿ"�jA���@��mO��3@����!?�>����@�2ނD�ٿ"�jA���@��mO��3@����!?�>����@�2ނD�ٿ"�jA���@��mO��3@����!?�>����@�2ނD�ٿ"�jA���@��mO��3@����!?�>����@�2ނD�ٿ"�jA���@��mO��3@����!?�>����@������ٿ��a���@�G؉>�3@%����!?��G��@aJ�+�ٿm�d���@�dT���3@]W
P��!?�(�F��@aJ�+�ٿm�d���@�dT���3@]W
P��!?�(�F��@��􎏤ٿp"��B�@K����3@C��x��!?�yɷ���@��Q�ٿ�pP���@u��>�3@��9�!?�ۆ���@qPT�ٿ�N p?��@� ��3@��f��!?���g=��@qPT�ٿ�N p?��@� ��3@��f��!?���g=��@qPT�ٿ�N p?��@� ��3@��f��!?���g=��@0>�P\�ٿڴ���@�c�	��3@_	���!?�Pd.�@�U���ٿ�`���@�,t��3@F�9>�!?���{�@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@>����ٿ��ܼ���@;)*��3@hQ;�ː!?�̚����@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@-a�*�ٿy��c$��@~���3@�;�n�!?B�C���@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@*O|�B�ٿ�_�����@8A��3@|�	��!?nz�Ō��@M���јٿ9�v�8��@US'��3@X�<��!?LV�bkA�@M���јٿ9�v�8��@US'��3@X�<��!?LV�bkA�@M���јٿ9�v�8��@US'��3@X�<��!?LV�bkA�@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@G>dL�ٿ���#t��@��ݷ@�3@���x�!?����@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@!�ȳ�ٿ�[-P ��@L�qIc�3@8�Ǎ�!?�1(
�@����*�ٿa�ۓ��@h�,��3@u�V�Q�!?1�����@����*�ٿa�ۓ��@h�,��3@u�V�Q�!?1�����@����*�ٿa�ۓ��@h�,��3@u�V�Q�!?1�����@����*�ٿa�ۓ��@h�,��3@u�V�Q�!?1�����@w�����ٿ_}��@�;��3@�a҅ʐ!?'y�`���@w�����ٿ_}��@�;��3@�a҅ʐ!?'y�`���@w�����ٿ_}��@�;��3@�a҅ʐ!?'y�`���@w�����ٿ_}��@�;��3@�a҅ʐ!?'y�`���@w�����ٿ_}��@�;��3@�a҅ʐ!?'y�`���@���ٿ.֠&��@�X�f��3@�j����!?� �R��@���ٿ.֠&��@�X�f��3@�j����!?� �R��@���ٿ.֠&��@�X�f��3@�j����!?� �R��@���ٿ.֠&��@�X�f��3@�j����!?� �R��@���ٿ.֠&��@�X�f��3@�j����!?� �R��@��X�ٿM=t݈��@$��|��3@*�4���!?u�����@?�[�ٿ)���XH�@��y8��3@�	���!?=Z���@�?��՞ٿ�y��b��@�����3@�u<L�!?&�����@YE;9�ٿ4��P<��@��3@��<���!?��]L�u�@YE;9�ٿ4��P<��@��3@��<���!?��]L�u�@YE;9�ٿ4��P<��@��3@��<���!?��]L�u�@YE;9�ٿ4��P<��@��3@��<���!?��]L�u�@)�:�ٿ�}w]��@��3@EaA�ΐ!?�9���r�@)�:�ٿ�}w]��@��3@EaA�ΐ!?�9���r�@)�:�ٿ�}w]��@��3@EaA�ΐ!?�9���r�@�GS2�ٿ!�[Q�f�@L��W,�3@�ֶD��!?�MnX1�@�GS2�ٿ!�[Q�f�@L��W,�3@�ֶD��!?�MnX1�@�GS2�ٿ!�[Q�f�@L��W,�3@�ֶD��!?�MnX1�@�GS2�ٿ!�[Q�f�@L��W,�3@�ֶD��!?�MnX1�@�%��ٿ��1Ϭ��@��Z�3@B�bfِ!?��53�@�%��ٿ��1Ϭ��@��Z�3@B�bfِ!?��53�@�%��ٿ��1Ϭ��@��Z�3@B�bfِ!?��53�@�{�m�ٿx�8�}�@Æ�(��3@���!?��D���@�{�m�ٿx�8�}�@Æ�(��3@���!?��D���@�{�m�ٿx�8�}�@Æ�(��3@���!?��D���@��E�[�ٿH|H����@�ͣ�X�3@J&�Kؐ!?�d���<�@��E�[�ٿH|H����@�ͣ�X�3@J&�Kؐ!?�d���<�@��E�[�ٿH|H����@�ͣ�X�3@J&�Kؐ!?�d���<�@��E�[�ٿH|H����@�ͣ�X�3@J&�Kؐ!?�d���<�@��E�[�ٿH|H����@�ͣ�X�3@J&�Kؐ!?�d���<�@�͖��ٿ{͖��@���5O�3@5a��!?$���e"�@�͖��ٿ{͖��@���5O�3@5a��!?$���e"�@�͖��ٿ{͖��@���5O�3@5a��!?$���e"�@�͖��ٿ{͖��@���5O�3@5a��!?$���e"�@��Y�E�ٿȊБ�D�@���=��3@�a�~<�!?>g�ߔH�@��Y�E�ٿȊБ�D�@���=��3@�a�~<�!?>g�ߔH�@��Y�E�ٿȊБ�D�@���=��3@�a�~<�!?>g�ߔH�@��Y�E�ٿȊБ�D�@���=��3@�a�~<�!?>g�ߔH�@uƺa.�ٿ�pGn�@��B��3@��	2�!?���DI�@uƺa.�ٿ�pGn�@��B��3@��	2�!?���DI�@uƺa.�ٿ�pGn�@��B��3@��	2�!?���DI�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@[�h�ٿdɎ��@�@-��k��3@]�.��!?�3�u3�@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�/�j�ٿ�d:W�@Ûk��3@����!?%I����@�O�`��ٿϑ���2�@ w���3@��V��!?�2�1&�@�O�`��ٿϑ���2�@ w���3@��V��!?�2�1&�@����ٿ���"�@�V ��3@���Ґ!?x������@����ٿ���"�@�V ��3@���Ґ!?x������@����ٿ���"�@�V ��3@���Ґ!?x������@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@���P�ٿ7:!(��@�?����3@��@ϐ!?��a� ��@'��}&�ٿ\�X^ߐ�@���L�3@«�Hِ!? ȝ��|�@���Oٿ�&�����@�C���3@hۦ�!?��cK���@�(7��ٿގ�KA��@���M�3@ t��!?��]~���@�(7��ٿގ�KA��@���M�3@ t��!?��]~���@H�Z�ٿ)*7��w�@�(+��3@ۦ<���!?�?����@H�Z�ٿ)*7��w�@�(+��3@ۦ<���!?�?����@�ؓGҞٿ�����9�@<�[�o�3@"�"��!?�l�\(��@�ؓGҞٿ�����9�@<�[�o�3@"�"��!?�l�\(��@�ؓGҞٿ�����9�@<�[�o�3@"�"��!?�l�\(��@�ؓGҞٿ�����9�@<�[�o�3@"�"��!?�l�\(��@�ؓGҞٿ�����9�@<�[�o�3@"�"��!?�l�\(��@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@C`]���ٿWy��f�@Nl~�3@ԡ��!?I���e�@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@q�P!��ٿ�"�{|��@)��ӏ�3@��А!?�A����@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@���71�ٿ�eY,��@��j�5�3@ape�!?߾?n��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@FQڜB�ٿ�i�ղ��@�R��0�3@������!?W��tu��@X��t��ٿCcl� ��@�Js:��3@/^��Ɛ!?Q��T��@X��t��ٿCcl� ��@�Js:��3@/^��Ɛ!?Q��T��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@uP���ٿ�k+�E�@{^�5 �3@��͐!?aa]�I��@=rܰ�ٿ�?kf��@0�O~��3@�Y5��!?Ú2$4��@=rܰ�ٿ�?kf��@0�O~��3@�Y5��!?Ú2$4��@=rܰ�ٿ�?kf��@0�O~��3@�Y5��!?Ú2$4��@=rܰ�ٿ�?kf��@0�O~��3@�Y5��!?Ú2$4��@��<y��ٿ�pQ0l:�@\/�%��3@-ł�Ԑ!?q.�Ѧ��@���+�ٿ�K�����@甤��3@��e��!?���(��@���+�ٿ�K�����@甤��3@��e��!?���(��@���+�ٿ�K�����@甤��3@��e��!?���(��@���+�ٿ�K�����@甤��3@��e��!?���(��@���+�ٿ�K�����@甤��3@��e��!?���(��@���+�ٿ�K�����@甤��3@��e��!?���(��@��>�ٿ�P�/��@z���3@"�ѧ�!?7�aS��@��>�ٿ�P�/��@z���3@"�ѧ�!?7�aS��@��>�ٿ�P�/��@z���3@"�ѧ�!?7�aS��@��>�ٿ�P�/��@z���3@"�ѧ�!?7�aS��@��>�ٿ�P�/��@z���3@"�ѧ�!?7�aS��@��[�ٿ>�`9�n�@R�o��3@�{=��!?����N#�@��[�ٿ>�`9�n�@R�o��3@�{=��!?����N#�@�O|�S�ٿ9��҂��@]����3@��Ga�!?f�B����@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@�m�)ãٿ�Ⱥt��@��gA�3@�^v�!?�n�9
,�@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@lȧt�ٿ%ݔ&0�@���4�3@���!?��"R��@�6F,!�ٿ�/��4�@]u^�3@p.�G��!?�)z�"��@�6F,!�ٿ�/��4�@]u^�3@p.�G��!?�)z�"��@�6F,!�ٿ�/��4�@]u^�3@p.�G��!?�)z�"��@�6F,!�ٿ�/��4�@]u^�3@p.�G��!?�)z�"��@ή�>�ٿ��BWPE�@<����3@n��"��!?����S��@ή�>�ٿ��BWPE�@<����3@n��"��!?����S��@ή�>�ٿ��BWPE�@<����3@n��"��!?����S��@JzA8͜ٿޑ�����@b�G	J�3@�sdĐ!?�t�:��@���
�ٿ�6���k�@����3@�7�A]�!?e������@���
�ٿ�6���k�@����3@�7�A]�!?e������@�D�t��ٿ���>Ѻ�@2���3@��cb�!?n)P�r��@�D�t��ٿ���>Ѻ�@2���3@��cb�!?n)P�r��@�D�t��ٿ���>Ѻ�@2���3@��cb�!?n)P�r��@�D�t��ٿ���>Ѻ�@2���3@��cb�!?n)P�r��@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@��R�Ǡٿb^�I���@��D��3@9LU۝�!?W�D���@\�����ٿ�r4��@�}K��3@�F+�}�!?l�&*d��@\�����ٿ�r4��@�}K��3@�F+�}�!?l�&*d��@\�����ٿ�r4��@�}K��3@�F+�}�!?l�&*d��@\�����ٿ�r4��@�}K��3@�F+�}�!?l�&*d��@���+�ٿS&�Ӧ��@`�	�3@��5XӐ!?���EȌ�@���+�ٿS&�Ӧ��@`�	�3@��5XӐ!?���EȌ�@���+�ٿS&�Ӧ��@`�	�3@��5XӐ!?���EȌ�@���+�ٿS&�Ӧ��@`�	�3@��5XӐ!?���EȌ�@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@��w��ٿ>��'�7�@O���`�3@ʀP��!?�T#��@ ���ٿSoJ��n�@��q=�3@$\,��!?��_�Ŵ�@ ���ٿSoJ��n�@��q=�3@$\,��!?��_�Ŵ�@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@�.f �ٿ6\'M^�@�\�l�3@�@�'ɐ!?0�d���@fW��ٿPH�)�P�@@�͋=�3@��~�!?b9K1�}�@fW��ٿPH�)�P�@@�͋=�3@��~�!?b9K1�}�@fW��ٿPH�)�P�@@�͋=�3@��~�!?b9K1�}�@fW��ٿPH�)�P�@@�͋=�3@��~�!?b9K1�}�@�9�l�ٿ?H�^�i�@��@
�3@��kݐ!?�t���?�@�9�l�ٿ?H�^�i�@��@
�3@��kݐ!?�t���?�@�9�l�ٿ?H�^�i�@��@
�3@��kݐ!?�t���?�@�9�l�ٿ?H�^�i�@��@
�3@��kݐ!?�t���?�@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@"�y�ٿ���<s��@[�9��3@�cJM��!?�'���@�\4ǡٿش�D�b�@Cd���3@����ǐ!?��G]�@m��P�ٿ�f�H�@����g�3@ׁ}�Ґ!?�1�'��@��z ��ٿ��z�S��@�5����3@��fYߐ!?]�ɹ�H�@��z ��ٿ��z�S��@�5����3@��fYߐ!?]�ɹ�H�@iR���ٿ�1�\�@'�O��3@<=��W�!?�
P?-:�@_2?N��ٿ��CO���@oC��3@z���4�!?��V^�@�[�ۭ�ٿ,n����@G �M��3@ݭ1Rk�!?���BX�@�[�ۭ�ٿ,n����@G �M��3@ݭ1Rk�!?���BX�@�[�ۭ�ٿ,n����@G �M��3@ݭ1Rk�!?���BX�@�3���ٿ�VFsW��@��,�3@C/�3`�!?���=�i�@�3���ٿ�VFsW��@��,�3@C/�3`�!?���=�i�@�3���ٿ�VFsW��@��,�3@C/�3`�!?���=�i�@1�>�ߪٿ�
׃*�@w)�P��3@�1���!?+��?��@y�`ǩٿ%y����@���p��3@i[_+ΐ!?i�q]>�@y�`ǩٿ%y����@���p��3@i[_+ΐ!?i�q]>�@y�`ǩٿ%y����@���p��3@i[_+ΐ!?i�q]>�@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@^d�T�ٿom�����@�l>��3@e�	�Ȑ!?f^6�|��@jDt��ٿ�epE���@�����3@ɵK���!?�\����@jDt��ٿ�epE���@�����3@ɵK���!?�\����@jDt��ٿ�epE���@�����3@ɵK���!?�\����@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@9��!��ٿ��%Z��@�c~D
�3@���^ܐ!?��9kX
�@��9M��ٿY$!�4�@}(n��3@o�J'�!?���b[+�@��9M��ٿY$!�4�@}(n��3@o�J'�!?���b[+�@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@����%�ٿ� t�p�@��`s�3@dHR�!?J't���@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@=Z��ٿ��Ja\��@q�O |�3@�>�SI�!?r�^$�1�@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@7}��:�ٿ���Y1�@9���3@�r`9��!?U�>.2��@-��c��ٿc��(���@����3@��oÊ�!?�����@-��c��ٿc��(���@����3@��oÊ�!?�����@U$���ٿ^��6��@�C�G�3@m��N�!?��T5�@U$���ٿ^��6��@�C�G�3@m��N�!?��T5�@U$���ٿ^��6��@�C�G�3@m��N�!?��T5�@	;c��ٿk_o����@/'�s�3@�j��!?ușw�@3�͗��ٿ�% mm�@}!��3@�	�m�!?x���l�@*��W�ٿ�_��@/���3@C�Y��!?��~�ʑ�@�0���ٿB�I�Q�@���Z�3@7�z�Ր!??#";�k�@��M
��ٿ�	"���@,�:�3@���!?�on����@jU*o��ٿ��b#�@y�����3@����!?p0��/H�@jU*o��ٿ��b#�@y�����3@����!?p0��/H�@jU*o��ٿ��b#�@y�����3@����!?p0��/H�@jU*o��ٿ��b#�@y�����3@����!?p0��/H�@jU*o��ٿ��b#�@y�����3@����!?p0��/H�@����ٿ�i��B�@OZ��3@@EOu֐!?�M��q�@����ٿ�i��B�@OZ��3@@EOu֐!?�M��q�@����ٿ�i��B�@OZ��3@@EOu֐!?�M��q�@����ٿ�i��B�@OZ��3@@EOu֐!?�M��q�@����ٿ�i��B�@OZ��3@@EOu֐!?�M��q�@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@���(e�ٿl�(H��@ws3x�3@��7_�!?
>s.��@�jQ �ٿ0�1���@2�Da�3@�Ed�!?��r����@k�lK��ٿƠb�D�@09x��3@���F��!?z	�[�W�@k�lK��ٿƠb�D�@09x��3@���F��!?z	�[�W�@���~�ٿ�E��7�@��Ӎ{�3@����Ԑ!?�S'��@���~�ٿ�E��7�@��Ӎ{�3@����Ԑ!?�S'��@̎�CX�ٿ�c��� �@�AՂ��3@��"���!?U[��u�@z��yB�ٿ����@գ��Z�3@�:�!?y�vq�@fe�\�ٿ��7���@�0f���3@�V��ې!?���)2��@����)�ٿ<c7���@f5(��3@6}���!?K�Jr��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@�u��G�ٿZ��=�L�@���*��3@�p��͐!?T�x|��@x4���ٿh�8MR(�@Qʞ�y�3@�����!?�a�R}0�@x4���ٿh�8MR(�@Qʞ�y�3@�����!?�a�R}0�@x4���ٿh�8MR(�@Qʞ�y�3@�����!?�a�R}0�@x4���ٿh�8MR(�@Qʞ�y�3@�����!?�a�R}0�@x4���ٿh�8MR(�@Qʞ�y�3@�����!?�a�R}0�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@�3����ٿߙ����@��>X4�3@E�!m�!?.�å�@}��(D�ٿF��
��@��=G�3@q���!?9R8���@}��(D�ٿF��
��@��=G�3@q���!?9R8���@}��(D�ٿF��
��@��=G�3@q���!?9R8���@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�d|�k�ٿ5���'c�@�УԷ�3@˻d��!?/�0�T�@�vY��ٿ�Z��@G�k��3@��&5��!?��`��@�vY��ٿ�Z��@G�k��3@��&5��!?��`��@�vY��ٿ�Z��@G�k��3@��&5��!?��`��@�vY��ٿ�Z��@G�k��3@��&5��!?��`��@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@Z�q�c�ٿ���Y�@B�#W��3@4���Đ!?�.m-;J�@��``�ٿ��Ђ���@�R���3@+��!?z<r��@��``�ٿ��Ђ���@�R���3@+��!?z<r��@S�B��ٿ�	$���@���le�3@��d���!?BI*/�G�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@��ٺ��ٿ�g����@e�O�3@���0��!?�x���9�@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�Oj�@�ٿ> �H��@����3@)�7<�!?v����@�w��ݠٿs>ï��@L����3@��M���!?�Jռ���@�w��ݠٿs>ï��@L����3@��M���!?�Jռ���@�w��ݠٿs>ï��@L����3@��M���!?�Jռ���@�w��ݠٿs>ï��@L����3@��M���!?�Jռ���@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@c��}�ٿ��ˎ�'�@}��5�3@%��^�!?�}��>��@M9e�ٿ���0#I�@Y́�3@U�%�G�!?���-JH�@M9e�ٿ���0#I�@Y́�3@U�%�G�!?���-JH�@9����ٿ�l]i��@H�4�3@|Q�L֐!?i.�.5�@9����ٿ�l]i��@H�4�3@|Q�L֐!?i.�.5�@9����ٿ�l]i��@H�4�3@|Q�L֐!?i.�.5�@9����ٿ�l]i��@H�4�3@|Q�L֐!?i.�.5�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�=6�=�ٿ�6Z�FK�@�ԼT5�3@��[�А!?+��o�q�@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@�.=�ٿ����@v�iU�3@	�V�ݐ!?J1�I���@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@����ٿ]�7]�4�@�B�3@���1�!?Pʶ��@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@�E�깢ٿ�a��6�@a<CU�3@ЅC*�!?�a?�r�@���ٿ�U�/��@����&�3@�})?�!?�e�%A��@���ٿ�U�/��@����&�3@�})?�!?�e�%A��@���ٿ�U�/��@����&�3@�})?�!?�e�%A��@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@i��}��ٿ�r���R�@���K�3@�Z���!?We�����@�}�k�ٿt'�aχ�@d�,8�3@$�OҐ!?����5��@�}�k�ٿt'�aχ�@d�,8�3@$�OҐ!?����5��@�}�k�ٿt'�aχ�@d�,8�3@$�OҐ!?����5��@�}�k�ٿt'�aχ�@d�,8�3@$�OҐ!?����5��@m��ţٿ�����@4�����3@�d�Q �!?�1�]���@m��ţٿ�����@4�����3@�d�Q �!?�1�]���@m��ţٿ�����@4�����3@�d�Q �!?�1�]���@m��ţٿ�����@4�����3@�d�Q �!?�1�]���@m��ţٿ�����@4�����3@�d�Q �!?�1�]���@�ܣ���ٿ"�f9��@�����3@o����!?�ѭ蜽�@�ܣ���ٿ"�f9��@�����3@o����!?�ѭ蜽�@�6'~�ٿ����=�@�h����3@�U� �!?�Q��.}�@�6'~�ٿ����=�@�h����3@�U� �!?�Q��.}�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@}�wϚٿ�?a|\�@� �3@rw���!?S�}d�@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@�z��ٿ/� �Yy�@�o����3@oT���!?�������@T��kW�ٿ]����@I�D�3@J�WԐ!?e3<K��@T��kW�ٿ]����@I�D�3@J�WԐ!?e3<K��@T��kW�ٿ]����@I�D�3@J�WԐ!?e3<K��@B�.�*�ٿ�^B]���@Y-��^�3@HU.˨�!?4,o-���@�gw��ٿ�0�B%��@Tl�]�3@SE�JƐ!?V�E�j�@|����ٿK��U��@�4��3@k��$�!?���x��@���>��ٿZy,���@}����3@��Tx1�!?F�-(�<�@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@�J�)��ٿ�q2)!�@����3@���F�!?S�m���@4b���ٿs�?����@�����3@h�`�!?���DS)�@4b���ٿs�?����@�����3@h�`�!?���DS)�@4b���ٿs�?����@�����3@h�`�!?���DS)�@4b���ٿs�?����@�����3@h�`�!?���DS)�@4b���ٿs�?����@�����3@h�`�!?���DS)�@��ip�ٿ�u��5�@ty[�#�3@���_��!?ld�����@��ip�ٿ�u��5�@ty[�#�3@���_��!?ld�����@�3�S��ٿd^T��@����z�3@	jh�͐!?^P���h�@�3�S��ٿd^T��@����z�3@	jh�͐!?^P���h�@F�g[G�ٿ7���O��@ނ�.�3@���j�!?�4Qt�@F�g[G�ٿ7���O��@ނ�.�3@���j�!?�4Qt�@F�g[G�ٿ7���O��@ނ�.�3@���j�!?�4Qt�@F�g[G�ٿ7���O��@ނ�.�3@���j�!?�4Qt�@7��;k�ٿ/;N����@(
�g�3@b�J.��!?������@7��;k�ٿ/;N����@(
�g�3@b�J.��!?������@7��;k�ٿ/;N����@(
�g�3@b�J.��!?������@7��;k�ٿ/;N����@(
�g�3@b�J.��!?������@7��;k�ٿ/;N����@(
�g�3@b�J.��!?������@b�x�8�ٿ<��p��@��#i��3@A�ؐ!?`���u��@b�x�8�ٿ<��p��@��#i��3@A�ؐ!?`���u��@b�x�8�ٿ<��p��@��#i��3@A�ؐ!?`���u��@b�x�8�ٿ<��p��@��#i��3@A�ؐ!?`���u��@G�M��ٿWٱK��@v(��3@M�|$��!?~ȓ_F��@G�M��ٿWٱK��@v(��3@M�|$��!?~ȓ_F��@CY/���ٿ��x���@0�^ ��3@����!?@١Jv��@CY/���ٿ��x���@0�^ ��3@����!?@١Jv��@�$6�C�ٿ\F����@+_�[e�3@�K��!?�7�Q#O�@���no�ٿ�w���B�@�T��3@o_í�!?��Hއ��@$�Ȱ�ٿ6��LP�@T�p%�3@�t��ΐ!?1ELa��@$�Ȱ�ٿ6��LP�@T�p%�3@�t��ΐ!?1ELa��@���Ҥٿ��SJ��@�,O��3@���禐!?u�g���@����ءٿ�y�6�6�@x� ���3@{+_�!?��s�@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�'��ٿ�G��O~�@���x�3@��!>�!?뢮���@�мA�ٿ�;����@�����3@�0j�)�!?�Qǁ7��@�мA�ٿ�;����@�����3@�0j�)�!?�Qǁ7��@�rX�ٿ�q!aH�@yK30	�3@�����!?J뇢C�@�rX�ٿ�q!aH�@yK30	�3@�����!?J뇢C�@�rX�ٿ�q!aH�@yK30	�3@�����!?J뇢C�@�rX�ٿ�q!aH�@yK30	�3@�����!?J뇢C�@,8�ٿܗY�\�@D��6�3@��n�.�!?i/Y���@,8�ٿܗY�\�@D��6�3@��n�.�!?i/Y���@W�x�ٿ�%B�w��@I��r��3@���!�!?�YG����@W�x�ٿ�%B�w��@I��r��3@���!�!?�YG����@W�x�ٿ�%B�w��@I��r��3@���!�!?�YG����@����ٿ����1�@+�89�3@Q�ت�!?�����@����ٿ����1�@+�89�3@Q�ت�!?�����@����ٿ����1�@+�89�3@Q�ت�!?�����@����ٿ����1�@+�89�3@Q�ت�!?�����@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�5�B�ٿ礼����@�B<e��3@xS�1�!?��8���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@�SA�j�ٿN0���k�@ܨ��3�3@;�[�!?]�l���@m����ٿ�M���@2^���3@� �ꦐ!?��N�[�@m����ٿ�M���@2^���3@� �ꦐ!?��N�[�@m����ٿ�M���@2^���3@� �ꦐ!?��N�[�@Ǯ���ٿnb��Tg�@G�ǑR�3@�*��!?ثǲ:�@Ǯ���ٿnb��Tg�@G�ǑR�3@�*��!?ثǲ:�@��'--�ٿˇ�?��@�P?��3@�F�Z[�!?Q5�
R�@��'--�ٿˇ�?��@�P?��3@�F�Z[�!?Q5�
R�@t����ٿυ�Q�@�9ᣏ�3@���}�!?����T�@4����ٿV�c=���@��h���3@�����!?�;�-�[�@4����ٿV�c=���@��h���3@�����!?�;�-�[�@�^��ٿ�����@�ol��3@�x_��!?�,�I}v�@�^��ٿ�����@�ol��3@�x_��!?�,�I}v�@j�f�I�ٿ�ͣm�?�@r�Jeb�3@�����!?�rF�@d�b��ٿt�\+�"�@�k'�3@5-8Eǐ!?��� �@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@�%0)O�ٿ���AE�@i� �3@� �Ԑ!?t-����@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@J�x7�ٿU�m'���@��j�3@�����!?�е�D��@��G�k�ٿ|ʋu��@��~#R�3@�a�&�!?�e���@��G�k�ٿ|ʋu��@��~#R�3@�a�&�!?�e���@��G�k�ٿ|ʋu��@��~#R�3@�a�&�!?�e���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�#�G��ٿ��I:9h�@�d���3@D���!?�#�P���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@�D�N�ٿٔ���@�R����3@
ԅ�!?��Ɠ���@��ic#�ٿzÕM}x�@�����3@M;,��!?k;MCM�@��ic#�ٿzÕM}x�@�����3@M;,��!?k;MCM�@��ic#�ٿzÕM}x�@�����3@M;,��!?k;MCM�@��ic#�ٿzÕM}x�@�����3@M;,��!?k;MCM�@��ic#�ٿzÕM}x�@�����3@M;,��!?k;MCM�@9��C��ٿ�]#�K��@j}:$�3@X�qÐ!?@L-n�@9��C��ٿ�]#�K��@j}:$�3@X�qÐ!?@L-n�@9��C��ٿ�]#�K��@j}:$�3@X�qÐ!?@L-n�@�@}�ٿ�	��sy�@�d���3@�_qҐ!?��`�&�@�@}�ٿ�	��sy�@�d���3@�_qҐ!?��`�&�@�@}�ٿ�	��sy�@�d���3@�_qҐ!?��`�&�@�@}�ٿ�	��sy�@�d���3@�_qҐ!?��`�&�@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@r�䃞ٿ�l>^�`�@�^A��3@�JO�!?wl�����@#�(�ٿ��qi��@I�4��3@����Ӑ!?��k�S�@#�(�ٿ��qi��@I�4��3@����Ӑ!?��k�S�@��v"�ٿ͝��t��@��n�3@��@��!?;2�ˑ�@��v"�ٿ͝��t��@��n�3@��@��!?;2�ˑ�@�[�N��ٿ�O:��r�@R�t��3@ E�>�!?@R�k��@=���<�ٿF�偁@�@��*��3@�m#��!?m�Jq��@']yMf�ٿ<��W�@ ����3@�vOݐ!?$�M	�@']yMf�ٿ<��W�@ ����3@�vOݐ!?$�M	�@']yMf�ٿ<��W�@ ����3@�vOݐ!?$�M	�@']yMf�ٿ<��W�@ ����3@�vOݐ!?$�M	�@^��Bp�ٿTQ�c�\�@�)P�3@F�:-�!?=H�U:�@^��Bp�ٿTQ�c�\�@�)P�3@F�:-�!?=H�U:�@^��Bp�ٿTQ�c�\�@�)P�3@F�:-�!?=H�U:�@^��Bp�ٿTQ�c�\�@�)P�3@F�:-�!?=H�U:�@aI/��ٿ�p�y���@�r4J�3@R�՜ϐ!?$�[���@aI/��ٿ�p�y���@�r4J�3@R�՜ϐ!?$�[���@�
�Ϣٿ��Q����@�ܝ�v�3@o�PNɐ!?�������@�
�Ϣٿ��Q����@�ܝ�v�3@o�PNɐ!?�������@�
�Ϣٿ��Q����@�ܝ�v�3@o�PNɐ!?�������@�
�Ϣٿ��Q����@�ܝ�v�3@o�PNɐ!?�������@�
�Ϣٿ��Q����@�ܝ�v�3@o�PNɐ!?�������@1sT�t�ٿ�Fkh��@'ͱ���3@^o4RŐ!?�G�ϰ�@1sT�t�ٿ�Fkh��@'ͱ���3@^o4RŐ!?�G�ϰ�@1sT�t�ٿ�Fkh��@'ͱ���3@^o4RŐ!?�G�ϰ�@1sT�t�ٿ�Fkh��@'ͱ���3@^o4RŐ!?�G�ϰ�@1sT�t�ٿ�Fkh��@'ͱ���3@^o4RŐ!?�G�ϰ�@|lE�ٿ�"B��[�@j��#��3@�ڧ@ܐ!?$�����@|lE�ٿ�"B��[�@j��#��3@�ڧ@ܐ!?$�����@I�)�؝ٿB-�'��@W�2��3@�wX���!?�
)'S�@I�)�؝ٿB-�'��@W�2��3@�wX���!?�
)'S�@�2�A~�ٿ#?��X��@����3@��H<��!?$JXж1�@�2�A~�ٿ#?��X��@����3@��H<��!?$JXж1�@�2�A~�ٿ#?��X��@����3@��H<��!?$JXж1�@�2�A~�ٿ#?��X��@����3@��H<��!?$JXж1�@C�=d�ٿr��N���@}�vC�3@�1$ݐ!?���T:O�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@鄠a?�ٿ�O�~V��@�Vz*{�3@�Ej3�!?��=j�@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@��Ε%�ٿ���BT"�@��Qs�3@O֛���!?�����@Nj�'��ٿY�G
9��@�^?1�3@�m�s�!?zx�,��@Nj�'��ٿY�G
9��@�^?1�3@�m�s�!?zx�,��@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@e��f8�ٿ�+Ĕ�O�@�B�f�3@:�x���!?�U%��E�@��]ԣ�ٿ�WnQ�M�@.�Z�3@�ཐ!?4�q����@��]ԣ�ٿ�WnQ�M�@.�Z�3@�ཐ!?4�q����@Xj�Q�ٿ!F�=�@����+�3@e�g��!?(/Z�>�@Xj�Q�ٿ!F�=�@����+�3@e�g��!?(/Z�>�@Xj�Q�ٿ!F�=�@����+�3@e�g��!?(/Z�>�@Xj�Q�ٿ!F�=�@����+�3@e�g��!?(/Z�>�@+��i�ٿST��x�@���h��3@�D3z�!?��?�I�@+��i�ٿST��x�@���h��3@�D3z�!?��?�I�@+��i�ٿST��x�@���h��3@�D3z�!?��?�I�@+��i�ٿST��x�@���h��3@�D3z�!?��?�I�@+��i�ٿST��x�@���h��3@�D3z�!?��?�I�@�;�m�ٿ�:�-p8�@,�!m�3@U��ݐ!?�-��;5�@�;�m�ٿ�:�-p8�@,�!m�3@U��ݐ!?�-��;5�@�;�m�ٿ�:�-p8�@,�!m�3@U��ݐ!?�-��;5�@�;�m�ٿ�:�-p8�@,�!m�3@U��ݐ!?�-��;5�@��K۝ٿgrnMI��@/����3@t�p���!?�l���@��K۝ٿgrnMI��@/����3@t�p���!?�l���@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�,� ��ٿ�A!v�@ߨX�3@	]!+ɐ!?���ɖ\�@�bg�ٿ�$-��@K	���3@��d���!?�`����@��Ir�ٿ�r��o�@��lI�3@�wX��!?cxh7��@��Ir�ٿ�r��o�@��lI�3@�wX��!?cxh7��@�ZH3��ٿ�0��C��@�\��-�3@4��ΐ!?=x�	(��@�ZH3��ٿ�0��C��@�\��-�3@4��ΐ!?=x�	(��@�ZH3��ٿ�0��C��@�\��-�3@4��ΐ!?=x�	(��@�ZH3��ٿ�0��C��@�\��-�3@4��ΐ!?=x�	(��@�ZH3��ٿ�0��C��@�\��-�3@4��ΐ!?=x�	(��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@B�N��ٿ	��v4�@Πx��3@�#���!?u��t8��@5�d��ٿ��q��@�~;��3@��ڢ��!?�C��"��@5�d��ٿ��q��@�~;��3@��ڢ��!?�C��"��@n�N�9�ٿ��qQA��@�OO�(�3@���5��!?���K�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@ݱa��ٿ�mR"�@̰���3@�v$���!?d	z�$�@B�M�ٿ+d�0a�@�b����3@��Ð!?L�����@�����ٿ���d���@I��Z�3@/�S��!?��}� a�@�����ٿ���d���@I��Z�3@/�S��!?��}� a�@	y�2'�ٿ���٧P�@����3@K�Ku|�!?k#�^�w�@	y�2'�ٿ���٧P�@����3@K�Ku|�!?k#�^�w�@��F��ٿ�4��}��@J�k�3@>�
_Ɛ!?�4R��1�@�f���ٿ�YcPF��@j����3@�ی{��!?+R�4�@�f���ٿ�YcPF��@j����3@�ی{��!?+R�4�@
�f,G�ٿ+/�<�=�@Y"R�3@&��|��!?c�Z�K��@
�f,G�ٿ+/�<�=�@Y"R�3@&��|��!?c�Z�K��@
�f,G�ٿ+/�<�=�@Y"R�3@&��|��!?c�Z�K��@
�f,G�ٿ+/�<�=�@Y"R�3@&��|��!?c�Z�K��@�i�8��ٿ��e]���@������3@x⬰�!?=�m=���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@�ʻ��ٿ5��^��@����3@�w���!?�y|���@��U-0�ٿ�q�ٺE�@�W}h�3@�Rx���!?`H���@��U-0�ٿ�q�ٺE�@�W}h�3@�Rx���!?`H���@�mw���ٿL�
��@�X7�3@H1J!?�:�&�@�mw���ٿL�
��@�X7�3@H1J!?�:�&�@d�G�ٿi�G���@�^����3@R���!?�ֽ���@d�G�ٿi�G���@�^����3@R���!?�ֽ���@d�G�ٿi�G���@�^����3@R���!?�ֽ���@d�G�ٿi�G���@�^����3@R���!?�ֽ���@d�G�ٿi�G���@�^����3@R���!?�ֽ���@d�G�ٿi�G���@�^����3@R���!?�ֽ���@p�UF8�ٿ��n����@��h�I�3@:�1��!?�����@p�UF8�ٿ��n����@��h�I�3@:�1��!?�����@p�UF8�ٿ��n����@��h�I�3@:�1��!?�����@�q��ٿӀn|�%�@�k��3@(m��!?7�M]d�@�'��t�ٿ�i��Բ�@�<'��3@�σ�!?=�#HcR�@�'��t�ٿ�i��Բ�@�<'��3@�σ�!?=�#HcR�@�'��t�ٿ�i��Բ�@�<'��3@�σ�!?=�#HcR�@�'��t�ٿ�i��Բ�@�<'��3@�σ�!?=�#HcR�@�'��t�ٿ�i��Բ�@�<'��3@�σ�!?=�#HcR�@:I���ٿ����A�@k�$�3@N��c��!?3����@:I���ٿ����A�@k�$�3@N��c��!?3����@:I���ٿ����A�@k�$�3@N��c��!?3����@:I���ٿ����A�@k�$�3@N��c��!?3����@�e�/y�ٿ������@_x��3@�.S���!?9�]�o~�@�e�/y�ٿ������@_x��3@�.S���!?9�]�o~�@�B�ٿ�C���&�@���}��3@��]�!?	`���a�@�B�ٿ�C���&�@���}��3@��]�!?	`���a�@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@�d�w/�ٿ�1"����@�K>�7�3@A�Z_a�!?Ns0���@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@��ty�ٿ`�ƉB��@ZB��W�3@�4ֈ��!?�~2�z �@w@��ҙٿ��t��@����3@����!?������@w@��ҙٿ��t��@����3@����!?������@w@��ҙٿ��t��@����3@����!?������@w@��ҙٿ��t��@����3@����!?������@w@��ҙٿ��t��@����3@����!?������@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@/�� �ٿXb���@%о[�3@�')��!?�*�S��@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@׹��.�ٿ��Ku�v�@x�\��3@j�����!?wJ���@�Y_�ٿVn�v�@�@
)V�Q�3@�%���!?I�3��@�Y_�ٿVn�v�@�@
)V�Q�3@�%���!?I�3��@�Y_�ٿVn�v�@�@
)V�Q�3@�%���!?I�3��@�1��?�ٿDt0�T��@x8��3@��A�ѐ!?Ԍ����@�1��?�ٿDt0�T��@x8��3@��A�ѐ!?Ԍ����@�1��?�ٿDt0�T��@x8��3@��A�ѐ!?Ԍ����@�����ٿ�a�`�n�@?IO�K�3@4x�~�!?���k��@�����ٿ�a�`�n�@?IO�K�3@4x�~�!?���k��@�����ٿ�a�`�n�@?IO�K�3@4x�~�!?���k��@�����ٿ�a�`�n�@?IO�K�3@4x�~�!?���k��@�����ٿ�a�`�n�@?IO�K�3@4x�~�!?���k��@��'j�ٿ����4�@2Hr��3@�(Pʦ�!?q���[	�@��'j�ٿ����4�@2Hr��3@�(Pʦ�!?q���[	�@��'j�ٿ����4�@2Hr��3@�(Pʦ�!?q���[	�@��'j�ٿ����4�@2Hr��3@�(Pʦ�!?q���[	�@��'j�ٿ����4�@2Hr��3@�(Pʦ�!?q���[	�@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@�j"+�ٿ��AT�B�@u���3@k��Ԑ!?	����@��RGa�ٿ��l�8 �@Dm��m�3@c��z��!?+���:��@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�-����ٿ�UIW�P�@F)���3@jg�]�!?���f�@�տ{�ٿ�-��}�@w�\��3@��O��!?�٤�K��@�)<�ݝٿ�Rr����@�`Z�)�3@��}�!?��Uř?�@�)<�ݝٿ�Rr����@�`Z�)�3@��}�!?��Uř?�@Ne����ٿ̺j�=�@�˃z�3@W�g���!?ŘO�@Ne����ٿ̺j�=�@�˃z�3@W�g���!?ŘO�@Ne����ٿ̺j�=�@�˃z�3@W�g���!?ŘO�@Ne����ٿ̺j�=�@�˃z�3@W�g���!?ŘO�@Ne����ٿ̺j�=�@�˃z�3@W�g���!?ŘO�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@v�Úٿ�0�t��@�z<F�3@��nӐ!?�-�y�@_�B�6�ٿf��h �@b��3@z�Wѐ!?��c<���@�mS��ٿMbd۱��@m���
�3@7�پԐ!?�WY����@�mS��ٿMbd۱��@m���
�3@7�پԐ!?�WY����@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@~Jr<�ٿy,�F,�@�tx��3@����Ԑ!?l�J<5�@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@�Pha�ٿ4"�����@�)����3@]%�Wʐ!?DgY9���@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@|EA1�ٿ�)� ��@����3@wV��!?)k/{,�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@P��@�ٿ�w�V���@�QljO�3@o���!?�d؏�6�@Xy��H�ٿ�jhO��@5G��3@�����!?B�pG��@��o���ٿ�3���@ω5�3@G��7��!?\�P��@��o���ٿ�3���@ω5�3@G��7��!?\�P��@��o���ٿ�3���@ω5�3@G��7��!?\�P��@��o���ٿ�3���@ω5�3@G��7��!?\�P��@��o���ٿ�3���@ω5�3@G��7��!?\�P��@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@���>�ٿ�S'�@Q��t#�3@<-Jx��!?!�����@��hD�ٿɛ�EE�@!�Y��3@�Q�Ő!?q�U����@��hD�ٿɛ�EE�@!�Y��3@�Q�Ő!?q�U����@��hD�ٿɛ�EE�@!�Y��3@�Q�Ő!?q�U����@?8�ߙٿ]D˿�@�f��n�3@���Ɛ!?E���w��@?8�ߙٿ]D˿�@�f��n�3@���Ɛ!?E���w��@x�G̝ٿfN?��@�I>���3@�����!?U�(�P�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@��t[��ٿ�"����@�c���3@���ǐ!?�1�0�@�AP+��ٿF���c�@Aq�C�3@bB]=Ȑ!?���ܼ�@"?�͗�ٿ��=i��@��+�i�3@-ݾ�!?�+\A��@"?�͗�ٿ��=i��@��+�i�3@-ݾ�!?�+\A��@"?�͗�ٿ��=i��@��+�i�3@-ݾ�!?�+\A��@�Q"��ٿ[��>��@F��1>�3@����*�!?�n�T��@�Q"��ٿ[��>��@F��1>�3@����*�!?�n�T��@�Q"��ٿ[��>��@F��1>�3@����*�!?�n�T��@�H�Y�ٿ����@Z%��3@H�;=�!?�+��K�@�H�Y�ٿ����@Z%��3@H�;=�!?�+��K�@�H�Y�ٿ����@Z%��3@H�;=�!?�+��K�@2���ٿ�x6�>��@.o}��3@��z�!?���4m!�@��ب�ٿJ�$H�>�@�J��t�3@ ���!?��if��@��ب�ٿJ�$H�>�@�J��t�3@ ���!?��if��@�udٿ���B��@w����3@K�&,�!?3�d�^�@�udٿ���B��@w����3@K�&,�!?3�d�^�@ٹ��ٿ9���[�@���j�3@K`n��!?R��ą�@ٹ��ٿ9���[�@���j�3@K`n��!?R��ą�@ٹ��ٿ9���[�@���j�3@K`n��!?R��ą�@��ۡٿ��蜾��@�bfD�3@B���!?7
�9��@��ۡٿ��蜾��@�bfD�3@B���!?7
�9��@��ۡٿ��蜾��@�bfD�3@B���!?7
�9��@)�S�[�ٿj����@s�I�y�3@3_�i`�!?��zd��@)�S�[�ٿj����@s�I�y�3@3_�i`�!?��zd��@)�S�[�ٿj����@s�I�y�3@3_�i`�!?��zd��@)�S�[�ٿj����@s�I�y�3@3_�i`�!?��zd��@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@�I>2�ٿ �#�X��@���3@��4�q�!?n��Z�@9q,y�ٿ9Gl�_#�@�J0�y�3@Lwlʗ�!?+5õS��@9q,y�ٿ9Gl�_#�@�J0�y�3@Lwlʗ�!?+5õS��@�S,#Śٿ5�m�@s���3@?�'͐!?�
��@�S,#Śٿ5�m�@s���3@?�'͐!?�
��@��Q�ٿ)<2T��@������3@��o��!?�6$�J�@��Q�ٿ)<2T��@������3@��o��!?�6$�J�@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@��싘ٿ�u�#i�@(z�8�3@N����!?�Uc�*��@>�t��ٿ��%���@.Tz��3@��А!?~�����@>�t��ٿ��%���@.Tz��3@��А!?~�����@���j��ٿaMO�	 �@�D��3@�B��ܐ!?K[R�"�@���j��ٿaMO�	 �@�D��3@�B��ܐ!?K[R�"�@���j��ٿaMO�	 �@�D��3@�B��ܐ!?K[R�"�@�R�P�ٿ��Z7��@��>��3@�"RP��!?�Ke ���@�R�P�ٿ��Z7��@��>��3@�"RP��!?�Ke ���@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@]nȚ\�ٿ�i8�G��@X���3@�ϴ���!?X1�3YV�@_qM�_�ٿẺ2w`�@�̣C��3@�����!?!oL���@��hS�ٿ-�0�_��@f���3@qs�ؐ!?Hx>��@��hS�ٿ-�0�_��@f���3@qs�ؐ!?Hx>��@��hS�ٿ-�0�_��@f���3@qs�ؐ!?Hx>��@��hS�ٿ-�0�_��@f���3@qs�ؐ!?Hx>��@n�7b�ٿ_�=��j�@T�BO��3@�a:ې!?]fG޿�@�tuդٿ��)$a]�@6��g�3@o�N#�!?C2�o7��@���åٿtXJ/+�@�1�3@J9?�!?�����*�@���åٿtXJ/+�@�1�3@J9?�!?�����*�@���åٿtXJ/+�@�1�3@J9?�!?�����*�@���åٿtXJ/+�@�1�3@J9?�!?�����*�@���åٿtXJ/+�@�1�3@J9?�!?�����*�@���åٿtXJ/+�@�1�3@J9?�!?�����*�@3����ٿ� ����@pV-MU�3@��^��!?��ֹ�@3����ٿ� ����@pV-MU�3@��^��!?��ֹ�@3����ٿ� ����@pV-MU�3@��^��!?��ֹ�@3����ٿ� ����@pV-MU�3@��^��!?��ֹ�@3����ٿ� ����@pV-MU�3@��^��!?��ֹ�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@w�m�ٿ�ؼG��@�:��;�3@��;��!?��d�@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@3���ٿ�5�����@s+N���3@$b@c|�!?�q���@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@��xݟٿ�@�g,Y�@����3@A�MŐ!?[�)�R��@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@8*ЍҚٿ���}�L�@����3@9�,Iɐ!?ݷi/|S�@�9��ٿ�G���9�@?!����3@^�)�А!?XW��@��@�9��ٿ�G���9�@?!����3@^�)�А!?XW��@��@�9��ٿ�G���9�@?!����3@^�)�А!?XW��@��@�9��ٿ�G���9�@?!����3@^�)�А!?XW��@��@�@�.Κٿ"�g��@�*�A$�3@ �ш�!?�ȶ���@�@�.Κٿ"�g��@�*�A$�3@ �ш�!?�ȶ���@���U�ٿn$�xm"�@������3@n�"M֐!?O֒��`�@���U�ٿn$�xm"�@������3@n�"M֐!?O֒��`�@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@���C�ٿ�ZuM�@�?^�J�3@������!?M~��@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@�¥z,�ٿj6��ŕ�@5�����3@����!?Gĥ-P�@M��J[�ٿ��%o��@�v��3@z�o8��!?�f����@U!Ke��ٿQY���@y@ 2^�3@u!��!?f�,,�R�@U!Ke��ٿQY���@y@ 2^�3@u!��!?f�,,�R�@U!Ke��ٿQY���@y@ 2^�3@u!��!?f�,,�R�@U!Ke��ٿQY���@y@ 2^�3@u!��!?f�,,�R�@�/���ٿ��(����@ѫ����3@�)�!?и�>���@�/���ٿ��(����@ѫ����3@�)�!?и�>���@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@�ɇ�ٿg�����@������3@۽M��!?��ws��@��� <�ٿ{@@O���@�A����3@��>���!?�b0Uá�@��� <�ٿ{@@O���@�A����3@��>���!?�b0Uá�@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�ן���ٿ�i Ɍ��@�xI��3@(�ِ!?V���@�[�a�ٿHg6��@�g2,��3@�a�x�!?�"o28�@���h)�ٿ��'��@�K�\��3@�F��!?t�7{/_�@���h)�ٿ��'��@�K�\��3@�F��!?t�7{/_�@���h)�ٿ��'��@�K�\��3@�F��!?t�7{/_�@���h)�ٿ��'��@�K�\��3@�F��!?t�7{/_�@���h)�ٿ��'��@�K�\��3@�F��!?t�7{/_�@�!~�כٿ�y�s�<�@�T.�d�3@��q���!?4�]=J�@�;}!�ٿ3@�L �@��ek�3@ކ_֐!?d����9�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@Lxj�ڝٿ�kg����@��>:��3@��l��!?l�k�@q���g�ٿ����:��@=O�J�3@�BO��!?�sPƮB�@q���g�ٿ����:��@=O�J�3@�BO��!?�sPƮB�@q���g�ٿ����:��@=O�J�3@�BO��!?�sPƮB�@})��̡ٿ>ϸ����@ь�!��3@�*�%j�!?F�e���@})��̡ٿ>ϸ����@ь�!��3@�*�%j�!?F�e���@})��̡ٿ>ϸ����@ь�!��3@�*�%j�!?F�e���@})��̡ٿ>ϸ����@ь�!��3@�*�%j�!?F�e���@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���՞�ٿ̗n�x[�@����3@'��!?'&���(�@���`�ٿ�%��]�@M��0�3@;��;Ȑ!?���]��@���`�ٿ�%��]�@M��0�3@;��;Ȑ!?���]��@���`�ٿ�%��]�@M��0�3@;��;Ȑ!?���]��@���`�ٿ�%��]�@M��0�3@;��;Ȑ!?���]��@���`�ٿ�%��]�@M��0�3@;��;Ȑ!?���]��@�ɶ�՚ٿQ� ���@�?�5r�3@�3��4�!?8����@�ɶ�՚ٿQ� ���@�?�5r�3@�3��4�!?8����@�ɶ�՚ٿQ� ���@�?�5r�3@�3��4�!?8����@�ɶ�՚ٿQ� ���@�?�5r�3@�3��4�!?8����@�ɶ�՚ٿQ� ���@�?�5r�3@�3��4�!?8����@aI��ٿ��NB�@����u�3@6#�� �!?�Xq��@aI��ٿ��NB�@����u�3@6#�� �!?�Xq��@aI��ٿ��NB�@����u�3@6#�� �!?�Xq��@aI��ٿ��NB�@����u�3@6#�� �!?�Xq��@�\_��ٿ�(>n  �@�t~g?�3@��Fc�!?��/m��@�\_��ٿ�(>n  �@�t~g?�3@��Fc�!?��/m��@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@�Y*+�ٿ���~G��@R;H��3@<�J�6�!?)ޢ�c/�@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@.��ٿƧY�Ē�@y=J��3@�!U��!?TI���@X����ٿ���ɝ��@/�o^��3@���ѱ�!?i1aG;��@X����ٿ���ɝ��@/�o^��3@���ѱ�!?i1aG;��@X����ٿ���ɝ��@/�o^��3@���ѱ�!?i1aG;��@X����ٿ���ɝ��@/�o^��3@���ѱ�!?i1aG;��@X����ٿ���ɝ��@/�o^��3@���ѱ�!?i1aG;��@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@ٜ����ٿ�Fƚ��@m[!��3@3ꉀ��!?r+�����@��U�Ϧٿ"�o�~�@������3@HY�U��!?���D�d�@[w��ٿ�2�g��@H�x��3@o�1;P�!?o,��� �@�[�Ԥٿ���'��@;o<� 4@v߀���!?���{��@ �� �ٿ��ԫz�@��+E4@��0�!?�v��k�@'��	�ٿN(�;��@�m|�3@v0��!?���Ku�@'��	�ٿN(�;��@�m|�3@v0��!?���Ku�@'��	�ٿN(�;��@�m|�3@v0��!?���Ku�@'��	�ٿN(�;��@�m|�3@v0��!?���Ku�@'��	�ٿN(�;��@�m|�3@v0��!?���Ku�@Z�"(�ٿ�8�r���@�*���3@鯆ۘ�!?q��C$g�@Z�"(�ٿ�8�r���@�*���3@鯆ۘ�!?q��C$g�@Z�"(�ٿ�8�r���@�*���3@鯆ۘ�!?q��C$g�@Z�"(�ٿ�8�r���@�*���3@鯆ۘ�!?q��C$g�@Z�"(�ٿ�8�r���@�*���3@鯆ۘ�!?q��C$g�@-	-��ٿ�c��%X�@O�٪�3@am���!?����D�@-	-��ٿ�c��%X�@O�٪�3@am���!?����D�@-	-��ٿ�c��%X�@O�٪�3@am���!?����D�@-	-��ٿ�c��%X�@O�٪�3@am���!?����D�@-	-��ٿ�c��%X�@O�٪�3@am���!?����D�@����ٿ[�����@�7��3@7�Gs�!?��9;�@	Y��ٿ %��@�p����3@��e� �!?1r��a��@&�q��ٿp�JФ��@�^�ǉ�3@1'8r�!?�¯�Bg�@&�q��ٿp�JФ��@�^�ǉ�3@1'8r�!?�¯�Bg�@������ٿ��`=�z�@-�l��3@������!?�'�@������ٿ��`=�z�@-�l��3@������!?�'�@������ٿ��`=�z�@-�l��3@������!?�'�@�N0%��ٿ�J����@Z�%��3@i��Ҟ�!?�z�>}�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@��>�ٿ0t_G�@IM���3@�wPlڐ!?�UwޖJ�@/���ٿ�Ǣ)��@���3@�u��!?)+ R��@/���ٿ�Ǣ)��@���3@�u��!?)+ R��@/���ٿ�Ǣ)��@���3@�u��!?)+ R��@/���ٿ�Ǣ)��@���3@�u��!?)+ R��@���ٿS��Y��@�X���3@�c�"�!?k�(���@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@HT�Ӡٿ1:+	
�@ȜN�X�3@
����!?AV����@��刴�ٿ3�8b��@5lx�p�3@`Ik?�!?��6�k��@��刴�ٿ3�8b��@5lx�p�3@`Ik?�!?��6�k��@��刴�ٿ3�8b��@5lx�p�3@`Ik?�!?��6�k��@��0��ٿ^E)���@��(�3@q�v��!?�G�eiy�@��NE�ٿ��=^��@�\���3@�S���!?l�ӾDO�@��NE�ٿ��=^��@�\���3@�S���!?l�ӾDO�@,�V�ٿ�^ڈ���@��ϗ��3@����!?�]W@��@,�V�ٿ�^ڈ���@��ϗ��3@����!?�]W@��@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�*��ٿ�0L
bB�@�T����3@HL�h
�!?�����@�ݑ���ٿ�tvvn�@B�K���3@(��<�!?�����@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@�,�G�ٿoK&Ƥ��@�&&�3@Bz71�!?~��G��@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���K�ٿ�gN_r�@���kY�3@��4�!?���~�@���.ٿ|���%�@��r�0�3@Oo=V�!?���k�y�@���.ٿ|���%�@��r�0�3@Oo=V�!?���k�y�@]�˛ٿ�#�s�@YZ��S�3@)��eʐ!?���i���@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�ԕ㧛ٿ;�zy<�@>#9��3@�2�h��!?�ĉV�`�@�Ƹ�ٿ��]�@k)��S�3@w/O��!?3�z��@�Ƹ�ٿ��]�@k)��S�3@w/O��!?3�z��@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@��m��ٿ��?�L�@�q����3@5n��!?v̑T���@g�=I�ٿ���$p[�@�B���3@*|+�Ð!?2k���@g�=I�ٿ���$p[�@�B���3@*|+�Ð!?2k���@g�=I�ٿ���$p[�@�B���3@*|+�Ð!?2k���@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@Sa�A�ٿ	F����@fBVe�3@��Bʐ!?ޜw4��@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�E�K��ٿHW.��@>��3@��;��!?}�q@)m�@�JN�ٿ9'b�|�@q
�N�3@�:���!?Q�?��@�JN�ٿ9'b�|�@q
�N�3@�:���!?Q�?��@��x�ٿ��F�]��@A����3@2�ٗ�!?fnC���@��x�ٿ��F�]��@A����3@2�ٗ�!?fnC���@��x�ٿ��F�]��@A����3@2�ٗ�!?fnC���@�;�s�ٿ��kZ/}�@��0��3@��{���!?0�4R*��@�S&�ٿ��3|sg�@�#w��3@��*��!?n�E�zZ�@�S&�ٿ��3|sg�@�#w��3@��*��!?n�E�zZ�@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@]'j�ٿpj1��P�@xWp�v�3@}���!?N��g��@-�Z��ٿkn����@~���S�3@L�r��!?B8*r�}�@�1�$��ٿ�p���@c����3@�����!?נR����@�1�$��ٿ�p���@c����3@�����!?נR����@�1�$��ٿ�p���@c����3@�����!?נR����@g��O�ٿEֱ�&r�@Eq�3@��!?L�T�@g��O�ٿEֱ�&r�@Eq�3@��!?L�T�@g��O�ٿEֱ�&r�@Eq�3@��!?L�T�@g��O�ٿEֱ�&r�@Eq�3@��!?L�T�@����<�ٿ/����q�@��!O�3@�PB��!?a(ۦ���@����<�ٿ/����q�@��!O�3@�PB��!?a(ۦ���@����<�ٿ/����q�@��!O�3@�PB��!?a(ۦ���@�H��q�ٿ�j��>��@
��G�3@!�#���!?���M��@�H��q�ٿ�j��>��@
��G�3@!�#���!?���M��@�V1a�ٿb����@��܅E�3@ѹ����!?q�$�@�V1a�ٿb����@��܅E�3@ѹ����!?q�$�@�V1a�ٿb����@��܅E�3@ѹ����!?q�$�@zRN^�ٿ�뷤&��@�V?�#�3@w/K���!?|��8%R�@zRN^�ٿ�뷤&��@�V?�#�3@w/K���!?|��8%R�@zRN^�ٿ�뷤&��@�V?�#�3@w/K���!?|��8%R�@zRN^�ٿ�뷤&��@�V?�#�3@w/K���!?|��8%R�@zRN^�ٿ�뷤&��@�V?�#�3@w/K���!?|��8%R�@u�w�ٿ�]M���@�y�n�3@���9��!?�9�9,P�@u�w�ٿ�]M���@�y�n�3@���9��!?�9�9,P�@u�w�ٿ�]M���@�y�n�3@���9��!?�9�9,P�@�oU��ٿ^�'L��@NY� ��3@��@@Ґ!?<|��h��@��Y�ٿĝ��@�[��c�3@���B��!?�����@��Y�ٿĝ��@�[��c�3@���B��!?�����@�߈a;�ٿ~,��%�@}�{��3@ߒSyÐ!?/gB���@�߈a;�ٿ~,��%�@}�{��3@ߒSyÐ!?/gB���@0GH���ٿ�2fޙ��@��.I-�3@V3�i��!?&X]qa�@LKV`a�ٿ�L���@��eW�3@����
�!?�M�$���@LKV`a�ٿ�L���@��eW�3@����
�!?�M�$���@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@4�ʚ�ٿ�o
Q��@���1��3@�I��!?��v#��@��Ҟ�ٿ�ܲl�\�@S�+g�3@P��J�!?��)�L,�@��Ҟ�ٿ�ܲl�\�@S�+g�3@P��J�!?��)�L,�@�S/�ٿd������@?��N�3@�>�!?��w����@�S/�ٿd������@?��N�3@�>�!?��w����@�S/�ٿd������@?��N�3@�>�!?��w����@�S/�ٿd������@?��N�3@�>�!?��w����@�S/�ٿd������@?��N�3@�>�!?��w����@�\�k�ٿ��}����@\c�^�3@K�J��!?��G^��@�\�k�ٿ��}����@\c�^�3@K�J��!?��G^��@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@��~.�ٿbޛ���@>�!<��3@�(��!?0C�aް�@=��ٿ��^�@��9�3@��T��!?d�L9��@=��ٿ��^�@��9�3@��T��!?d�L9��@Ef��A�ٿ����y)�@�|J��3@(vA��!?���@A��@���И�ٿ�6I���@B�I 4@������!?�����@���И�ٿ�6I���@B�I 4@������!?�����@���И�ٿ�6I���@B�I 4@������!?�����@���И�ٿ�6I���@B�I 4@������!?�����@���И�ٿ�6I���@B�I 4@������!?�����@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@h��:O�ٿ���h�#�@ ���3@6�)Ӑ!?�.�|��@ǐ�L��ٿ䦧�R��@����3@'E����!?���){�@ǐ�L��ٿ䦧�R��@����3@'E����!?���){�@ǐ�L��ٿ䦧�R��@����3@'E����!?���){�@ǐ�L��ٿ䦧�R��@����3@'E����!?���){�@i�����ٿ��K�@�,q�3@�V.T/�!?��x����@i�����ٿ��K�@�,q�3@�V.T/�!?��x����@i�����ٿ��K�@�,q�3@�V.T/�!?��x����@�ut�ٿ����I7�@)<�0��3@ �"��!?�S>���@��$�j�ٿG�,���@ߌsN�3@��e=�!? �d���@��$�j�ٿG�,���@ߌsN�3@��e=�!? �d���@	ݝ�|�ٿI��z���@޽m���3@׫&�!?���v�@I�f^B�ٿ&#e�:�@75WT�3@]��"%�!?.�v�@I�f^B�ٿ&#e�:�@75WT�3@]��"%�!?.�v�@���ŗٿ��Ȑ�O�@S��]��3@4�v��!?d�{����@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@�4���ٿ�{�����@�b�%X�3@&�G4�!?�n��@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@��D�ٿ�4�xX��@�c�=��3@Tд�!?(]��(�@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@�5�Y�ٿ�����@����3@/wz��!?w%G��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���bѡٿ�:0%V�@�'^���3@5�����!?�E��@���ٿ��Y��@�����3@2>���!?�d_�"&�@���ٿ��Y��@�����3@2>���!?�d_�"&�@���ٿ��Y��@�����3@2>���!?�d_�"&�@���ٿ��Y��@�����3@2>���!?�d_�"&�@���ٿ��Y��@�����3@2>���!?�d_�"&�@�宽�ٿ%_V�#R�@�o�l_�3@���^)�!?��ZP ��@u9
�ܗٿ2��<�F�@�����3@>Il@�!?��'�!~�@zzP�ٿm`� ��@b(nG��3@�/�W��!?F�
%ʧ�@!A�x`�ٿgd��IA�@������3@^L�O�!?j�����@��A��ٿ�#6M�@�����3@��6��!?�
��(�@�zJ�0�ٿ�tr���@*5����3@��>��!?Rɕo?��@�zJ�0�ٿ�tr���@*5����3@��>��!?Rɕo?��@�o	k�ٿc������@��d���3@����!?�ZP�U��@�o	k�ٿc������@��d���3@����!?�ZP�U��@�5.��ٿ�t	t�2�@�z1�3@�;"��!?F�[I��@�5.��ٿ�t	t�2�@�z1�3@�;"��!?F�[I��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@*8F'M�ٿ5�B�z��@8'`@��3@�g0ܯ�!?��*C��@�*wu�ٿg@�В �@r�/L��3@ـb��!?]	#�$��@�*wu�ٿg@�В �@r�/L��3@ـb��!?]	#�$��@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@u����ٿڅl��`�@�c#�3@�y�7ΐ!?s2����@��@π�ٿ�f�����@~K*��3@j2���!?�p���@��l�ٿ3�_�2L�@*����3@b�|��!?:�v�K��@��l�ٿ3�_�2L�@*����3@b�|��!?:�v�K��@��l�ٿ3�_�2L�@*����3@b�|��!?:�v�K��@&�	��ٿ��?�L�@�qY���3@D�ԐF�!?�(YB46�@&�	��ٿ��?�L�@�qY���3@D�ԐF�!?�(YB46�@�;�pr�ٿn�Ѽ��@��T���3@j���X�!?��@���@�;�pr�ٿn�Ѽ��@��T���3@j���X�!?��@���@�;�pr�ٿn�Ѽ��@��T���3@j���X�!?��@���@�;�pr�ٿn�Ѽ��@��T���3@j���X�!?��@���@�;�pr�ٿn�Ѽ��@��T���3@j���X�!?��@���@B��$�ٿZ�|L���@pUվ�3@9+=�א!?�|%�}��@B��$�ٿZ�|L���@pUվ�3@9+=�א!?�|%�}��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@�Йm��ٿ�Z����@��	J��3@�����!?)o
>)��@���:�ٿ�ٰ�*x�@�nz�3@s���!?��m�?��@���:�ٿ�ٰ�*x�@�nz�3@s���!?��m�?��@���:�ٿ�ٰ�*x�@�nz�3@s���!?��m�?��@���:�ٿ�ٰ�*x�@�nz�3@s���!?��m�?��@��"o̞ٿN�J���@���8��3@[�Xwː!?�ݯ�c�@A'���ٿ�]F!]��@AB�H�3@Q�7@��!?;6o��@�n��ٿ�C�CS�@��7��3@����!?,�뙺.�@�n��ٿ�C�CS�@��7��3@����!?,�뙺.�@�n��ٿ�C�CS�@��7��3@����!?,�뙺.�@�n��ٿ�C�CS�@��7��3@����!?,�뙺.�@�n��ٿ�C�CS�@��7��3@����!?,�뙺.�@Z�?b��ٿR��_�@�T�T�3@$0�ڐ!?��y,��@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�}���ٿmD��@9X��3@o5唡�!?_��\�@�|��ݟٿ`�E����@�����3@��#�!?��{�T��@�|��ݟٿ`�E����@�����3@��#�!?��{�T��@�|��ݟٿ`�E����@�����3@��#�!?��{�T��@�|��ݟٿ`�E����@�����3@��#�!?��{�T��@�|��ݟٿ`�E����@�����3@��#�!?��{�T��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@y��yڞٿ�m�����@I�&Q�3@CЙC
�!?jG�{f��@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@��6���ٿ�D�"��@���^�3@�Wِ!?^K+T�@X���V�ٿFe'h=�@.��G�3@?��Z�!?*�����@{�8:N�ٿ4�Ն�@������3@X-=�!?���G�@{�8:N�ٿ4�Ն�@������3@X-=�!?���G�@{�8:N�ٿ4�Ն�@������3@X-=�!?���G�@cQ)��ٿ�
� �@�2^gW�3@������!?�� N���@cQ)��ٿ�
� �@�2^gW�3@������!?�� N���@cQ)��ٿ�
� �@�2^gW�3@������!?�� N���@cQ)��ٿ�
� �@�2^gW�3@������!?�� N���@��L��ٿ_{��7��@��[� �3@�"RՐ!?
ѡ��=�@���7Ȝٿ���跺�@�����3@w����!?�+�j��@���7Ȝٿ���跺�@�����3@w����!?�+�j��@���7Ȝٿ���跺�@�����3@w����!?�+�j��@�r�xl�ٿDn=�o�@�:��3@2um�ې!?�&@�=�@�r�xl�ٿDn=�o�@�:��3@2um�ې!?�&@�=�@�b[���ٿ������@"�9�W�3@wW6�!??�!y��@�b[���ٿ������@"�9�W�3@wW6�!??�!y��@�b[���ٿ������@"�9�W�3@wW6�!??�!y��@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@9��i�ٿ�.~"01�@�0�"��3@K����!?)�p����@�_�10�ٿ���yX�@�����3@�R�!?ҿEG���@�_�10�ٿ���yX�@�����3@�R�!?ҿEG���@�_�10�ٿ���yX�@�����3@�R�!?ҿEG���@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@`Z�P�ٿ2��9�@r6�#��3@��Ix��!?�$��S��@�L��P�ٿ{N�7\��@�+-I��3@�۲<��!?#��_-��@�L��P�ٿ{N�7\��@�+-I��3@�۲<��!?#��_-��@�8;b��ٿ� ~ƽ�@c6K�-�3@d�١�!?sa+���@��j��ٿyQI-9�@��n�@�3@F�v�Đ!?B�y����@��j��ٿyQI-9�@��n�@�3@F�v�Đ!?B�y����@��j��ٿyQI-9�@��n�@�3@F�v�Đ!?B�y����@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@�-n��ٿaUj��@��&��3@\�u��!?E��ƅ��@iЏ�ٿ�X�c-��@�k�3@��|�ϐ!?}U��N�@iЏ�ٿ�X�c-��@�k�3@��|�ϐ!?}U��N�@�/=�a�ٿs_k~��@i?7�3@�]�hΐ!?�P���,�@�'#T�ٿ�^ U���@��.��3@ͩ%�Ő!?�t K"]�@�'#T�ٿ�^ U���@��.��3@ͩ%�Ő!?�t K"]�@�'#T�ٿ�^ U���@��.��3@ͩ%�Ő!?�t K"]�@�'#T�ٿ�^ U���@��.��3@ͩ%�Ő!?�t K"]�@�ct�ٿ�iaņ�@�Ӣ���3@��eu��!?�y5RE�@�ct�ٿ�iaņ�@�Ӣ���3@��eu��!?�y5RE�@�ct�ٿ�iaņ�@�Ӣ���3@��eu��!?�y5RE�@�ct�ٿ�iaņ�@�Ӣ���3@��eu��!?�y5RE�@{c�ӣٿ(���{�@�@��3@��L��!?�gݹ`�@{c�ӣٿ(���{�@�@��3@��L��!?�gݹ`�@{c�ӣٿ(���{�@�@��3@��L��!?�gݹ`�@{c�ӣٿ(���{�@�@��3@��L��!?�gݹ`�@{c�ӣٿ(���{�@�@��3@��L��!?�gݹ`�@F�U�ٿ�^v2��@�#eה�3@��(Ґ!?��h�gk�@F�U�ٿ�^v2��@�#eה�3@��(Ґ!?��h�gk�@F�U�ٿ�^v2��@�#eה�3@��(Ґ!?��h�gk�@F�U�ٿ�^v2��@�#eה�3@��(Ґ!?��h�gk�@�.ޔ�ٿa2���@�*m��3@�[HՐ!?���N�@�.ޔ�ٿa2���@�*m��3@�[HՐ!?���N�@�.ޔ�ٿa2���@�*m��3@�[HՐ!?���N�@�.ޔ�ٿa2���@�*m��3@�[HՐ!?���N�@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@YwL�	�ٿϛ�7�0�@��3@�Z����!?f5�8E��@�?[N�ٿ>I��?��@�����3@�mǯi�!?�� �%�@�?[N�ٿ>I��?��@�����3@�mǯi�!?�� �%�@�?[N�ٿ>I��?��@�����3@�mǯi�!?�� �%�@Mh��t�ٿD�7I��@�f*D��3@@�y:��!?��1Y�@,���U�ٿH���ǿ�@N[l�z�3@�ġ;�!?6��� �@,���U�ٿH���ǿ�@N[l�z�3@�ġ;�!?6��� �@q�8�ٿIs5vQ�@�u����3@~qh��!?M��ΤJ�@q�8�ٿIs5vQ�@�u����3@~qh��!?M��ΤJ�@�νu>�ٿ̀�w�9�@�F�z��3@vm����!?��fʳ�@/�0�ٿt�-/O�@�����3@���!?�f�}]�@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@}���ٿ��IvD�@��Dz��3@9Mȫ�!?\Ε���@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@2��Ƥٿ�J����@��U���3@jn-��!?�"z�u�@@4F�ΞٿcJ�?#�@�� �3@G~�!?��Ĉ�`�@@4F�ΞٿcJ�?#�@�� �3@G~�!?��Ĉ�`�@w��ҚٿΥ$�l�@oԀx�3@k�o���!?_�z}��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@�N˭�ٿ���
�F�@����3@�Lw��!?�!q�k��@��]��ٿf3y==I�@���{J�3@[K��ѐ!?*��CH�@��]��ٿf3y==I�@���{J�3@[K��ѐ!?*��CH�@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��{8٢ٿ A��*��@l %4��3@zB�K͐!?U������@��V>�ٿ�+�����@D��'��3@Ԇ�� �!?#I�/+��@/�(o#�ٿA�0��\�@�78v��3@{u���!?s�3Of�@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@��
�ɣٿ	?k��@.~�(��3@� d��!?���>j��@�,���ٿQwzF�@3�q�m�3@l�k �!?�)��/��@��-5�ٿ�o��3�@w�j/�3@=>�Ɛ!?y�5���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@r�����ٿ�3��/�@��WK�3@��I`!?�Fɸ���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�	�ޙٿY�7��@� h���3@C3�f�!??O˯���@�P{�V�ٿ�,)H�X�@l ���3@Ҳ����!?�L�ۋ��@����ٿ�H�tO0�@��aZ�3@��cd��!?��WV�Q�@����ٿ�H�tO0�@��aZ�3@��cd��!?��WV�Q�@����ٿ�H�tO0�@��aZ�3@��cd��!?��WV�Q�@����ٿ�H�tO0�@��aZ�3@��cd��!?��WV�Q�@����ٿ�H�tO0�@��aZ�3@��cd��!?��WV�Q�@�q2�Пٿ��Y��@	�-�e�3@�W��!?�X�5���@�q2�Пٿ��Y��@	�-�e�3@�W��!?�X�5���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�ӏ���ٿS���f�@�����3@k�Ұߐ!?���h���@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@�аgȡٿ?d�m�@��:K��3@��Ӑ!?6��� �@FW_�ŝٿA��1u�@w�c���3@�b�O��!?�r`ב��@FW_�ŝٿA��1u�@w�c���3@�b�O��!?�r`ב��@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@���f��ٿaŇ�@�_�Z��3@�8���!?��}Y���@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@�y0c�ٿ&;%���@ ����3@L��>q�!?�Ւ����@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@e��Q�ٿ�x�����@�G(�3@��V^�!?r8��a��@��v��ٿ+M��U��@-�Y{��3@�u%ߐ!?�f�`��@g��&��ٿ;nR=�K�@�Z#Ӹ�3@7���!?���n�@g��&��ٿ;nR=�K�@�Z#Ӹ�3@7���!?���n�@g��&��ٿ;nR=�K�@�Z#Ӹ�3@7���!?���n�@d���ٿ����|��@�#����3@q����!?D����@�@d���ٿ����|��@�#����3@q����!?D����@�@&���3�ٿ��C��@ȯ�}�3@�˄���!?�ן:�@&���3�ٿ��C��@ȯ�}�3@�˄���!?�ן:�@&���3�ٿ��C��@ȯ�}�3@�˄���!?�ן:�@�jy��ٿ���k�T�@V����3@vO r'�!?�|���/�@��G�j�ٿ�)į�w�@�M��3@�=JwÐ!?���<?��@��G�j�ٿ�)į�w�@�M��3@�=JwÐ!?���<?��@��G�j�ٿ�)į�w�@�M��3@�=JwÐ!?���<?��@��G�j�ٿ�)į�w�@�M��3@�=JwÐ!?���<?��@~[-�+�ٿ2�{�T��@��|��3@��e��!?Y��Y��@~[-�+�ٿ2�{�T��@��|��3@��e��!?Y��Y��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@4[����ٿ�F�%N�@��L��3@3��1��!?�*�-��@5Y�4�ٿ�g����@��#��3@ӌ��!?ؚJt�~�@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�HL��ٿ��)V��@u�y�[�3@�����!?p�����@�ۥ�ٿ-�|l7��@�xt���3@JҒ�!?X��3��@�ۥ�ٿ-�|l7��@�xt���3@JҒ�!?X��3��@�ۥ�ٿ-�|l7��@�xt���3@JҒ�!?X��3��@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@���2��ٿ�CP6���@�/����3@P�)Ő!?<��W�r�@Nz|�ٿ�VL���@�ٱx2�3@�8�Ԑ!?9!c��@��a��ٿ�5�"���@�w/Z�3@�i���!?�_xk�P�@��a��ٿ�5�"���@�w/Z�3@�i���!?�_xk�P�@����,�ٿ�l�2�@ -�>�3@�{H�`�!?�Z�V���@����,�ٿ�l�2�@ -�>�3@�{H�`�!?�Z�V���@����,�ٿ�l�2�@ -�>�3@�{H�`�!?�Z�V���@�Q"R.�ٿ�x?Ȉ��@��n6��3@b��a�!?&���P�@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@f�!�ٿ8^C����@�����3@i�◐!?t�GX��@���P�ٿF}R��@XSap��3@�Ӕg��!?�2�ܔ��@���P�ٿF}R��@XSap��3@�Ӕg��!?�2�ܔ��@7,d&$�ٿ&KV}��@�q��%�3@��=O��!?j6>���@ye��0�ٿ6eߒb>�@��1���3@�;�-�!?r�v��<�@ye��0�ٿ6eߒb>�@��1���3@�;�-�!?r�v��<�@�hW<=�ٿ!٦E�)�@fv����3@�:y1��!?
�v�Z�@�hW<=�ٿ!٦E�)�@fv����3@�:y1��!?
�v�Z�@�hW<=�ٿ!٦E�)�@fv����3@�:y1��!?
�v�Z�@hh���ٿ�ĘI��@T$�qx�3@��i���!?����p�@hh���ٿ�ĘI��@T$�qx�3@��i���!?����p�@hh���ٿ�ĘI��@T$�qx�3@��i���!?����p�@�|�@b�ٿ{I����@ӕ\�B�3@���!?�T��{B�@�|�@b�ٿ{I����@ӕ\�B�3@���!?�T��{B�@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@%�u��ٿ�S麲��@*F�{��3@�G����!?1��y��@˚9�ٿ- ʿ;|�@,v����3@~	�3w�!?��@���@��
Ǟٿd@#���@aSV���3@�C���!?xk��x��@��
Ǟٿd@#���@aSV���3@�C���!?xk��x��@%��d9�ٿƙJ���@U�����3@�����!?�9���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@��$ �ٿ	��{H��@P�V��3@���!�!?"��=���@����b�ٿ-:J��@���3@K��!?"��?��@����b�ٿ-:J��@���3@K��!?"��?��@����b�ٿ-:J��@���3@K��!?"��?��@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@eq�r�ٿ�NA⅖�@�����3@\q\X�!?u�<����@Zoo�B�ٿJa+@��@��w�3@��/#��!?�B����@Zoo�B�ٿJa+@��@��w�3@��/#��!?�B����@Zoo�B�ٿJa+@��@��w�3@��/#��!?�B����@l�s|4�ٿ�|8);�@��`��3@����o�!?����(�@l�s|4�ٿ�|8);�@��`��3@����o�!?����(�@l�s|4�ٿ�|8);�@��`��3@����o�!?����(�@�����ٿ5� ����@��no�3@�	��h�!?�����6�@��fx�ٿT�̛���@��\B��3@�@��l�!?D�i�:�@��fx�ٿT�̛���@��\B��3@�@��l�!?D�i�:�@��fx�ٿT�̛���@��\B��3@�@��l�!?D�i�:�@��fx�ٿT�̛���@��\B��3@�@��l�!?D�i�:�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@r�!"��ٿA�h���@:���C�3@�5�Ҥ�!?����9Q�@{z$,��ٿgLD���@��0��3@�!ŀ�!?�7�*J�@x+郛ٿqv�&@L�@�����3@sF�M�!?�ȡ�I�@�(�ٿ%�Q3���@� ���3@7�ζ�!?f�_Ԙ��@�(�ٿ%�Q3���@� ���3@7�ζ�!?f�_Ԙ��@�(�ٿ%�Q3���@� ���3@7�ζ�!?f�_Ԙ��@�(�ٿ%�Q3���@� ���3@7�ζ�!?f�_Ԙ��@�(�ٿ%�Q3���@� ���3@7�ζ�!?f�_Ԙ��@���2#�ٿ���*�@���+��3@��!��!?�-�����@���2#�ٿ���*�@���+��3@��!��!?�-�����@���2#�ٿ���*�@���+��3@��!��!?�-�����@���2#�ٿ���*�@���+��3@��!��!?�-�����@���2#�ٿ���*�@���+��3@��!��!?�-�����@��g��ٿ&�pp�@��3 �3@.Ng���!?��]y}�@��g��ٿ&�pp�@��3 �3@.Ng���!?��]y}�@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@\=G��ٿ�}M��<�@J?����3@Sh!?�ν�}��@�����ٿe�G���@�HV�3@BϮΐ!?���$��@�����ٿe�G���@�HV�3@BϮΐ!?���$��@�����ٿe�G���@�HV�3@BϮΐ!?���$��@��I�ʦٿZ�{3��@��!e�3@2�����!?�XOA\�@��I�ʦٿZ�{3��@��!e�3@2�����!?�XOA\�@��I�ʦٿZ�{3��@��!e�3@2�����!?�XOA\�@{}?�2�ٿ�/�cN�@�lc�a�3@�;<
��!?9�؎Y�@{}?�2�ٿ�/�cN�@�lc�a�3@�;<
��!?9�؎Y�@{}?�2�ٿ�/�cN�@�lc�a�3@�;<
��!?9�؎Y�@{}?�2�ٿ�/�cN�@�lc�a�3@�;<
��!?9�؎Y�@�����ٿ7A����@��
X`�3@�	*�!?�)�Rv��@�����ٿ7A����@��
X`�3@�	*�!?�)�Rv��@ڔ�'�ٿ���j&��@���	�3@�%VC�!?�kK$���@ڔ�'�ٿ���j&��@���	�3@�%VC�!?�kK$���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@=�bn�ٿ�T����@������3@N�7�Z�!?^Z���@��W.q�ٿt���'j�@/��A�3@a/wo.�!?>�c��@��W.q�ٿt���'j�@/��A�3@a/wo.�!?>�c��@B2�7-�ٿ�K:\�J�@�(�\�3@��O� �!?Ab�����@B2�7-�ٿ�K:\�J�@�(�\�3@��O� �!?Ab�����@*����ٿ UcU�F�@�{{�3@��]W�!?�(���@��e�ٿ�Ǥ4F��@��8�3@L�I�!?Y�����@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@kk�3��ٿS�^�q�@���b�3@U���Z�!?�an4��@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@��M���ٿ�������@�7d�n�3@5��f��!?�ы�:�@�ܧ��ٿ���;��@��wu�3@c\V���!?*:�9��@�ܧ��ٿ���;��@��wu�3@c\V���!?*:�9��@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@\;[X$�ٿ��U��@�F-��3@���-֐!?�xq���@�o���ٿ��V��/�@V��I��3@�X�<ΐ!?6!��J�@�o���ٿ��V��/�@V��I��3@�X�<ΐ!?6!��J�@�o���ٿ��V��/�@V��I��3@�X�<ΐ!?6!��J�@�o���ٿ��V��/�@V��I��3@�X�<ΐ!?6!��J�@�ؾp��ٿ�b~���@�����3@\�i���!?F�7GU�@�-z�^�ٿ�X%�<�@�0s{�3@�����!?��ERNj�@�-z�^�ٿ�X%�<�@�0s{�3@�����!?��ERNj�@�-z�^�ٿ�X%�<�@�0s{�3@�����!?��ERNj�@�-z�^�ٿ�X%�<�@�0s{�3@�����!?��ERNj�@M΅ϬٿԜUc�@�C܇�3@�0�A��!?�+��y��@M΅ϬٿԜUc�@�C܇�3@�0�A��!?�+��y��@M΅ϬٿԜUc�@�C܇�3@�0�A��!?�+��y��@M΅ϬٿԜUc�@�C܇�3@�0�A��!?�+��y��@�	i�ٿ�7x�z�@h����3@����!?^'��2�@�	i�ٿ�7x�z�@h����3@����!?^'��2�@W�N��ٿAw�5��@쩟���3@fw{�!?��a�w�@����ٿ��|��@�~����3@��k��!?ٶ�,�@����ٿ��|��@�~����3@��k��!?ٶ�,�@����ٿ��|��@�~����3@��k��!?ٶ�,�@����ٿ��|��@�~����3@��k��!?ٶ�,�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@�JUų�ٿ�m�g��@,zī��3@6y�ސ!?y�֏+�@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@`	���ٿ�ڈ���@�mJ���3@�zu��!?�'���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@.5���ٿ����P�@bq���3@
��	��!?��7���@�ߵ���ٿ��d���@ Dˏ]�3@c�(�!?��$2���@e�<e�ٿ���5��@RV���3@�M�K�!?��t�f��@e�<e�ٿ���5��@RV���3@�M�K�!?��t�f��@��G�ٿ-,����@'ǚq�3@3�i�!?�G�Y��@��G�ٿ-,����@'ǚq�3@3�i�!?�G�Y��@��D1�ٿ���2�{�@o�E �3@'�*,��!?5�ʉ��@��D1�ٿ���2�{�@o�E �3@'�*,��!?5�ʉ��@��D1�ٿ���2�{�@o�E �3@'�*,��!?5�ʉ��@��:��ٿ��ic��@I���3@��fļ�!?��b����@��:��ٿ��ic��@I���3@��fļ�!?��b����@j5�M�ٿ�$���:�@k�6�b�3@��|y��!?��1���@��=�ٿ���	�t�@À���3@���!?���˘�@T�Ŧפٿ�Dadʆ�@2��Jn�3@\LꟐ!?c�Fa��@T�Ŧפٿ�Dadʆ�@2��Jn�3@\LꟐ!?c�Fa��@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�]Ԥ��ٿ'�T��@.@����3@�a֯�!?~����@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@�vr>�ٿU�\��@��{�3@�4���!?��@�l��@CaǏΣٿ���Ae@�@( =��3@�ǡ�	�!?$��*�@��}�ٿ}��b��@]�T>�3@�]Bŭ�!?�	���@��}�ٿ}��b��@]�T>�3@�]Bŭ�!?�	���@��}�ٿ}��b��@]�T>�3@�]Bŭ�!?�	���@��}�ٿ}��b��@]�T>�3@�]Bŭ�!?�	���@�R�Lǡٿ�"R�2�@8ƽ��3@c��̐!?�3\�Q�@�R�Lǡٿ�"R�2�@8ƽ��3@c��̐!?�3\�Q�@�R�Lǡٿ�"R�2�@8ƽ��3@c��̐!?�3\�Q�@�R�Lǡٿ�"R�2�@8ƽ��3@c��̐!?�3\�Q�@�R�Lǡٿ�"R�2�@8ƽ��3@c��̐!?�3\�Q�@��j�ٿ�1�^�Z�@��5� �3@TشY
�!?i��)>�@��j�ٿ�1�^�Z�@��5� �3@TشY
�!?i��)>�@K�K�ٿ7���4y�@����3@t%>�!?Q��QHI�@K�K�ٿ7���4y�@����3@t%>�!?Q��QHI�@K�K�ٿ7���4y�@����3@t%>�!?Q��QHI�@K�K�ٿ7���4y�@����3@t%>�!?Q��QHI�@��=��ٿ{���}�@�N���3@L��99�!?���;��@��=��ٿ{���}�@�N���3@L��99�!?���;��@�����ٿ��sg�O�@k�ɴ�3@��4�!?d�J�R"�@�����ٿ��sg�O�@k�ɴ�3@��4�!?d�J�R"�@�����ٿ��sg�O�@k�ɴ�3@��4�!?d�J�R"�@� %P�ٿ8�Ru���@���ɉ�3@�{��1�!?�J�p���@� %P�ٿ8�Ru���@���ɉ�3@�{��1�!?�J�p���@�H۽�ٿCst`��@��{�U�3@.�E{��!?Ua���@�H۽�ٿCst`��@��{�U�3@.�E{��!?Ua���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@E`�˛ٿK:�*�w�@������3@T%��!?��}$���@T�� Ǟٿ��"D��@8
[�j�3@M\����!?��y@�*�@T�� Ǟٿ��"D��@8
[�j�3@M\����!?��y@�*�@T�� Ǟٿ��"D��@8
[�j�3@M\����!?��y@�*�@T�� Ǟٿ��"D��@8
[�j�3@M\����!?��y@�*�@T�� Ǟٿ��"D��@8
[�j�3@M\����!?��y@�*�@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@UGt�ٿ�u��y�@m�'���3@���h�!?�c; ��@Ah�]ԝٿٞ��k$�@*G���3@F�Yf��!?�C�N���@Ah�]ԝٿٞ��k$�@*G���3@F�Yf��!?�C�N���@Y��Υٿ�>���@�ቀ��3@�ɋ�y�!?�����@Y��Υٿ�>���@�ቀ��3@�ɋ�y�!?�����@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@'���͟ٿ����N_�@	��7�3@��Z��!?������@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�a)E�ٿ��'�@�KY��3@��ِ!?[�\��p�@�i�9�ٿ������@]���w�3@��5��!?�R&m�|�@�i�9�ٿ������@]���w�3@��5��!?�R&m�|�@�i�9�ٿ������@]���w�3@��5��!?�R&m�|�@�i�9�ٿ������@]���w�3@��5��!?�R&m�|�@�i�9�ٿ������@]���w�3@��5��!?�R&m�|�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�.M�7�ٿ�7Ab��@�-�+�3@R���Ґ!?���&ly�@�cIٞٿ4�2�@�0vv�3@)�����!?M�s|��@�cIٞٿ4�2�@�0vv�3@)�����!?M�s|��@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@�=kq�ٿ��ؽ\�@AY����3@$��8�!?ik�[K�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@>��@��ٿ�:�?&]�@=uTT\�3@I��8�!?s��2�@�	~���ٿ ��p���@��$��3@x�T��!?�ŉ��0�@�	~���ٿ ��p���@��$��3@x�T��!?�ŉ��0�@�	~���ٿ ��p���@��$��3@x�T��!?�ŉ��0�@�	~���ٿ ��p���@��$��3@x�T��!?�ŉ��0�@�ǜҝٿ�`���@��'E��3@��Lj�!?�l���s�@�ǜҝٿ�`���@��'E��3@��Lj�!?�l���s�@�ǜҝٿ�`���@��'E��3@��Lj�!?�l���s�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@�p��ٿn��U��@����3@���!?�N��^�@7��Sd�ٿ|Moy*�@��X��3@ԣ;���!?E��0ͼ�@7��Sd�ٿ|Moy*�@��X��3@ԣ;���!?E��0ͼ�@7��Sd�ٿ|Moy*�@��X��3@ԣ;���!?E��0ͼ�@7��Sd�ٿ|Moy*�@��X��3@ԣ;���!?E��0ͼ�@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@��'��ٿ��៑�@�T�M��3@q�i�!?�q�M���@������ٿdwM��@����3@�>���!?r��?��@������ٿdwM��@����3@�>���!?r��?��@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@Z_�G��ٿ�elB��@�Ru[�3@);��͐!?�,����@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@�*`N��ٿ`gŕ�@��muK�3@���!?��OLɒ�@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@oG=3��ٿ����@ ���3@�B1��!?0զ��@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@���ɸ�ٿ��|����@|�]=��3@�n_�!?��x���@h�r��ٿ��C�� �@3Q�z��3@:�ېא!?��T�D��@h�r��ٿ��C�� �@3Q�z��3@:�ېא!?��T�D��@h�r��ٿ��C�� �@3Q�z��3@:�ېא!?��T�D��@����Λٿs�n���@���'�3@��[�ϐ!?i5n߿�@_z7b5�ٿ��U�� �@%󉍕�3@��j�Đ!?���'���@�� A�ٿ��3��@E���3@F�sYԐ!?��I¬I�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@2���Y�ٿ!��P���@���m�3@7д��!?���6�@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@_�e6�ٿ}���@x��g�3@�\� �!?TA8u��@I��i�ٿ�32���@�g
Q�3@�h)�
�!?�zE�W'�@��p�g�ٿ�Ĥ֦��@A�\�3@� �+̐!?�l����@�qf�R�ٿ������@�y{+�3@3 Q]��!?��x/Eg�@�qf�R�ٿ������@�y{+�3@3 Q]��!?��x/Eg�@�v�ěٿh���e�@�I�*��3@M ����!?R@�#��@�v�ěٿh���e�@�I�*��3@M ����!?R@�#��@�v�ěٿh���e�@�I�*��3@M ����!?R@�#��@�v�ěٿh���e�@�I�*��3@M ����!?R@�#��@�S�|�ٿ�p>xܲ�@nq����3@�lt�!?�ď ��@�S�|�ٿ�p>xܲ�@nq����3@�lt�!?�ď ��@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@��F���ٿ�	Ut��@�����3@2+1��!?+�E ?B�@%v�_�ٿqV��m7�@����6�3@X{���!?�����@%v�_�ٿqV��m7�@����6�3@X{���!?�����@%v�_�ٿqV��m7�@����6�3@X{���!?�����@���a��ٿN�w�{��@�I�q�3@n`��!?'r��%��@���a��ٿN�w�{��@�I�q�3@n`��!?'r��%��@��l��ٿ�4��d�@ X�/�3@����!?�Mj���@}��1��ٿ<)�uN�@C=��]�3@r_R6�!?.�����@}��1��ٿ<)�uN�@C=��]�3@r_R6�!?.�����@O#jw��ٿ@�t���@��\(��3@�__@�!?6�sD��@O#jw��ٿ@�t���@��\(��3@�__@�!?6�sD��@n!�fZ�ٿ�=���@s4����3@��Qv��!?��*ԟ�@n!�fZ�ٿ�=���@s4����3@��Qv��!?��*ԟ�@n!�fZ�ٿ�=���@s4����3@��Qv��!?��*ԟ�@AF	�ٿ����@�#�
��3@�!:А!?��PI�3�@AF	�ٿ����@�#�
��3@�!:А!?��PI�3�@AF	�ٿ����@�#�
��3@�!:А!?��PI�3�@AF	�ٿ����@�#�
��3@�!:А!?��PI�3�@L,�8u�ٿ��#��@����3@NRZo��!?6�Aԩ6�@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@@@TK�ٿ���<��@%F���3@�>�Đ!?F������@Һ�n�ٿ��cv��@�/ޫ��3@��/'��!?,g���@Һ�n�ٿ��cv��@�/ޫ��3@��/'��!?,g���@Һ�n�ٿ��cv��@�/ޫ��3@��/'��!?,g���@Һ�n�ٿ��cv��@�/ޫ��3@��/'��!?,g���@Һ�n�ٿ��cv��@�/ޫ��3@��/'��!?,g���@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@4��.ݤٿm�q���@�&W��3@�e���!?�{̇F{�@�Y�̢ٿ����`s�@�E�>#�3@��;��!?��(���@�Y�̢ٿ����`s�@�E�>#�3@��;��!?��(���@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@)�9yT�ٿ~�����@Zsy ��3@,��ݐ!?vJ��@ct���ٿ�V�U�@z@"S}�3@���S�!?�� ~��@ct���ٿ�V�U�@z@"S}�3@���S�!?�� ~��@ct���ٿ�V�U�@z@"S}�3@���S�!?�� ~��@ct���ٿ�V�U�@z@"S}�3@���S�!?�� ~��@�A`GŚٿ�&���I�@�PW�F�3@��A��!?e�'�v��@�A`GŚٿ�&���I�@�PW�F�3@��A��!?e�'�v��@�A`GŚٿ�&���I�@�PW�F�3@��A��!?e�'�v��@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@唇[��ٿN@&��@��`���3@�6O�!?��t���@*��T�ٿ���`�@狺��3@���!?�_����@D�Z��ٿ8�����@����i�3@�T"��!?�|`7�i�@D�Z��ٿ8�����@����i�3@�T"��!?�|`7�i�@D�Z��ٿ8�����@����i�3@�T"��!?�|`7�i�@D�Z��ٿ8�����@����i�3@�T"��!?�|`7�i�@����ٿ�ˋ�2�@쩿x�3@σ�EԐ!?�����@����ٿ�ˋ�2�@쩿x�3@σ�EԐ!?�����@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@�|�'͝ٿoy��3��@@�ܕ��3@>X�3��!?��Z@��@]��B�ٿ+z��k�@.et��3@���N�!?:��r��@]��B�ٿ+z��k�@.et��3@���N�!?:��r��@v�>Ȁ�ٿ�@V}�h�@Oi�E�3@s�2#��!?�X3P5S�@v�>Ȁ�ٿ�@V}�h�@Oi�E�3@s�2#��!?�X3P5S�@v�>Ȁ�ٿ�@V}�h�@Oi�E�3@s�2#��!?�X3P5S�@R�~ު�ٿYq5�=��@W�����3@��%��!?�J�����@R�~ު�ٿYq5�=��@W�����3@��%��!?�J�����@�o��\�ٿs��~�Y�@�j
G�3@���ϐ!?������@k�vo��ٿI�L�@��W��3@��j��!?�j����@k�vo��ٿI�L�@��W��3@��j��!?�j����@k�vo��ٿI�L�@��W��3@��j��!?�j����@Y�Z��ٿ�_��{b�@�3W���3@�����!?V/��3��@Y�Z��ٿ�_��{b�@�3W���3@�����!?V/��3��@Y�Z��ٿ�_��{b�@�3W���3@�����!?V/��3��@�mQ��ٿ7�9#|��@�+A���3@o�o;��!?��=BK�@�mQ��ٿ7�9#|��@�+A���3@o�o;��!?��=BK�@��>Y�ٿ[��VY�@���T~�3@A�ce��!?	=����@��>Y�ٿ[��VY�@���T~�3@A�ce��!?	=����@��>Y�ٿ[��VY�@���T~�3@A�ce��!?	=����@|�%c
�ٿ�p��;�@A����3@����y�!?��/��@|�%c
�ٿ�p��;�@A����3@����y�!?��/��@|�%c
�ٿ�p��;�@A����3@����y�!?��/��@|�%c
�ٿ�p��;�@A����3@����y�!?��/��@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@Q����ٿK�Q��[�@�s���3@L-A�r�!?�bUM���@��g��ٿ��u���@i����3@�$'���!?]ĸ߃��@��g��ٿ��u���@i����3@�$'���!?]ĸ߃��@��q�ٿ�)��(�@�/; J�3@���;��!?��N�_c�@��q�ٿ�)��(�@�/; J�3@���;��!?��N�_c�@��q�ٿ�)��(�@�/; J�3@���;��!?��N�_c�@��q�ٿ�)��(�@�/; J�3@���;��!?��N�_c�@��q�ٿ�)��(�@�/; J�3@���;��!?��N�_c�@���_ϧٿu��nS�@��6�3@cJK@`�!?���Rb�@���_ϧٿu��nS�@��6�3@cJK@`�!?���Rb�@�KpVz�ٿg:�H�@,�ز%�3@i���>�!?�!J��@�F�㈡ٿ��s�{��@��s)�3@�媗|�!?�"z�#M�@���"P�ٿl�i���@�m�Х�3@6(~b��!?���~v�@���"P�ٿl�i���@�m�Х�3@6(~b��!?���~v�@���"P�ٿl�i���@�m�Х�3@6(~b��!?���~v�@�I�/�ٿ�,���@2%�3@�k�[�!?GYo�t3�@y�'�ٿ�� �^��@�����3@uY>d��!?�����@y�'�ٿ�� �^��@�����3@uY>d��!?�����@y�'�ٿ�� �^��@�����3@uY>d��!?�����@y�'�ٿ�� �^��@�����3@uY>d��!?�����@y�'�ٿ�� �^��@�����3@uY>d��!?�����@� ��L�ٿޭDy�a�@����3@�Ͼ ��!?&�y&���@� ��L�ٿޭDy�a�@����3@�Ͼ ��!?&�y&���@� ��L�ٿޭDy�a�@����3@�Ͼ ��!?&�y&���@� ��L�ٿޭDy�a�@����3@�Ͼ ��!?&�y&���@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@�O��ٿ,�� �7�@�	<I�3@\͕�ܐ!?�F����@nmݠٿ�z����@�Ɩ�'�3@���Z͐!?ǻkMF��@\�<��ٿ"���o��@��];�3@��p(��!?]�1z��@\�<��ٿ"���o��@��];�3@��p(��!?]�1z��@�R�Y^�ٿ�Y���h�@�o����3@f
��!�!?�y��s�@�R�Y^�ٿ�Y���h�@�o����3@f
��!�!?�y��s�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@�O����ٿf�҃�D�@���/��3@!�x֐!?s�@�E�@��8�ٿ�����@���>�3@���ߐ!?:���z�@��8�ٿ�����@���>�3@���ߐ!?:���z�@�B␝ٿLd6�e"�@hU����3@���q��!? ���ې�@�B␝ٿLd6�e"�@hU����3@���q��!? ���ې�@�B␝ٿLd6�e"�@hU����3@���q��!? ���ې�@�/�?�ٿ��^��@�cr�3@��xh��!?�O����@�/�?�ٿ��^��@�cr�3@��xh��!?�O����@ z�W�ٿ:.w���@�*�w�3@y)1�l�!?���#�@ z�W�ٿ:.w���@�*�w�3@y)1�l�!?���#�@ z�W�ٿ:.w���@�*�w�3@y)1�l�!?���#�@i�aK�ٿ{��@�&�H��3@K�_{�!?�ւ-&-�@i�aK�ٿ{��@�&�H��3@K�_{�!?�ւ-&-�@i�aK�ٿ{��@�&�H��3@K�_{�!?�ւ-&-�@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@c��ٿ8�2q�@x�����3@�� ː!?�s�K��@4�� �ٿ\��Rq�@V��WR�3@S7K7��!?�l^�A�@4�� �ٿ\��Rq�@V��WR�3@S7K7��!?�l^�A�@4�� �ٿ\��Rq�@V��WR�3@S7K7��!?�l^�A�@+���ϧٿ/*oUY^�@}I+�v�3@j�44\�!?Q�����@z�@���ٿ.sI^D��@l�2��3@-\MY�!?���h���@z�@���ٿ.sI^D��@l�2��3@-\MY�!?���h���@{�Σٿ})<�*��@�;����3@m4��w�!?��T|��@{�Σٿ})<�*��@�;����3@m4��w�!?��T|��@J{hbj�ٿ(��tQ��@V ���3@F>3�:�!?KL�S��@J{hbj�ٿ(��tQ��@V ���3@F>3�:�!?KL�S��@J{hbj�ٿ(��tQ��@V ���3@F>3�:�!?KL�S��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@���~/�ٿV(�Z}�@�ٖ*8�3@���i�!?5�$ڊ��@`��zޣٿ2��r�3�@�7j��3@*[풐!?�=��J�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@6\���ٿһ�pS�@�X�o�3@p��r��!?};�0Z�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@a���ٿ#���
��@B�P��3@��D��!?q-��B�@�{|�ٿ~��G��@"�����3@�bā�!?�ڛl�@�{|�ٿ~��G��@"�����3@�bā�!?�ڛl�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@�����ٿ��}i�@*B{7�3@Ԉ�F�!?!z�w�@,V�ڞٿs�׍�#�@+bP��3@`��u�!?����4��@,V�ڞٿs�׍�#�@+bP��3@`��u�!?����4��@,V�ڞٿs�׍�#�@+bP��3@`��u�!?����4��@,V�ڞٿs�׍�#�@+bP��3@`��u�!?����4��@,V�ڞٿs�׍�#�@+bP��3@`��u�!?����4��@���~��ٿ��ܒ��@4�l'��3@|����!?�"F�
��@���~��ٿ��ܒ��@4�l'��3@|����!?�"F�
��@���~��ٿ��ܒ��@4�l'��3@|����!?�"F�
��@�!��ٿ�{���@�a^c�3@��|Ð!?T����@�!��ٿ�{���@�a^c�3@��|Ð!?T����@�!��ٿ�{���@�a^c�3@��|Ð!?T����@�!��ٿ�{���@�a^c�3@��|Ð!?T����@�!��ٿ�{���@�a^c�3@��|Ð!?T����@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@��[�ٿ���I��@���2�3@%lx�ސ!?yķ���@y�[:�ٿ��3���@P�"��3@�n�2�!?H�~�]�@y�[:�ٿ��3���@P�"��3@�n�2�!?H�~�]�@y�[:�ٿ��3���@P�"��3@�n�2�!?H�~�]�@y�[:�ٿ��3���@P�"��3@�n�2�!?H�~�]�@6�s�ٿ�)�1S�@�����3@6�b��!?�E ~���@6�s�ٿ�)�1S�@�����3@6�b��!?�E ~���@6�s�ٿ�)�1S�@�����3@6�b��!?�E ~���@6�s�ٿ�)�1S�@�����3@6�b��!?�E ~���@G�		�ٿv6�[kr�@��l��3@HgdӐ!?]`�@G�		�ٿv6�[kr�@��l��3@HgdӐ!?]`�@G�		�ٿv6�[kr�@��l��3@HgdӐ!?]`�@G�		�ٿv6�[kr�@��l��3@HgdӐ!?]`�@��L�ٿ���BzP�@;�ZX��3@u ݿ�!?��I�b�@! Зv�ٿ�EJ��@ϔ z��3@� }���!?u�kfW�@! Зv�ٿ�EJ��@ϔ z��3@� }���!?u�kfW�@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@*��r�ٿ�n #�@�ol��3@�y&���!?u��?��@N�-vQ�ٿ�{�};�@� ���3@��ϐ!?��i_��@N�-vQ�ٿ�{�};�@� ���3@��ϐ!?��i_��@N�-vQ�ٿ�{�};�@� ���3@��ϐ!?��i_��@N�-vQ�ٿ�{�};�@� ���3@��ϐ!?��i_��@N�-vQ�ٿ�{�};�@� ���3@��ϐ!?��i_��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@����ٿ�Т6��@>���'�3@���筐!?&�Jt��@	y��{�ٿgQ�KY��@T���3@�[G��!?lr�����@�X%$f�ٿ�B8�M��@�W���3@K�����!?@O����@8�m��ٿ�>�Y�@�c��3@�,Gν�!?Z
��t��@��,���ٿ:����@u�`�L�3@���!?HZYu��@��,���ٿ:����@u�`�L�3@���!?HZYu��@��,���ٿ:����@u�`�L�3@���!?HZYu��@F����ٿ��t��&�@�w+���3@[	aQ4�!?{�'G��@F����ٿ��t��&�@�w+���3@[	aQ4�!?{�'G��@��C�W�ٿ�C� 	H�@S���3@A$�!?���d@��@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@��[u�ٿ��v"���@�|���3@z���֐!?s�@���@�
A��ٿ��%��]�@<ε�g�3@,�X��!?65���6�@�
A��ٿ��%��]�@<ε�g�3@,�X��!?65���6�@Sr�ߤٿR��C^=�@b��w��3@��h��!?+=[c&�@Sr�ߤٿR��C^=�@b��w��3@��h��!?+=[c&�@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@�ߋ��ٿg!.j��@��F���3@B� ��!?������@R�#�r�ٿ�W��4�@�ק]D�3@�>ؐ!?�On���@��7��ٿ7!Q+�I�@�����3@��J�
�!?�4����@��7��ٿ7!Q+�I�@�����3@��J�
�!?�4����@(zʦ�ٿTW�-�@o5m#��3@���̐!?,7�-g��@(zʦ�ٿTW�-�@o5m#��3@���̐!?,7�-g��@(zʦ�ٿTW�-�@o5m#��3@���̐!?,7�-g��@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@ROX���ٿ��Z�+�@�J���3@�4^���!?ͤNH���@����[�ٿn4����@E�b��3@'��,�!? 8��.�@����[�ٿn4����@E�b��3@'��,�!? 8��.�@����[�ٿn4����@E�b��3@'��,�!? 8��.�@����[�ٿn4����@E�b��3@'��,�!? 8��.�@"k���ٿ}�y/���@a�rz`�3@@hM!��!?)VA�}�@"k���ٿ}�y/���@a�rz`�3@@hM!��!?)VA�}�@����ٿn-\��@��F��3@-����!?2�VOG��@����ٿn-\��@��F��3@-����!?2�VOG��@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@�e�R�ٿ��}���@��R�3@&�?;�!?��S�@{\yy�ٿiRŧ��@�F��3@t�qH<�!?�z�7F��@ʳ5�ٿo���@���H��3@n�� �!?�#��{�@ʳ5�ٿo���@���H��3@n�� �!?�#��{�@�QxU�ٿ�� �%�@y�����3@[k�@�!?����_�@,4ae�ٿn�ߢ���@yx�� �3@�|�Ö�!?}d7�@�@,4ae�ٿn�ߢ���@yx�� �3@�|�Ö�!?}d7�@�@,4ae�ٿn�ߢ���@yx�� �3@�|�Ö�!?}d7�@�@,4ae�ٿn�ߢ���@yx�� �3@�|�Ö�!?}d7�@�@?[X��ٿ�x�鐯�@�nV���3@=�d�!?sr��q�@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�����ٿ��p׊�@�9V�f�3@h�8 !�!?4y ���@�CZjԥٿ��JRQ�@cq�cx�3@��	}�!?����h��@�CZjԥٿ��JRQ�@cq�cx�3@��	}�!?����h��@�CZjԥٿ��JRQ�@cq�cx�3@��	}�!?����h��@�CZjԥٿ��JRQ�@cq�cx�3@��	}�!?����h��@�CZjԥٿ��JRQ�@cq�cx�3@��	}�!?����h��@�S2xءٿފ��|�@O9�(��3@�%Gʐ!?Ib��6�@�S2xءٿފ��|�@O9�(��3@�%Gʐ!?Ib��6�@�S2xءٿފ��|�@O9�(��3@�%Gʐ!?Ib��6�@�S2xءٿފ��|�@O9�(��3@�%Gʐ!?Ib��6�@�ƾ��ٿjw���@1�83J�3@����א!?���|1��@�ƾ��ٿjw���@1�83J�3@����א!?���|1��@P��8�ٿb��TG[�@<�P�3@o3���!?�����@P��8�ٿb��TG[�@<�P�3@o3���!?�����@V���
�ٿ�؈���@��o-�3@ŏj]�!?���En��@V���
�ٿ�؈���@��o-�3@ŏj]�!?���En��@V���
�ٿ�؈���@��o-�3@ŏj]�!?���En��@�u��ٿ�L_Cj�@�d�j��3@Ш=�+�!?O^Neb8�@�u��ٿ�L_Cj�@�d�j��3@Ш=�+�!?O^Neb8�@�u��ٿ�L_Cj�@�d�j��3@Ш=�+�!?O^Neb8�@ߓ<�,�ٿe7CNq�@%���,�3@�?٫��!?�W*�Z��@ߓ<�,�ٿe7CNq�@%���,�3@�?٫��!?�W*�Z��@ߓ<�,�ٿe7CNq�@%���,�3@�?٫��!?�W*�Z��@ߓ<�,�ٿe7CNq�@%���,�3@�?٫��!?�W*�Z��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@�}��e�ٿ�bHY��@��y��3@HQ��_�!?>d�4��@��"�ܣٿRȯ׳]�@0���3@�����!?�5;I`�@��"�ܣٿRȯ׳]�@0���3@�����!?�5;I`�@��"�ܣٿRȯ׳]�@0���3@�����!?�5;I`�@��"�ܣٿRȯ׳]�@0���3@�����!?�5;I`�@��"�ܣٿRȯ׳]�@0���3@�����!?�5;I`�@
m1��ٿ��B�Q�@d�]�3@�&���!?�3��A$�@��6�K�ٿ�E��h�@���c;�3@B
�n�!?�bʠ�^�@B�h�ٿqH��@"M�3@֖���!?Ƶ�;�@B�h�ٿqH��@"M�3@֖���!?Ƶ�;�@B�h�ٿqH��@"M�3@֖���!?Ƶ�;�@'t�&�ٿAeK!��@���X�3@[�0�!?i	-��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@�<n%�ٿ���	�C�@(�-�z�3@nvӐ!?Gխ.9��@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@%Ӆ���ٿ�TzQ�@徜ľ�3@Qq�q��!?�����m�@��f���ٿ�~�s��@"�#p�3@W�ҏ�!?q0��
�@��f���ٿ�~�s��@"�#p�3@W�ҏ�!?q0��
�@y˯���ٿzd����@�9`��3@�ڡ��!?��LK�
�@y˯���ٿzd����@�9`��3@�ڡ��!?��LK�
�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@���Y�ٿ�W ��@�Eh�3@�8ǐ!?S���$�@lT?��ٿw��"��@�Me��3@������!?��JN;��@lT?��ٿw��"��@�Me��3@������!?��JN;��@lT?��ٿw��"��@�Me��3@������!?��JN;��@����ٿvE���@�0ؚ�3@t�5ڐ!?���
�@����ٿvE���@�0ؚ�3@t�5ڐ!?���
�@����ٿvE���@�0ؚ�3@t�5ڐ!?���
�@����ٿvE���@�0ؚ�3@t�5ڐ!?���
�@O���7�ٿ"8>�u��@ˉ����3@����!?ͬy�W�@O���7�ٿ"8>�u��@ˉ����3@����!?ͬy�W�@O���7�ٿ"8>�u��@ˉ����3@����!?ͬy�W�@O���7�ٿ"8>�u��@ˉ����3@����!?ͬy�W�@O���7�ٿ"8>�u��@ˉ����3@����!?ͬy�W�@O���ٿ��D���@�MW�L�3@ԕ{i�!?I�,����@��E�ٿ�j��c�@'!&(�3@�B�Ր!?y��z�@g'#(�ٿ^�%���@�Br�3@�&���!?���#�@g'#(�ٿ^�%���@�Br�3@�&���!?���#�@g'#(�ٿ^�%���@�Br�3@�&���!?���#�@�3�u��ٿ���m<�@�\G���3@Ж���!?�d����@]Y��ޜٿ,��v�@ag]��3@Mu��_�!?���@X�+�ٿ6r�Л�@��*�p�3@d��,W�!?������@X�+�ٿ6r�Л�@��*�p�3@d��,W�!?������@X�+�ٿ6r�Л�@��*�p�3@d��,W�!?������@��C��ٿ�$F��q�@3����3@�^\��!?`�-I�h�@�8��ٿ�O �P��@����3@*�͢��!?��w���@�8��ٿ�O �P��@����3@*�͢��!?��w���@�8��ٿ�O �P��@����3@*�͢��!?��w���@�8��ٿ�O �P��@����3@*�͢��!?��w���@�8��ٿ�O �P��@����3@*�͢��!?��w���@�8��ٿ�O �P��@����3@*�͢��!?��w���@Zٖ��ٿ�݅w���@���	��3@�^��k�!?~eoA]*�@Zٖ��ٿ�݅w���@���	��3@�^��k�!?~eoA]*�@Zٖ��ٿ�݅w���@���	��3@�^��k�!?~eoA]*�@/iI�R�ٿ��E���@�mU��3@?�[Ӂ�!?b8<�H�@/iI�R�ٿ��E���@�mU��3@?�[Ӂ�!?b8<�H�@/iI�R�ٿ��E���@�mU��3@?�[Ӂ�!?b8<�H�@jL��ٿab��!��@��B�T�3@?���!?/�@jL��ٿab��!��@��B�T�3@?���!?/�@jL��ٿab��!��@��B�T�3@?���!?/�@jL��ٿab��!��@��B�T�3@?���!?/�@V!뵨ٿ�	���@?���3@DK���!?����D�@V!뵨ٿ�	���@?���3@DK���!?����D�@V!뵨ٿ�	���@?���3@DK���!?����D�@V!뵨ٿ�	���@?���3@DK���!?����D�@V!뵨ٿ�	���@?���3@DK���!?����D�@V!뵨ٿ�	���@?���3@DK���!?����D�@��F��ٿ�3Ɏ�+�@\D�M�3@h��'�!?H�����@��F��ٿ�3Ɏ�+�@\D�M�3@h��'�!?H�����@��F��ٿ�3Ɏ�+�@\D�M�3@h��'�!?H�����@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@��/t[�ٿ_�[bu�@�َ{�3@�}1+�!?�1�RA�@?�{�v�ٿ����b�@�Բ}E�3@�� 	�!?����j�@?�{�v�ٿ����b�@�Բ}E�3@�� 	�!?����j�@?�{�v�ٿ����b�@�Բ}E�3@�� 	�!?����j�@?�{�v�ٿ����b�@�Բ}E�3@�� 	�!?����j�@?�{�v�ٿ����b�@�Բ}E�3@�� 	�!?����j�@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�^&Uؤٿ��c��_�@�����3@�9�bؐ!?��w��@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@�r/\+�ٿY�Ǽk��@���)�3@�L����!?�LQ���@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@��y���ٿ�E���@OtH1�3@���[Ր!?�S����@���H��ٿ����h��@��G��3@��RṐ!?~	����@s`nH��ٿU��(c��@i�5c��3@�+p��!?�k�h��@s`nH��ٿU��(c��@i�5c��3@�+p��!?�k�h��@s`nH��ٿU��(c��@i�5c��3@�+p��!?�k�h��@�e�\O�ٿB�<���@�eXdF�3@M�ƛ�!?n���e�@�;^AK�ٿ3]����@%�d:l�3@2DѶx�!?j?bM���@�;^AK�ٿ3]����@%�d:l�3@2DѶx�!?j?bM���@��4��ٿJ�:K��@��f�h�3@F��ʥ�!?UB��3��@��4��ٿJ�:K��@��f�h�3@F��ʥ�!?UB��3��@�G��ٿ�4�Kp�@��a�s�3@���晐!?dt�:l��@�G��ٿ�4�Kp�@��a�s�3@���晐!?dt�:l��@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@
�K���ٿF�^�\�@�G��/�3@�����!?��s�2�@�yr�v�ٿ�J��y�@�2�US�3@�R�6��!?�����@�yr�v�ٿ�J��y�@�2�US�3@�R�6��!?�����@�yr�v�ٿ�J��y�@�2�US�3@�R�6��!?�����@�yr�v�ٿ�J��y�@�2�US�3@�R�6��!?�����@�yr�v�ٿ�J��y�@�2�US�3@�R�6��!?�����@���
�ٿ}b}�[�@��T��3@���ݐ!?Ŗ~�+��@���
�ٿ}b}�[�@��T��3@���ݐ!?Ŗ~�+��@���
�ٿ}b}�[�@��T��3@���ݐ!?Ŗ~�+��@���
�ٿ}b}�[�@��T��3@���ݐ!?Ŗ~�+��@���
�ٿ}b}�[�@��T��3@���ݐ!?Ŗ~�+��@��#��ٿ������@,f����3@�12��!?�tO� �@��#��ٿ������@,f����3@�12��!?�tO� �@��#��ٿ������@,f����3@�12��!?�tO� �@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@C�*T��ٿugs���@�t�}4@Q7\Ȑ!?���՝��@�$�x
�ٿה]�'��@��rJ��3@R��Ő!?g�`�IR�@�$�x
�ٿה]�'��@��rJ��3@R��Ő!?g�`�IR�@�$Q�ٿ�����a�@Tw�5�3@��=�!?�/*4���@�$Q�ٿ�����a�@Tw�5�3@��=�!?�/*4���@�$Q�ٿ�����a�@Tw�5�3@��=�!?�/*4���@�$Q�ٿ�����a�@Tw�5�3@��=�!?�/*4���@�O����ٿQl2u��@��ʎl�3@��0�!?�;3U���@�O����ٿQl2u��@��ʎl�3@��0�!?�;3U���@�O����ٿQl2u��@��ʎl�3@��0�!?�;3U���@�:۵��ٿH�:�R��@�����3@l����!?ë�%I�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@���L�ٿ-�4/��@����3@t���!?!��ˬ�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@����n�ٿ�Pf��@V��p�3@r�r��!?���tj�@o�A{�ٿk#E<��@�w�,��3@'��M�!?�=%���@o�A{�ٿk#E<��@�w�,��3@'��M�!?�=%���@o�A{�ٿk#E<��@�w�,��3@'��M�!?�=%���@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@��A	v�ٿ~�?�Pj�@�Ӈa�3@���֐!?Pu0j�@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@D	[v�ٿ���A�@ks]��3@i���ې!?��`��@.�@�ٿ-7Y���@��d��3@��:R�!?�]�|��@���J��ٿ�H�����@�����3@ �^c�!?��[�B��@���J��ٿ�H�����@�����3@ �^c�!?��[�B��@��>DS�ٿh�:+A�@=sh�3@+�ﮩ�!?WG�e�@��>DS�ٿh�:+A�@=sh�3@+�ﮩ�!?WG�e�@��>DS�ٿh�:+A�@=sh�3@+�ﮩ�!?WG�e�@��>DS�ٿh�:+A�@=sh�3@+�ﮩ�!?WG�e�@��>DS�ٿh�:+A�@=sh�3@+�ﮩ�!?WG�e�@Nt�	G�ٿZEt���@��.}�3@��=��!?Z�[�H�@Nt�	G�ٿZEt���@��.}�3@��=��!?Z�[�H�@�D�f֚ٿm��,OH�@�)'�3@:�afY�!?��V���@�D�f֚ٿm��,OH�@�)'�3@:�afY�!?��V���@����ٿI���ʀ�@�rW�o�3@��C�^�!?Is!X��@����ٿI���ʀ�@�rW�o�3@��C�^�!?Is!X��@k��'�ٿ��'9�@uο_k�3@��qR�!?yso���@k��'�ٿ��'9�@uο_k�3@��qR�!?yso���@�$��ٿ��"c��@��y�t 4@Y�K_Đ!?���QK�@�$��ٿ��"c��@��y�t 4@Y�K_Đ!?���QK�@�$��ٿ��"c��@��y�t 4@Y�K_Đ!?���QK�@KE��ٿ�gY�I�@��%7�3@�f~�!?Z$��0��@Հ׺�ٿ�}�X�@V[
��3@�AA�ސ!?�#�^(��@ٶ:�ٿ�0p����@MT$4��3@-u���!?��{�+�@ٶ:�ٿ�0p����@MT$4��3@-u���!?��{�+�@����o�ٿ�(�s���@g���'�3@g�/͐!?_e�E_�@E<>�ٿ����X9�@��n%�3@>���!?l����Z�@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@*/b�ģٿ�\��G��@�,�Z�3@ i�]��!?�x�M��@@�đ�ٿ��-��@'�>�3@��]�!?��1�s��@@�đ�ٿ��-��@'�>�3@��]�!?��1�s��@@�đ�ٿ��-��@'�>�3@��]�!?��1�s��@@�đ�ٿ��-��@'�>�3@��]�!?��1�s��@@�đ�ٿ��-��@'�>�3@��]�!?��1�s��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@���CV�ٿmR5��@<����3@�"+�!?�;��-��@.O�� �ٿ�	�dsu�@�Zz�l�3@+㟪�!?g��M���@.O�� �ٿ�	�dsu�@�Zz�l�3@+㟪�!?g��M���@.O�� �ٿ�	�dsu�@�Zz�l�3@+㟪�!?g��M���@.O�� �ٿ�	�dsu�@�Zz�l�3@+㟪�!?g��M���@.O�� �ٿ�	�dsu�@�Zz�l�3@+㟪�!?g��M���@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��P�;�ٿ1KO��|�@]��TO�3@ub�N�!?͓���u�@��e\��ٿ7V
ov�@U1�x�3@������!? �Ӵ�5�@��e\��ٿ7V
ov�@U1�x�3@������!? �Ӵ�5�@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@)N�x�ٿ����L��@��-�3@�!�A�!?��u����@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@j��E�ٿ"k�7�P�@;
L	&�3@*�j�Đ!?�{#� ��@�j��ٿ3oSj�}�@��:T�3@#`㜠�!?��T�o�@��][�ٿB��{a��@��A+��3@�9�w�!?M��%|��@��][�ٿB��{a��@��A+��3@�9�w�!?M��%|��@��][�ٿB��{a��@��A+��3@�9�w�!?M��%|��@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@� ǝ[�ٿ�O��@�,i���3@?﹬ΐ!?j�w���@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@x�򮘕ٿ�����\�@@K?��3@ae�C��!?�0��z�@&��ٿ�ز5���@������3@^"%qp�!?=葸�O�@P/��Қٿg<�nc�@�T$~��3@��N�G�!?,5<��@P/��Қٿg<�nc�@�T$~��3@��N�G�!?,5<��@P/��Қٿg<�nc�@�T$~��3@��N�G�!?,5<��@P/��Қٿg<�nc�@�T$~��3@��N�G�!?,5<��@P/��Қٿg<�nc�@�T$~��3@��N�G�!?,5<��@W���v�ٿAb ����@V�oj)�3@av�U=�!?z:?<��@W���v�ٿAb ����@V�oj)�3@av�U=�!?z:?<��@���4j�ٿEJ��0�@�� ��3@��G�!?+��$d��@�˝R
�ٿ�Ӧ����@��Nq. 4@�D��S�!?B���EY�@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@n9��k�ٿ�z	(�@w��N�3@�~�s�!?,����@
�����ٿmԄx�y�@f����3@O����!?��n���@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@O�fʥٿ̎�P� �@IE6��3@��Î�!?�>����@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@Ҋ+�ٿ�3 ~�f�@Mz]���3@T���!?�^s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@g�8��ٿ���b��@���&��3@�ok,�!?�4.�s��@�*�jɘٿl�t0���@"բ�j�3@��/�!?P'	.�@�*�jɘٿl�t0���@"բ�j�3@��/�!?P'	.�@�*�jɘٿl�t0���@"բ�j�3@��/�!?P'	.�@�*�jɘٿl�t0���@"բ�j�3@��/�!?P'	.�@�*�jɘٿl�t0���@"բ�j�3@��/�!?P'	.�@wdS�ٿ!��4��@����3@���ѐ!?s51��K�@wdS�ٿ!��4��@����3@���ѐ!?s51��K�@wdS�ٿ!��4��@����3@���ѐ!?s51��K�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@�l���ٿ����)�@9�A2�3@L����!?�6~XN�@��qSW�ٿ�M@q���@��dM�3@7��2��!?0�{���@��qSW�ٿ�M@q���@��dM�3@7��2��!?0�{���@��qSW�ٿ�M@q���@��dM�3@7��2��!?0�{���@��qSW�ٿ�M@q���@��dM�3@7��2��!?0�{���@��qSW�ٿ�M@q���@��dM�3@7��2��!?0�{���@���~åٿ��|}�x�@������3@�eа�!?x�!�
��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@ ��EK�ٿ�^���@��&�-�3@���$��!?5�X^n��@����x�ٿ��:�8�@�O�l��3@�yTaܐ!?Wl	u��@����x�ٿ��:�8�@�O�l��3@�yTaܐ!?Wl	u��@����x�ٿ��:�8�@�O�l��3@�yTaܐ!?Wl	u��@�r'"%�ٿ�+�)J�@x��=�3@_�6+��!?Sa�\��@�����ٿ-���S��@��xY	�3@�Ч���!?t�.�.(�@�����ٿ-���S��@��xY	�3@�Ч���!?t�.�.(�@�����ٿ-���S��@��xY	�3@�Ч���!?t�.�.(�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@A�Q(��ٿ��"�]S�@�7&��3@��>�ǐ!?x'4#�@D5F.
�ٿOa(� �@����3@�?G�Y�!?�e���@D5F.
�ٿOa(� �@����3@�?G�Y�!?�e���@��$�ٿK
�2���@��y��3@��^�q�!?n	�&_f�@��$�ٿK
�2���@��y��3@��^�q�!?n	�&_f�@�ER�q�ٿ{�͊6��@��Y{�3@�c�!?,����y�@�ER�q�ٿ{�͊6��@��Y{�3@�c�!?,����y�@��i~ӫٿ�*ƌ�U�@���}�3@���~Ð!?\(H��q�@��i~ӫٿ�*ƌ�U�@���}�3@���~Ð!?\(H��q�@��i~ӫٿ�*ƌ�U�@���}�3@���~Ð!?\(H��q�@��i~ӫٿ�*ƌ�U�@���}�3@���~Ð!?\(H��q�@��_�͟ٿ�E�@7"�@����3@�54�!?�6E��H�@��_�͟ٿ�E�@7"�@����3@�54�!?�6E��H�@��_�͟ٿ�E�@7"�@����3@�54�!?�6E��H�@���h�ٿCԏJ�b�@g����3@i�Ot�!?�۲����@���h�ٿCԏJ�b�@g����3@i�Ot�!?�۲����@���h�ٿCԏJ�b�@g����3@i�Ot�!?�۲����@���h�ٿCԏJ�b�@g����3@i�Ot�!?�۲����@�0��ġٿ8%2Wqy�@������3@xK����!?�L"�6�@�0��ġٿ8%2Wqy�@������3@xK����!?�L"�6�@�0��ġٿ8%2Wqy�@������3@xK����!?�L"�6�@�0��ġٿ8%2Wqy�@������3@xK����!?�L"�6�@��f�ٿ��A�F��@z?SN�3@�|����!?�8F�V$�@3W�N��ٿu��!̜�@�����3@�"`�!?a,��)�@3W�N��ٿu��!̜�@�����3@�"`�!?a,��)�@3W�N��ٿu��!̜�@�����3@�"`�!?a,��)�@3W�N��ٿu��!̜�@�����3@�"`�!?a,��)�@^��o.�ٿ������@u����3@8P�ސ!?�s&���@^��o.�ٿ������@u����3@8P�ސ!?�s&���@d�j>�ٿ�?��;)�@���G�3@j,�[��!?��?-��@Y�4%��ٿ�}��\��@`�s���3@z�4OҐ!?�+�|�@Ѹ�E�ٿ���h�@ ��i�3@X���!?��+Ř4�@��f���ٿ����"W�@ ��3@�y�ݒ�!?���
�@��f���ٿ����"W�@ ��3@�y�ݒ�!?���
�@��f���ٿ����"W�@ ��3@�y�ݒ�!?���
�@�X#�!�ٿ(�,�k�@��S3�3@#Y�D��!?)G(���@�6�/�ٿT�%ӯ��@ˉ���3@,��
�!?��0���@�6�/�ٿT�%ӯ��@ˉ���3@,��
�!?��0���@�6�/�ٿT�%ӯ��@ˉ���3@,��
�!?��0���@�6�/�ٿT�%ӯ��@ˉ���3@,��
�!?��0���@�6�/�ٿT�%ӯ��@ˉ���3@,��
�!?��0���@�J�E�ٿ��:�z��@��9E�3@����!?��^I�@�J�E�ٿ��:�z��@��9E�3@����!?��^I�@�J�E�ٿ��:�z��@��9E�3@����!?��^I�@�J�E�ٿ��:�z��@��9E�3@����!?��^I�@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@���)��ٿ1�UQ���@�ߪf�3@�a�!?���H��@�����ٿ`�o�@�}� 4@R�А!?���F^�@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@�X'I�ٿRɵ�%��@Tv�c!�3@T"�'�!?Y�u��@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@����Ϣٿ�$�����@�*^�`�3@,�\�!?�;_4���@��2��ٿ���Ɍa�@P��1�3@�$O#��!?�-8+���@��2��ٿ���Ɍa�@P��1�3@�$O#��!?�-8+���@��2��ٿ���Ɍa�@P��1�3@�$O#��!?�-8+���@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@��t�*�ٿ �>�KJ�@X,�rM�3@�/!]��!?�1�;H�@Rԓ�ŝٿ�Q�Z�
�@���!�3@䜗��!?�{?����@Rԓ�ŝٿ�Q�Z�
�@���!�3@䜗��!?�{?����@Rԓ�ŝٿ�Q�Z�
�@���!�3@䜗��!?�{?����@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@8����ٿ�э?	��@�v�3@ʳ��!?.j6Ϯ��@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@�cY�ٿ9�ZB��@�12#�3@\7�(֐!?j[�;}�@y�Jy�ٿ��5�uw�@[i(���3@X�̐!?�f�p0�@y�Jy�ٿ��5�uw�@[i(���3@X�̐!?�f�p0�@}\6�ٿ�&�GJ�@���:s�3@4��ސ!?6�>�jm�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@��:
�ٿg�4�U��@��ˡ�3@}B�W�!?�̒��v�@�I�|��ٿ��;!Z�@/Y7t3�3@��Cq��!?:X�gΓ�@ t���ٿ�Je�>��@���3@-�^�!?������@:ҜQi�ٿ_@�*��@?Yy���3@�����!?r�����@:ҜQi�ٿ_@�*��@?Yy���3@�����!?r�����@:ҜQi�ٿ_@�*��@?Yy���3@�����!?r�����@:ҜQi�ٿ_@�*��@?Yy���3@�����!?r�����@`�
��ٿ��6X�@/C�5��3@���!?���6��@`�
��ٿ��6X�@/C�5��3@���!?���6��@�����ٿ(.C�&�@p�����3@3����!?̥uO���@�����ٿ(.C�&�@p�����3@3����!?̥uO���@�����ٿ(.C�&�@p�����3@3����!?̥uO���@�����ٿ(.C�&�@p�����3@3����!?̥uO���@�����ٿ(.C�&�@p�����3@3����!?̥uO���@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@4)�_��ٿ����~�@.B�[�3@�����!?��K$��@�v��@�ٿ��R�@���y9�3@�ŗJ�!?��4��@���8O�ٿp�y��@X8d �4@�����!?�½vX��@����Ֆٿ�>�n��@�� �u�3@VKf�N�!?+�&���@����Ֆٿ�>�n��@�� �u�3@VKf�N�!?+�&���@����Ֆٿ�>�n��@�� �u�3@VKf�N�!?+�&���@����Ֆٿ�>�n��@�� �u�3@VKf�N�!?+�&���@�SJ�̑ٿ�45N�@�����3@|���!?��z�4�@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@5a�4}�ٿ�xsx�h�@wR��3@�G��!?�	1y���@��H�a�ٿh�E{RR�@�so�R�3@t�N�!?5�/���@��H�a�ٿh�E{RR�@�so�R�3@t�N�!?5�/���@��H�a�ٿh�E{RR�@�so�R�3@t�N�!?5�/���@��H�a�ٿh�E{RR�@�so�R�3@t�N�!?5�/���@�2,�h�ٿ�f�"^��@BL����3@�H}sw�!?����{�@�2,�h�ٿ�f�"^��@BL����3@�H}sw�!?����{�@�2,�h�ٿ�f�"^��@BL����3@�H}sw�!?����{�@O����ٿ�!�1��@�gZ��3@X���!?6�G�O�@O����ٿ�!�1��@�gZ��3@X���!?6�G�O�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@����=�ٿ��j޳�@�YP��3@��4�א!?�=IY.�@�v�{�ٿ`+%�$^�@F~�1��3@rH#ʐ!?T��8���@:/�ٿ7.�Z>�@b) ��3@̞�V!�!?x���Z��@:/�ٿ7.�Z>�@b) ��3@̞�V!�!?x���Z��@o�D��ٿ���ے��@T�^d�3@�����!?��.-�v�@����ٿlEQ�B�@E�Pf��3@WV9�`�!?-c����@����ٿlEQ�B�@E�Pf��3@WV9�`�!?-c����@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@Uc=���ٿ��T�1�@"aP��3@\���!?WC�h	�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@��p��ٿ'.YCC�@<����3@*
2�!?�c�++�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@�O�ٿX&�� �@h�m�3@j¢t��!?���2w�@���ٿ诵�'�@�U�F1�3@3p��Ð!?x8L��G�@���ٿ诵�'�@�U�F1�3@3p��Ð!?x8L��G�@���ٿ诵�'�@�U�F1�3@3p��Ð!?x8L��G�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@��ўٿˠhS]�@iTk��3@�	K��!?���r�@�r��ٿ�g�y�@���Ʀ�3@{ oo��!?sO�$sn�@�r��ٿ�g�y�@���Ʀ�3@{ oo��!?sO�$sn�@�r��ٿ�g�y�@���Ʀ�3@{ oo��!?sO�$sn�@�r��ٿ�g�y�@���Ʀ�3@{ oo��!?sO�$sn�@u����ٿPz�$�@�:��n�3@�[ihѐ!?N�{MUt�@������ٿO��ps��@�x�̏�3@5wMpߐ!?��[4��@������ٿO��ps��@�x�̏�3@5wMpߐ!?��[4��@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@���kܥٿ㫨+��@�0��3@�����!?�Qc���@8�3S��ٿ�t�Y��@ux��3@5��䀐!?
k�����@8�3S��ٿ�t�Y��@ux��3@5��䀐!?
k�����@8�3S��ٿ�t�Y��@ux��3@5��䀐!?
k�����@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@���#�ٿ��U���@
�
��3@c��M��!?=t�n!�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@~f���ٿ�A��	�@�{��3@6ige�!?����^�@��;l8�ٿ.�'��@>{"��3@�Y\�p�!?�3Vq���@��;l8�ٿ.�'��@>{"��3@�Y\�p�!?�3Vq���@<�_(��ٿ<��g��@�o|ɻ�3@��BN��!?�E��=�@<�_(��ٿ<��g��@�o|ɻ�3@��BN��!?�E��=�@<�_(��ٿ<��g��@�o|ɻ�3@��BN��!?�E��=�@<�_(��ٿ<��g��@�o|ɻ�3@��BN��!?�E��=�@<�_(��ٿ<��g��@�o|ɻ�3@��BN��!?�E��=�@�A�E�ٿ2�|���@�װk��3@�H�R�!?���k4��@�A�E�ٿ2�|���@�װk��3@�H�R�!?���k4��@41��Кٿ��)56��@(:��7�3@�d��!?y�M�@B6̶v�ٿ�s{���@!'���3@�����!?�ۡ�v�@��8~�ٿ�������@�5�3�3@I@���!?�:�����@��8~�ٿ�������@�5�3�3@I@���!?�:�����@��8~�ٿ�������@�5�3�3@I@���!?�:�����@��8~�ٿ�������@�5�3�3@I@���!?�:�����@��8~�ٿ�������@�5�3�3@I@���!?�:�����@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@Wn���ٿ���-c�@�����3@����!?5��i8�@zXY�ٿ}��]�@_�4'��3@��+�!?}�SB�@�p-��ٿ�d�Q���@(ݒ�p�3@A�\�3�!?𥆪U�@�p-��ٿ�d�Q���@(ݒ�p�3@A�\�3�!?𥆪U�@�+�ǣٿ:o����@��
k�3@6���	�!?�\c����@�+�ǣٿ:o����@��
k�3@6���	�!?�\c����@�+�ǣٿ:o����@��
k�3@6���	�!?�\c����@Nݏ��ٿ?>r���@����3@Y��!?1��2M�@Nݏ��ٿ?>r���@����3@Y��!?1��2M�@Nݏ��ٿ?>r���@����3@Y��!?1��2M�@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@�!�3"�ٿ�0k
���@$
�n(�3@�׉��!?]S����@>��@��ٿ����z�@y����3@V���p�!?{Ǜx�@>��@��ٿ����z�@y����3@V���p�!?{Ǜx�@>��@��ٿ����z�@y����3@V���p�!?{Ǜx�@�[���ٿ(ۅ���@�(����3@^ڗKʐ!?pk�U$�@�[���ٿ(ۅ���@�(����3@^ڗKʐ!?pk�U$�@�[���ٿ(ۅ���@�(����3@^ڗKʐ!?pk�U$�@�[���ٿ(ۅ���@�(����3@^ڗKʐ!?pk�U$�@�[���ٿ(ۅ���@�(����3@^ڗKʐ!?pk�U$�@(I+��ٿ'���@��m��3@�M9ݐ!?��d�s��@K�����ٿ������@��	ݶ�3@K-c3m�!?}���^Y�@��꼘ٿ����#�@e>M��3@��ظ�!?|�m���@��꼘ٿ����#�@e>M��3@��ظ�!?|�m���@�EM��ٿ#��f�@ �\��3@�9RÐ!?��ݮ��@�EM��ٿ#��f�@ �\��3@�9RÐ!?��ݮ��@�EM��ٿ#��f�@ �\��3@�9RÐ!?��ݮ��@�EM��ٿ#��f�@ �\��3@�9RÐ!?��ݮ��@�EM��ٿ#��f�@ �\��3@�9RÐ!?��ݮ��@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@� 36�ٿ�}i���@�!}&��3@�/x��!?G<dP �@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@|t�ݠ�ٿ'l`se��@N���3@��-�!?��̒�#�@Μx�]�ٿ���7��@a���m�3@�<��k�!?z?�v��@Μx�]�ٿ���7��@a���m�3@�<��k�!?z?�v��@8����ٿɾG��k�@z�� H�3@�����!?��m{3d�@���J��ٿ�ǒe��@{�n��3@��s�z�!?�{��e�@���J��ٿ�ǒe��@{�n��3@��s�z�!?�{��e�@���J��ٿ�ǒe��@{�n��3@��s�z�!?�{��e�@���J��ٿ�ǒe��@{�n��3@��s�z�!?�{��e�@,��\ݨٿ�KK���@�n&�3@�s��`�!?:e�n<�@,��\ݨٿ�KK���@�n&�3@�s��`�!?:e�n<�@,��\ݨٿ�KK���@�n&�3@�s��`�!?:e�n<�@,��\ݨٿ�KK���@�n&�3@�s��`�!?:e�n<�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@���Ʃ�ٿ��e5c�@Й,���3@�y3�!?%z\Uo�@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@&��ly�ٿ�㋿(��@�)e���3@�ى��!?Z�5_���@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@��@��ٿBO��Њ�@���S|�3@E�L�ѐ!?~͵�;�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@�I��ٿ�VI���@�����3@oEcЪ�!?vUݞ<�@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@%�.�ٿ��32 ��@���b�3@ ��驐!?c�����@�r�̤ٿ��`P�p�@Tئ��3@�ڕNw�!?w!�s"L�@�r�̤ٿ��`P�p�@Tئ��3@�ڕNw�!?w!�s"L�@�r�̤ٿ��`P�p�@Tئ��3@�ڕNw�!?w!�s"L�@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@����ٿ��ݏS�@�6��3@��*���!?�!9Z��@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�|@g�ٿ6򮷂g�@�qD���3@��~`ڐ!?"�#mu�@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@�Q�Q�ٿ�Q~�T��@:t����3@+s��!?F
u�]��@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@u�N?�ٿ�����@&�����3@{���!?�y�<>x�@��#Ţ�ٿ��`A�@�~�fg�3@b�D��!?kN����@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@�7���ٿh޹YG��@Ƶ����3@�E9��!?P^?V�@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@]F)Yןٿ���_$/�@`��\/�3@�{ﱐ!?-�^���@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�_�Q��ٿ�ZGD�@�����3@l�$���!?�s�!JK�@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@�)�,�ٿ�43J=d�@���!��3@Bg/}��!?�4:�.��@��0�}�ٿ�XV�w��@��I���3@A�$l�!?%�Gw��@��0�}�ٿ�XV�w��@��I���3@A�$l�!?%�Gw��@��0�}�ٿ�XV�w��@��I���3@A�$l�!?%�Gw��@��0�}�ٿ�XV�w��@��I���3@A�$l�!?%�Gw��@�7���ٿB�K��@�V��3@K��>��!?�~ ��#�@�7���ٿB�K��@�V��3@K��>��!?�~ ��#�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@�"|�ٿg���x��@�>�7�3@�7w�Ր!?x-�{2�@B2��ٿ�U����@�]���3@��*�!?�<��_�@B2��ٿ�U����@�]���3@��*�!?�<��_�@B2��ٿ�U����@�]���3@��*�!?�<��_�@B2��ٿ�U����@�]���3@��*�!?�<��_�@B2��ٿ�U����@�]���3@��*�!?�<��_�@B2��ٿ�U����@�]���3@��*�!?�<��_�@� �<�ٿ�^4��D�@=J�ϱ�3@�d|	֐!?���C�@� �<�ٿ�^4��D�@=J�ϱ�3@�d|	֐!?���C�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@S�U4�ٿ��W�G��@ũ�[_�3@%j��̐!?c*[V�@��I)�ٿ�cr����@�k^8m�3@5�ӏk�!?�w���@��I)�ٿ�cr����@�k^8m�3@5�ӏk�!?�w���@��I)�ٿ�cr����@�k^8m�3@5�ӏk�!?�w���@��I)�ٿ�cr����@�k^8m�3@5�ӏk�!?�w���@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@���V�ٿ� PZU��@�G&
��3@�W�H}�!?���#�@b�q7̣ٿ�꜠��@���-��3@���S��!?��^�+c�@b�q7̣ٿ�꜠��@���-��3@���S��!?��^�+c�@b�q7̣ٿ�꜠��@���-��3@���S��!?��^�+c�@b�q7̣ٿ�꜠��@���-��3@���S��!?��^�+c�@b�q7̣ٿ�꜠��@���-��3@���S��!?��^�+c�@�$џ��ٿ�c����@Xn{P��3@���!?,|��w�@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@<m=NǢٿ ����@L��<�3@�.G���!?af����@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@�o�j�ٿI��҂�@� ����3@l�t��!?N�y%��@����x�ٿY��+�*�@9o��3@b.���!?� ����@����x�ٿY��+�*�@9o��3@b.���!?� ����@�׎��ٿK�[%��@}��A�3@�gg&��!?�/��U�@�׎��ٿK�[%��@}��A�3@�gg&��!?�/��U�@�׎��ٿK�[%��@}��A�3@�gg&��!?�/��U�@�׎��ٿK�[%��@}��A�3@�gg&��!?�/��U�@�d���ٿ�䷡4�@�Kv��3@�թ1��!?��2��@9VA�N�ٿ��9+��@�&5�	�3@�?�[s�!?9�ƊX�@��nN�ٿ�m����@�
4L��3@�� ��!?´��*5�@��nN�ٿ�m����@�
4L��3@�� ��!?´��*5�@��nN�ٿ�m����@�
4L��3@�� ��!?´��*5�@��nN�ٿ�m����@�
4L��3@�� ��!?´��*5�@��nN�ٿ�m����@�
4L��3@�� ��!?´��*5�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@����m�ٿ%e�f�@�i��3@˕���!?,~�b	�@��)X��ٿՠ�ő�@�1Pp!�3@a�<c��!?�#b0���@*J]��ٿJ ����@[bZ|9�3@Y��hϐ!?Coq�[K�@�y�.�ٿcV!ZZ�@���@��3@��� �!?��+�@�!��ٿ9��'��@!ߛZd�3@xD
�!?����<�@�!��ٿ9��'��@!ߛZd�3@xD
�!?����<�@�!��ٿ9��'��@!ߛZd�3@xD
�!?����<�@�!��ٿ9��'��@!ߛZd�3@xD
�!?����<�@�!��ٿ9��'��@!ߛZd�3@xD
�!?����<�@T�����ٿ�u)��@�Y�P��3@�@��!?[�*�]�@T�����ٿ�u)��@�Y�P��3@�@��!?[�*�]�@T�����ٿ�u)��@�Y�P��3@�@��!?[�*�]�@T�����ٿ�u)��@�Y�P��3@�@��!?[�*�]�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@�h���ٿ����4|�@^���3@�?Z-��!?S�{`x�@ҧ84��ٿ`/�=O�@��y�*�3@�v���!?Sp1�"�@ҧ84��ٿ`/�=O�@��y�*�3@�v���!?Sp1�"�@ҧ84��ٿ`/�=O�@��y�*�3@�v���!?Sp1�"�@ҧ84��ٿ`/�=O�@��y�*�3@�v���!?Sp1�"�@ҧ84��ٿ`/�=O�@��y�*�3@�v���!?Sp1�"�@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@xbڭH�ٿS�h����@Ң�J��3@2I��!?��g��@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@�Y3v�ٿ����(��@K�?Y�3@3X��!?�t�)�@T��ܣٿ�=@p
��@�DZ��3@:4_Ő!?�x�^���@]=����ٿM�T�P2�@9�Õ��3@�2���!?v�DK���@]=����ٿM�T�P2�@9�Õ��3@�2���!?v�DK���@�Q5eF�ٿ=�����@��"G�3@e���ɐ!?/�����@�Q5eF�ٿ=�����@��"G�3@e���ɐ!?/�����@�Q5eF�ٿ=�����@��"G�3@e���ɐ!?/�����@�lΡ2�ٿ��<��@QV&=�3@�D�χ�!?~[%��q�@�lΡ2�ٿ��<��@QV&=�3@�D�χ�!?~[%��q�@�lΡ2�ٿ��<��@QV&=�3@�D�χ�!?~[%��q�@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@�J�K��ٿ��(f(��@�*^$��3@{5(p��!?.XU���@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@H���ٿqW]*+�@WĈ�|�3@�{ϐ!?GW�pIG�@|r���ٿHͷ�&�@b���+�3@��}3o�!?��_��+�@|r���ٿHͷ�&�@b���+�3@��}3o�!?��_��+�@|r���ٿHͷ�&�@b���+�3@��}3o�!?��_��+�@|r���ٿHͷ�&�@b���+�3@��}3o�!?��_��+�@|r���ٿHͷ�&�@b���+�3@��}3o�!?��_��+�@v�]0J�ٿ]&���@.�-f�3@�L`ؘ�!?S�� �\�@����ŝٿB�r��1�@���3@��)��!?*(�I��@����ŝٿB�r��1�@���3@��)��!?*(�I��@����ŝٿB�r��1�@���3@��)��!?*(�I��@W����ٿ�h�#"��@�-o��3@�>�Yΐ!?���A��@W����ٿ�h�#"��@�-o��3@�>�Yΐ!?���A��@W����ٿ�h�#"��@�-o��3@�>�Yΐ!?���A��@�>�	�ٿ�a��fE�@/t����3@��9#А!?�ϯ��!�@�>�	�ٿ�a��fE�@/t����3@��9#А!?�ϯ��!�@�>�	�ٿ�a��fE�@/t����3@��9#А!?�ϯ��!�@��Q0B�ٿuc�v�5�@S�NT�3@؝q���!?�P�`�@c�Q�j�ٿ�h�.��@fK��3@X�2u�!?��Y�R�@��gz��ٿU�)��@˿����3@�D
WŐ!?x��/�&�@��gz��ٿU�)��@˿����3@�D
WŐ!?x��/�&�@��gz��ٿU�)��@˿����3@�D
WŐ!?x��/�&�@��gz��ٿU�)��@˿����3@�D
WŐ!?x��/�&�@��gz��ٿU�)��@˿����3@�D
WŐ!?x��/�&�@�vX���ٿ��>�I�@(�mE�3@`,!��!?�U^����@�vX���ٿ��>�I�@(�mE�3@`,!��!?�U^����@�C�ѥٿD�����@�0�y�3@'F�ߐ!?s��r��@�V��>�ٿ�Z�ˆ��@2N��3@�qM���!?z0�G���@�V��>�ٿ�Z�ˆ��@2N��3@�qM���!?z0�G���@�V��>�ٿ�Z�ˆ��@2N��3@�qM���!?z0�G���@�V��>�ٿ�Z�ˆ��@2N��3@�qM���!?z0�G���@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@�p���ٿe���[��@�:�{n�3@�d�!?]z�:��@��,���ٿ?X�=�/�@�^`�3@��˜�!??:W�R7�@��,���ٿ?X�=�/�@�^`�3@��˜�!??:W�R7�@��,���ٿ?X�=�/�@�^`�3@��˜�!??:W�R7�@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@2+#o��ٿ9�:+s&�@�[Q�3@���vِ!?����@ڕ2&�ٿ�����(�@3"��D�3@H?gÐ!?ٻr�i3�@�|�ћٿxĈ���@�\`���3@�H��!?�~O�}�@�|�ћٿxĈ���@�\`���3@�H��!?�~O�}�@�|�ћٿxĈ���@�\`���3@�H��!?�~O�}�@��$O��ٿ��Ӏ��@t��N�3@����!?�Y�F���@��$O��ٿ��Ӏ��@t��N�3@����!?�Y�F���@��$O��ٿ��Ӏ��@t��N�3@����!?�Y�F���@2��P��ٿ\���G��@���3@?,��Ր!?�׹��{�@2��P��ٿ\���G��@���3@?,��Ր!?�׹��{�@2��P��ٿ\���G��@���3@?,��Ր!?�׹��{�@�譆�ٿs�����@��Ą��3@�z��ː!?�Oj0���@)�(�ٿ�e�@*��a>�3@�O�xې!?)q��@��;:�ٿwt
 fV�@�x�#�3@D[����!?i�Q��b�@��;:�ٿwt
 fV�@�x�#�3@D[����!?i�Q��b�@��;:�ٿwt
 fV�@�x�#�3@D[����!?i�Q��b�@ P �ٿ�����@S����3@�ᨠ�!?���9��@ P �ٿ�����@S����3@�ᨠ�!?���9��@ P �ٿ�����@S����3@�ᨠ�!?���9��@��p�ٿI���T�@���P�3@pZ%4ܐ!?m��"��@��p�ٿI���T�@���P�3@pZ%4ܐ!?m��"��@�w�2ŗٿ����a��@��!=�3@YkD��!?��h�@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@�����ٿ�昞��@����3@�����!?�+Q����@9�5�s�ٿ�S����@��p6�3@��򲄐!?�l��,��@ROZ�Şٿ�v��zE�@V�����3@�n�4��!?7o_�x�@ROZ�Şٿ�v��zE�@V�����3@�n�4��!?7o_�x�@ROZ�Şٿ�v��zE�@V�����3@�n�4��!?7o_�x�@iq�6�ٿN�a���@�ʞ��3@����!?��7��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@j;R�ɘٿKLb9��@�����3@�g���!?YPfo��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@�N@ �ٿ������@����3@6J�q��!?�ͬ��@{��ٿ7�K7,��@s$o�3@Y�d�!?m�7����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@����ٿ�A�aa	�@U��3@�N����!?M�����@���̟ٿ�����\�@Hz�l��3@�]Y��!?[���
b�@����ٿDo�8��@�3g���3@ �8�!?ʱ�5��@����ٿDo�8��@�3g���3@ �8�!?ʱ�5��@����ٿDo�8��@�3g���3@ �8�!?ʱ�5��@����ٿDo�8��@�3g���3@ �8�!?ʱ�5��@V���ٿQDƉRF�@��:��3@B���!?�|��i��@V���ٿQDƉRF�@��:��3@B���!?�|��i��@V���ٿQDƉRF�@��:��3@B���!?�|��i��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@k܄aW�ٿ*�v\��@g�n�y�3@�S�!?��2zB��@�����ٿ]A����@�z�*�3@2̡��!?�E�ño�@��
ޠٿ�HW9��@����(�3@)ֳ���!?�/š@g�@��"ޣٿ:��L�}�@����3@���̐!?���]&-�@��"ޣٿ:��L�}�@����3@���̐!?���]&-�@��"ޣٿ:��L�}�@����3@���̐!?���]&-�@��"ޣٿ:��L�}�@����3@���̐!?���]&-�@��3���ٿr�����@�Y���3@딛m!?S�7�@��3���ٿr�����@�Y���3@딛m!?S�7�@��3���ٿr�����@�Y���3@딛m!?S�7�@��3���ٿr�����@�Y���3@딛m!?S�7�@��3���ٿr�����@�Y���3@딛m!?S�7�@��3���ٿr�����@�Y���3@딛m!?S�7�@��}̡ٿ����?��@.�~���3@�W�'�!?����@�@��}̡ٿ����?��@.�~���3@�W�'�!?����@�@��}̡ٿ����?��@.�~���3@�W�'�!?����@�@�x��ʣٿ�AFC�"�@�!��3@:�CJӐ!?>}O��@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@R�oY�ٿE)x���@P�t��3@f9��!?1���d0�@v?g'�ٿU�!�Q��@K��f�3@��L�!?��A)O�@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@�ٸ�F�ٿ�mpOL�@*^N���3@�����!?�"���@,
^� �ٿ�4 ���@�y�pW�3@y�ސ!?�?�e���@,
^� �ٿ�4 ���@�y�pW�3@y�ސ!?�?�e���@,
^� �ٿ�4 ���@�y�pW�3@y�ސ!?�?�e���@,
^� �ٿ�4 ���@�y�pW�3@y�ސ!?�?�e���@,
^� �ٿ�4 ���@�y�pW�3@y�ސ!?�?�e���@U,���ٿ,f@b��@���9�3@	�i��!?�֪\#s�@U,���ٿ,f@b��@���9�3@	�i��!?�֪\#s�@U,���ٿ,f@b��@���9�3@	�i��!?�֪\#s�@ԛ2%�ٿ(��r���@�F|w-�3@C�w'Ð!?R@W_�@ԛ2%�ٿ(��r���@�F|w-�3@C�w'Ð!?R@W_�@+
<A�ٿZ�VΈ�@քp��3@H�:#��!?��Ff��@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@�?�(��ٿlP�jy��@=�(-��3@%��ݶ�!?�$eKt�@Y9��n�ٿ�Z|�]�@5[̈]�3@s뼞�!?�N<���@Y9��n�ٿ�Z|�]�@5[̈]�3@s뼞�!?�N<���@�L���ٿq%����@�څ�3@���J��!?�z�.v��@�L���ٿq%����@�څ�3@���J��!?�z�.v��@���C�ٿB:��1��@�&���3@���� �!?\�߸t!�@���C�ٿB:��1��@�&���3@���� �!?\�߸t!�@���C�ٿB:��1��@�&���3@���� �!?\�߸t!�@���C�ٿB:��1��@�&���3@���� �!?\�߸t!�@ֵ@��ٿq
�
u�@^����3@>�&/��!?�0�x�@ֵ@��ٿq
�
u�@^����3@>�&/��!?�0�x�@ֵ@��ٿq
�
u�@^����3@>�&/��!?�0�x�@ֵ@��ٿq
�
u�@^����3@>�&/��!?�0�x�@�Ӟ���ٿ��p��@��1M��3@w��А!?E��T4�@�Ӟ���ٿ��p��@��1M��3@w��А!?E��T4�@�^q��ٿ*Tqx�@�T�-X�3@'���7�!?e?g�B��@f
h���ٿޯ���@��T�3@�*�3Z�!?g�2k��@f
h���ٿޯ���@��T�3@�*�3Z�!?g�2k��@f
h���ٿޯ���@��T�3@�*�3Z�!?g�2k��@f
h���ٿޯ���@��T�3@�*�3Z�!?g�2k��@���:�ٿ��\�@EH��z�3@�M@S�!?�����@���:�ٿ��\�@EH��z�3@�M@S�!?�����@���:�ٿ��\�@EH��z�3@�M@S�!?�����@��	��ٿ9��|�@�YK7��3@��r�2�!?����f��@��	��ٿ9��|�@�YK7��3@��r�2�!?����f��@��	��ٿ9��|�@�YK7��3@��r�2�!?����f��@��	��ٿ9��|�@�YK7��3@��r�2�!?����f��@�4���ٿ�mk2:��@��{;��3@�1}��!?��u<		�@�4���ٿ�mk2:��@��{;��3@�1}��!?��u<		�@G�I(f�ٿ���	�@��!�3@�s�g�!?1)�/�@�8�p�ٿ$�#�"��@FSeI��3@�ܱ휐!?J_�Ј2�@�#H��ٿ�����@�|��3@/�d��!?��ge\��@�da1�ٿ�ɳ���@��B�3@׵���!??3��Y��@�da1�ٿ�ɳ���@��B�3@׵���!??3��Y��@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@D��y֢ٿ�ӭ�{J�@�m"��3@���Kې!?��z��p�@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@��5.�ٿ,��b|~�@z� m��3@�.��A�!?'��[��@ʫ�݊�ٿ�b�I���@e��>�3@��:�ѐ!?O�'�@ʫ�݊�ٿ�b�I���@e��>�3@��:�ѐ!?O�'�@ʫ�݊�ٿ�b�I���@e��>�3@��:�ѐ!?O�'�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@?sC�b�ٿ�����@�wd��3@����ِ!?�
8�ԇ�@��s�ٿ���v�@�m#S��3@�`༠�!?k:��q�@��s�ٿ���v�@�m#S��3@�`༠�!?k:��q�@��s�ٿ���v�@�m#S��3@�`༠�!?k:��q�@��x!��ٿ,Y$ρ*�@�V'�=�3@sZ��ʐ!?Ǜ�����@��x!��ٿ,Y$ρ*�@�V'�=�3@sZ��ʐ!?Ǜ�����@��x!��ٿ,Y$ρ*�@�V'�=�3@sZ��ʐ!?Ǜ�����@��x!��ٿ,Y$ρ*�@�V'�=�3@sZ��ʐ!?Ǜ�����@��x!��ٿ,Y$ρ*�@�V'�=�3@sZ��ʐ!?Ǜ�����@��%�U�ٿR����C�@;B?�3@��C!?ҫ����@�>fh+�ٿC|�aE9�@(�� �3@��j��!?�����U�@�>fh+�ٿC|�aE9�@(�� �3@��j��!?�����U�@�_���ٿ������@�!�i��3@E�O� �!?Q��x�t�@�_���ٿ������@�!�i��3@E�O� �!?Q��x�t�@�_���ٿ������@�!�i��3@E�O� �!?Q��x�t�@�_���ٿ������@�!�i��3@E�O� �!?Q��x�t�@�۲��ٿvq��%�@|�:��3@�m&�!?g j|���@�۲��ٿvq��%�@|�:��3@�m&�!?g j|���@ь�ݢٿ?b�Z+�@�S�H��3@�=ٔ��!?�1	����@ь�ݢٿ?b�Z+�@�S�H��3@�=ٔ��!?�1	����@ь�ݢٿ?b�Z+�@�S�H��3@�=ٔ��!?�1	����@ь�ݢٿ?b�Z+�@�S�H��3@�=ٔ��!?�1	����@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@3Q��ٿ���D�n�@hy�� �3@��l_	�!?�qV�ԩ�@��iX�ٿM)|��@�x'm��3@�n�dː!?�U����@��iX�ٿM)|��@�x'm��3@�n�dː!?�U����@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@N�)�ʛٿq$�Q>�@kD��3@Xo���!?���}�@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@3��'�ٿ�đx�U�@�ǀ��3@7�ǳ�!?�f�jy��@S�zɝٿv�c
=�@X �F�3@��Zʐ!?�H&q��@%j�2��ٿ'��$��@J��s��3@x�Wj��!?�|��7+�@%j�2��ٿ'��$��@J��s��3@x�Wj��!?�|��7+�@%j�2��ٿ'��$��@J��s��3@x�Wj��!?�|��7+�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�J�>�ٿp�
�V�@����3@���f��!?���g�@�@�:�Ǜٿyb�� ��@�E�v��3@�ѐ!?~�_�e]�@�:�Ǜٿyb�� ��@�E�v��3@�ѐ!?~�_�e]�@�:�Ǜٿyb�� ��@�E�v��3@�ѐ!?~�_�e]�@�:�Ǜٿyb�� ��@�E�v��3@�ѐ!?~�_�e]�@�:�Ǜٿyb�� ��@�E�v��3@�ѐ!?~�_�e]�@�Z���ٿ���阄�@�تWP�3@2h[@�!?	�<�)��@ ��v-�ٿ���4��@��XI�3@;b��!?�l0���@���şٿ��Ё��@�E�`h�3@$�>^Ր!?\"�%*��@���şٿ��Ё��@�E�`h�3@$�>^Ր!?\"�%*��@���şٿ��Ё��@�E�`h�3@$�>^Ր!?\"�%*��@���şٿ��Ё��@�E�`h�3@$�>^Ր!?\"�%*��@�vz۟ٿ�[��x�@vM-
�3@�Ja��!?%7�%��@�vz۟ٿ�[��x�@vM-
�3@�Ja��!?%7�%��@�vz۟ٿ�[��x�@vM-
�3@�Ja��!?%7�%��@���>v�ٿ!�7����@��}X��3@��f �!?��j��@���>v�ٿ!�7����@��}X��3@��f �!?��j��@���>v�ٿ!�7����@��}X��3@��f �!?��j��@���>v�ٿ!�7����@��}X��3@��f �!?��j��@�i��ϛٿW�a�@�(_z�3@z�y��!?4o�2%�@�i��ϛٿW�a�@�(_z�3@z�y��!?4o�2%�@�i��ϛٿW�a�@�(_z�3@z�y��!?4o�2%�@�i��ϛٿW�a�@�(_z�3@z�y��!?4o�2%�@��"�G�ٿ�Z����@�A�z��3@���K��!?�=��"��@��"�G�ٿ�Z����@�A�z��3@���K��!?�=��"��@��"�G�ٿ�Z����@�A�z��3@���K��!?�=��"��@��"�G�ٿ�Z����@�A�z��3@���K��!?�=��"��@��"�G�ٿ�Z����@�A�z��3@���K��!?�=��"��@�i(�ٿ���֙�@]�u���3@B߆9��!?������@��t*�ٿ�+�Njy�@�2�(�3@zy��ѐ!?��.�K%�@�D�ʑ�ٿ�м���@Ws(��3@��Y���!?C���@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@�rՊ�ٿ^���1L�@2��!I�3@���m�!?Y)�c[��@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@����ܛٿ��|��@=� ��3@�w�b�!?.��jaA�@UW��יٿ4:c%z��@�b���3@�t�y��!?D���L�@�1�p��ٿ���L9��@U� (�3@����!?��k�
�@�1�p��ٿ���L9��@U� (�3@����!?��k�
�@��Ɖ�ٿS1$�'R�@�!b}��3@p�i��!?��,��r�@��Ɖ�ٿS1$�'R�@�!b}��3@p�i��!?��,��r�@&oe�ٿ!�g����@M��u�3@�����!?��K���@����ġٿ��75�%�@�G�rA�3@��8}�!?��#��@y��'�ٿt-�Y&��@��u��3@�;c���!?�3]S�T�@y��'�ٿt-�Y&��@��u��3@�;c���!?�3]S�T�@y��'�ٿt-�Y&��@��u��3@�;c���!?�3]S�T�@y��'�ٿt-�Y&��@��u��3@�;c���!?�3]S�T�@��1�ٿtY �0��@#�Nu�3@tUU���!?�b|���@��1�ٿtY �0��@#�Nu�3@tUU���!?�b|���@��1�ٿtY �0��@#�Nu�3@tUU���!?�b|���@��1�ٿtY �0��@#�Nu�3@tUU���!?�b|���@��1�ٿtY �0��@#�Nu�3@tUU���!?�b|���@\ �@�ٿ�S�Ь��@Dg��3�3@{@�'�!?��J�Tx�@\ �@�ٿ�S�Ь��@Dg��3�3@{@�'�!?��J�Tx�@\ �@�ٿ�S�Ь��@Dg��3�3@{@�'�!?��J�Tx�@\ �@�ٿ�S�Ь��@Dg��3�3@{@�'�!?��J�Tx�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@n�@�7�ٿ�k�q\�@�����3@���ؐ!?sH�!�,�@��W��ٿE�N$��@^Ov��3@����Ő!?�0;��@��W��ٿE�N$��@^Ov��3@����Ő!?�0;��@?"�}��ٿ��mt��@TނC�3@��Eǐ!?kt��}�@JXllÝٿ�ak����@y~��3@��C�!?��-!.�@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@����ٿM'�F��@�U��b�3@�l��!?�j�ڷ��@��PS�ٿI�hs4'�@Z"õ��3@���U�!?�kH����@��PS�ٿI�hs4'�@Z"õ��3@���U�!?�kH����@��PS�ٿI�hs4'�@Z"õ��3@���U�!?�kH����@��PS�ٿI�hs4'�@Z"õ��3@���U�!?�kH����@��PS�ٿI�hs4'�@Z"õ��3@���U�!?�kH����@��c��ٿ�M�����@.��l��3@�+%�X�!?:J�$� �@7����ٿyD=�*E�@���r�3@Cِ!? �@�8��@7����ٿyD=�*E�@���r�3@Cِ!? �@�8��@7����ٿyD=�*E�@���r�3@Cِ!? �@�8��@���@�ٿLV�,dL�@�G"5��3@�cLJߐ!?_yL���@���@�ٿLV�,dL�@�G"5��3@�cLJߐ!?_yL���@q�����ٿ<K�����@��W�
�3@�2��!?޺,@��@q�����ٿ<K�����@��W�
�3@�2��!?޺,@��@q�����ٿ<K�����@��W�
�3@�2��!?޺,@��@��sģٿ���D��@��ڬ��3@M��ߐ!?�N�NȻ�@��sģٿ���D��@��ڬ��3@M��ߐ!?�N�NȻ�@��sģٿ���D��@��ڬ��3@M��ߐ!?�N�NȻ�@��sģٿ���D��@��ڬ��3@M��ߐ!?�N�NȻ�@��sģٿ���D��@��ڬ��3@M��ߐ!?�N�NȻ�@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@�g3��ٿ�9�U~��@����3@+E�Tϐ!?��� G��@��)�ٿ������@N�;/�3@��t��!?� �����@��)�ٿ������@N�;/�3@��t��!?� �����@��)�ٿ������@N�;/�3@��t��!?� �����@��)�ٿ������@N�;/�3@��t��!?� �����@��)�ٿ������@N�;/�3@��t��!?� �����@W�h�ߠٿw�P�D�@���!a�3@�`���!?G<�UX��@W�h�ߠٿw�P�D�@���!a�3@�`���!?G<�UX��@��o�P�ٿ�6Q �R�@��\?��3@ ��ΐ!?�l�����@��o�P�ٿ�6Q �R�@��\?��3@ ��ΐ!?�l�����@��o�P�ٿ�6Q �R�@��\?��3@ ��ΐ!?�l�����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@�ܨNݥٿ+��h;�@���؋�3@g�S�Ȑ!?�9P����@i�Ļݞٿ6�tM^��@l�4���3@;T���!?�J�P}�@i�Ļݞٿ6�tM^��@l�4���3@;T���!?�J�P}�@i�Ļݞٿ6�tM^��@l�4���3@;T���!?�J�P}�@Z׌�L�ٿ�wrkl��@�LX?��3@Ҭȅ��!?R*^�-��@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@;C�a0�ٿ36���)�@�Â-��3@�:X��!?��4���@�3� b�ٿ�7z^d��@�M�
�3@�{�;А!?-�����@�3� b�ٿ�7z^d��@�M�
�3@�{�;А!?-�����@�3� b�ٿ�7z^d��@�M�
�3@�{�;А!?-�����@�3� b�ٿ�7z^d��@�M�
�3@�{�;А!?-�����@�3� b�ٿ�7z^d��@�M�
�3@�{�;А!?-�����@޸� ��ٿtɒ&��@B97�3@J����!?��ʽ�@޸� ��ٿtɒ&��@B97�3@J����!?��ʽ�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@A��bL�ٿG� �-�@U����3@�ij�!?'ı�|�@���ϡٿO��.�@"X�x�3@��7��!?�j���b�@���ϡٿO��.�@"X�x�3@��7��!?�j���b�@���ϡٿO��.�@"X�x�3@��7��!?�j���b�@�t���ٿ?����@+i�'I�3@�'%E��!?$��=ν�@�5�ٿdN_��c�@�=�Ֆ�3@�FR�ː!?~�M��3�@�5�ٿdN_��c�@�=�Ֆ�3@�FR�ː!?~�M��3�@�5�ٿdN_��c�@�=�Ֆ�3@�FR�ː!?~�M��3�@�5�ٿdN_��c�@�=�Ֆ�3@�FR�ː!?~�M��3�@�5�ٿdN_��c�@�=�Ֆ�3@�FR�ː!?~�M��3�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@bU6�Пٿ�� �3�@�=7�G�3@�Әo�!??�deG�@;>\�l�ٿ����@O�_\��3@C���!?�`2=j��@;>\�l�ٿ����@O�_\��3@C���!?�`2=j��@;>\�l�ٿ����@O�_\��3@C���!?�`2=j��@;>\�l�ٿ����@O�_\��3@C���!?�`2=j��@0mI��ٿ��3�5��@y�CiJ�3@e�Eސ!?�?���b�@0mI��ٿ��3�5��@y�CiJ�3@e�Eސ!?�?���b�@0mI��ٿ��3�5��@y�CiJ�3@e�Eސ!?�?���b�@}v	�ٿ,��6��@�����3@�����!?��Jr��@�����ٿk��s��@{C����3@���Fː!?_ D��n�@�����ٿk��s��@{C����3@���Fː!?_ D��n�@�����ٿk��s��@{C����3@���Fː!?_ D��n�@�N��ɟٿtŸ!{�@��?@�3@����֐!?�c���n�@�N��ɟٿtŸ!{�@��?@�3@����֐!?�c���n�@�N��ɟٿtŸ!{�@��?@�3@����֐!?�c���n�@�N��ɟٿtŸ!{�@��?@�3@����֐!?�c���n�@�x��E�ٿ�^�T��@�BH�c�3@�����!?�]H  ��@�x��E�ٿ�^�T��@�BH�c�3@�����!?�]H  ��@�+����ٿ�	=F��@ek���3@(F7ѐ!?Wx��H1�@�+����ٿ�	=F��@ek���3@(F7ѐ!?Wx��H1�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@��z4�ٿk>��x�@�uf��3@���}�!?A��tH�@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@Ӹ�&Şٿ�U!#1�@��3qp�3@�D�i��!?��7��@���\�ٿ�zL���@�����3@/|��ؐ!?g7���@���\�ٿ�zL���@�����3@/|��ؐ!?g7���@�)L}�ٿ���r��@�luU�3@�{�k֐!?T�v�)��@�)L}�ٿ���r��@�luU�3@�{�k֐!?T�v�)��@�)L}�ٿ���r��@�luU�3@�{�k֐!?T�v�)��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@	�ט*�ٿ����?��@V�gV��3@YJ���!?�6}_��@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@�ũ:�ٿ3��s&��@�=�a��3@N�&ɐ!?Q�Ὀ�@8w(h�ٿ���&�$�@�}v]��3@;�ȱ�!?��
���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@�T0�8�ٿ+��m�E�@2����3@�E�n��!?���n���@Ac9���ٿ�9��c�@ɡ�Y��3@AI�樐!?&]^��@Ac9���ٿ�9��c�@ɡ�Y��3@AI�樐!?&]^��@Ac9���ٿ�9��c�@ɡ�Y��3@AI�樐!?&]^��@Ac9���ٿ�9��c�@ɡ�Y��3@AI�樐!?&]^��@�{O��ٿ[˻]�@��ʱf�3@W���ߐ!?Ʉ�P>�@�{O��ٿ[˻]�@��ʱf�3@W���ߐ!?Ʉ�P>�@�{O��ٿ[˻]�@��ʱf�3@W���ߐ!?Ʉ�P>�@�{O��ٿ[˻]�@��ʱf�3@W���ߐ!?Ʉ�P>�@�t�v�ٿ���A���@b<f��3@E�Ē�!?Z���el�@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�?�b7�ٿ�у(��@g|���3@�"!?F��w���@�R�˟ٿR�>45��@b|,��3@�K냑�!?���(��@�R�˟ٿR�>45��@b|,��3@�K냑�!?���(��@�R�˟ٿR�>45��@b|,��3@�K냑�!?���(��@�R�˟ٿR�>45��@b|,��3@�K냑�!?���(��@&��$�ٿ�Ա]#�@,����3@^ڔ��!?��K�8��@&��$�ٿ�Ա]#�@,����3@^ڔ��!?��K�8��@&��$�ٿ�Ա]#�@,����3@^ڔ��!?��K�8��@��G�ҚٿsN�s��@�q�!�3@eB��!?#gt7�I�@��G�ҚٿsN�s��@�q�!�3@eB��!?#gt7�I�@��G�ҚٿsN�s��@�q�!�3@eB��!?#gt7�I�@��G�ҚٿsN�s��@�q�!�3@eB��!?#gt7�I�@��G�ҚٿsN�s��@�q�!�3@eB��!?#gt7�I�@�  �ٿi8�e���@UZ�8�3@T�j��!?��7o�@$�>�0�ٿ�Aho��@E��w�3@%���!?��y\��@*�-7�ٿ�M����@aS�~��3@p�g/�!?�W�s���@*�-7�ٿ�M����@aS�~��3@p�g/�!?�W�s���@*�-7�ٿ�M����@aS�~��3@p�g/�!?�W�s���@*�-7�ٿ�M����@aS�~��3@p�g/�!?�W�s���@9:�u\�ٿ'���$�@r�$`E�3@_hU�!?:��7�@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@Oi�ˈ�ٿ?\�d��@�NX��3@�s�0ؐ!?�������@
�B�Y�ٿ�����@��%a��3@{.�Ǵ�!?��c���@�/���ٿ��O~�@ �4� �3@����!?�^��ܲ�@�/���ٿ��O~�@ �4� �3@����!?�^��ܲ�@�/���ٿ��O~�@ �4� �3@����!?�^��ܲ�@�/���ٿ��O~�@ �4� �3@����!?�^��ܲ�@Ƨ�c�ٿ��9��M�@��z��3@g�C��!?u�`uq��@Ƨ�c�ٿ��9��M�@��z��3@g�C��!?u�`uq��@Ƨ�c�ٿ��9��M�@��z��3@g�C��!?u�`uq��@Ƨ�c�ٿ��9��M�@��z��3@g�C��!?u�`uq��@Ƨ�c�ٿ��9��M�@��z��3@g�C��!?u�`uq��@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@I4fE�ٿ����D�@\�*�O�3@~�ǐ!?������@T��mt�ٿcL0�M�@�|"���3@�UI��!?s8Pv�w�@T��mt�ٿcL0�M�@�|"���3@�UI��!?s8Pv�w�@T��mt�ٿcL0�M�@�|"���3@�UI��!?s8Pv�w�@T��mt�ٿcL0�M�@�|"���3@�UI��!?s8Pv�w�@u �IСٿA��P�@dc���3@K��S��!?1�����@u �IСٿA��P�@dc���3@K��S��!?1�����@u �IСٿA��P�@dc���3@K��S��!?1�����@r!�Ӟٿ%�=��@R�
�S�3@#��C��!?eg.Z&�@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@���΢ٿn8?����@���?��3@[a�7ݐ!?�sR(��@����ٿ�}[��@�Q�hf�3@5��!?a�Ԟ�O�@�9�^�ٿ:�Q|ZO�@,~�c��3@і��F�!?�v�Yy��@�n�0��ٿ5��2���@���R_�3@V�\��!?\��w.[�@$��ٿA��2H�@�k/�3@,͍��!?�oq�7�@���/�ٿ��!�v��@�CF�=�3@Q)��!?��ʐ�@�7*�ٿ�l�/Z��@@�5x�3@��#�Ɛ!?V��g���@�7*�ٿ�l�/Z��@@�5x�3@��#�Ɛ!?V��g���@�7*�ٿ�l�/Z��@@�5x�3@��#�Ɛ!?V��g���@�^��ٿL��"%��@�$%�:�3@CP<���!?o�6o��@�^��ٿL��"%��@�$%�:�3@CP<���!?o�6o��@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@��گ.�ٿ��VϮ��@�յNN�3@f=���!?����M�@~X��͠ٿ�8����@�@����3@�=����!?gW�o���@~X��͠ٿ�8����@�@����3@�=����!?gW�o���@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@�I/~��ٿ킄�P��@���g�3@P۠'�!?�ry3��@ &q�(�ٿ���r*�@،����3@j�щ�!?$r�V�@D��c�ٿ"RB��M�@�>:y��3@�+U�!?���?�@D��c�ٿ"RB��M�@�>:y��3@�+U�!?���?�@,1<�ٿ�T8x��@�6�O��3@��;7͐!?1�z�B�@,1<�ٿ�T8x��@�6�O��3@��;7͐!?1�z�B�@,1<�ٿ�T8x��@�6�O��3@��;7͐!?1�z�B�@�_t��ٿ��&�@�6��3@.�|��!?�6�'�@p��A�ٿI������@q5��"�3@P�҃ɐ!?\�ߊ�@p��A�ٿI������@q5��"�3@P�҃ɐ!?\�ߊ�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@A�����ٿ4���T�@��Cu�3@���\4�!?�Vy�.�@�'�袝ٿ`q�h3��@J���v�3@w�Zr�!?Mo-%e�@����ٿ�x�vX��@ۧ6��3@&��-R�!?, 3�5�@����ٿ�x�vX��@ۧ6��3@&��-R�!?, 3�5�@����ٿ�x�vX��@ۧ6��3@&��-R�!?, 3�5�@R���K�ٿ,�CV4�@�sϩ�3@9��Y	�!?��\�H�@�^M#Ģٿ����V��@�w�U�3@��~��!?�`4��@禐)Z�ٿ��Ht(8�@N1Z�/�3@J�[���!?�oe@�T�@禐)Z�ٿ��Ht(8�@N1Z�/�3@J�[���!?�oe@�T�@禐)Z�ٿ��Ht(8�@N1Z�/�3@J�[���!?�oe@�T�@bm��1�ٿ�vҺ
B�@¨E>��3@��w��!?�d��%�@bm��1�ٿ�vҺ
B�@¨E>��3@��w��!?�d��%�@bm��1�ٿ�vҺ
B�@¨E>��3@��w��!?�d��%�@\�nצٿ��q�x��@2`�3�3@�d��j�!?!�L�4��@\�nצٿ��q�x��@2`�3�3@�d��j�!?!�L�4��@\�nצٿ��q�x��@2`�3�3@�d��j�!?!�L�4��@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@i�_`A�ٿ�#�@�@m����3@y1J���!?2_(���@�z�!�ٿ3K~��@�I@$�3@o��j��!?��.����@�z�!�ٿ3K~��@�I@$�3@o��j��!?��.����@V�;"�ٿ4[����@l!�
�3@qw�G��!?�QTb��@�IPB�ٿQ��#�@��o���3@?�&�O�!?��e*t��@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@����ٿ6�����@A�fj�3@|����!?��2"���@�&��o�ٿC���+�@}�޽]�3@�����!?gԧ"*�@����c�ٿU~{>��@6юs��3@�&w��!?Ă<Z'�@4`��ٿNN����@����M�3@�z�ơ�!?�ls��@�@4`��ٿNN����@����M�3@�z�ơ�!?�ls��@�@H��q�ٿ5>�>���@���K]�3@(]���!?zM���@'|%��ٿ��44�@Q����3@��E���!?C6� ��@/���ٿ��{����@̣���3@�_&/ܐ!?KD�	�@V�)E��ٿ�����@C����3@����k�!?��K���@V�)E��ٿ�����@C����3@����k�!?��K���@V�)E��ٿ�����@C����3@����k�!?��K���@V�)E��ٿ�����@C����3@����k�!?��K���@V�)E��ٿ�����@C����3@����k�!?��K���@"��	��ٿ}e�X��@���)��3@�d��!?�"y+wr�@k~^�ٿ�;\��	�@�ʺ��3@ΏF���!?�7Ġ	��@k~^�ٿ�;\��	�@�ʺ��3@ΏF���!?�7Ġ	��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@�9�Ϣٿ��r�*�@�L�Q�3@6�/I��!?\�?��@��j.�ٿ�$f�ԙ�@��U�1�3@���Ԑ!?2�No|�@��V�ٿ$7d��@*V(F	�3@%�M��!?�(����@��V�ٿ$7d��@*V(F	�3@%�M��!?�(����@��V�ٿ$7d��@*V(F	�3@%�M��!?�(����@��gl��ٿ��\cfA�@=vF�}�3@�U�5��!?4���3$�@�m�ٿ>{���@8H:�3@c�W`��!?�^La�@�m�ٿ>{���@8H:�3@c�W`��!?�^La�@�m�ٿ>{���@8H:�3@c�W`��!?�^La�@�m�ٿ>{���@8H:�3@c�W`��!?�^La�@�m�ٿ>{���@8H:�3@c�W`��!?�^La�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@u3�-�ٿ혫�T#�@��OWP�3@d).���!?Ԑ���R�@`�o]��ٿ�p��@�y��o�3@5&�_��!?���w��@`�o]��ٿ�p��@�y��o�3@5&�_��!?���w��@`�o]��ٿ�p��@�y��o�3@5&�_��!?���w��@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@3¬�ٿ�Ut�D��@)`�-�3@Ɛʗ��!?�qF���@	�:­�ٿ(m��{��@rP���3@�s��6�!?�tD�#�@	�:­�ٿ(m��{��@rP���3@�s��6�!?�tD�#�@@��T�ٿ��Xa��@�n���3@Db��q�!?�d�JDz�@/�Zd��ٿD�}テ�@�\��J�3@T�T.�!?�1�O�@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�����ٿ�~�1�@��� ��3@T���E�!?��]���@�Q��ٿؽn���@!����3@h$�'�!?Vh��@�Q��ٿؽn���@!����3@h$�'�!?Vh��@�Q��ٿؽn���@!����3@h$�'�!?Vh��@�Q��ٿؽn���@!����3@h$�'�!?Vh��@Z8�$�ٿo�"6��@�:=��3@�y�V��!?IU�u��@Z8�$�ٿo�"6��@�:=��3@�y�V��!?IU�u��@Z8�$�ٿo�"6��@�:=��3@�y�V��!?IU�u��@Z8�$�ٿo�"6��@�:=��3@�y�V��!?IU�u��@���K��ٿm�5%|�@lo�U��3@v<�j�!?��Wat��@���K��ٿm�5%|�@lo�U��3@v<�j�!?��Wat��@���K��ٿm�5%|�@lo�U��3@v<�j�!?��Wat��@;�ba�ٿ[�����@���"��3@�
5M��!?,6����@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@C��_Рٿz�ػ!��@��}�3@�����!?����0��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@?�N �ٿ�2����@�J���3@OQ���!?�&z&��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@:6-H~�ٿ���Xݢ�@�5k�G�3@u��Lߐ!?_O�uf��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��#�I�ٿ�gO-ɺ�@<��1�3@���E��!?#Ԙ�l��@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@��p���ٿ�#��}v�@7k�&�3@	|�ΐ!?�a�3���@(�Q��ٿe]R��@'���K�3@�ɯ���!?)����R�@(�Q��ٿe]R��@'���K�3@�ɯ���!?)����R�@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@o�F��ٿO�_`���@ g����3@��h��!?�Ψ6���@�!L���ٿ�P�.�@R�)�3@�z��!?>�<�p��@K@8�|�ٿg%���@.T�rp�3@"����!?���_�@K@8�|�ٿg%���@.T�rp�3@"����!?���_�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@7B>`��ٿ%��l�$�@j:����3@����ѐ!?�|9Y�@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�$�J��ٿ]���\�@$݇���3@,}y���!?�[����@�09�ٿ'�oO�/�@��(�3@�]�Y�!?2V!�XC�@I��4�ٿ��ݨ�@`=��5�3@��Ga�!?b�j�@I��4�ٿ��ݨ�@`=��5�3@��Ga�!?b�j�@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@��y�ʠٿ���=+�@Bcd=T�3@�5���!?��$��@8]���ٿ��D�P�@�2�Z�3@Q
�t�!?aʡ=�@8]���ٿ��D�P�@�2�Z�3@Q
�t�!?aʡ=�@�.g1ٛٿ ��)`��@=%x���3@�����!?	��Y��@�.g1ٛٿ ��)`��@=%x���3@�����!?	��Y��@�.g1ٛٿ ��)`��@=%x���3@�����!?	��Y��@.n�'�ٿtw����@�Ǳ��3@YƮ���!?�Dg���@.n�'�ٿtw����@�Ǳ��3@YƮ���!?�Dg���@.n�'�ٿtw����@�Ǳ��3@YƮ���!?�Dg���@.n�'�ٿtw����@�Ǳ��3@YƮ���!?�Dg���@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@����ٿ�/�"�@���N�3@=��_	�!?���I��@�ƶ��ٿ�F:R8�@�<����3@��j�!?���d��@�ƶ��ٿ�F:R8�@�<����3@��j�!?���d��@נ�M�ٿ�#��Y��@!��G��3@��q:ѐ!?������@נ�M�ٿ�#��Y��@!��G��3@��q:ѐ!?������@z��-��ٿUp�":7�@��]\��3@g_�K��!?�d�/]�@z��-��ٿUp�":7�@��]\��3@g_�K��!?�d�/]�@z��-��ٿUp�":7�@��]\��3@g_�K��!?�d�/]�@z��-��ٿUp�":7�@��]\��3@g_�K��!?�d�/]�@8����ٿ��ʛ��@�,���3@��5K�!?6ӛ���@M�b�ٿ�vRo��@�����3@��G��!?��;��@&��=Šٿ�P�KS�@E�^���3@�3ii1�!?'�ic-�@&��=Šٿ�P�KS�@E�^���3@�3ii1�!?'�ic-�@ɦ,�(�ٿ<��U��@���J��3@�M����!?��JT��@�)���ٿ�t��w�@��w���3@!�0��!?D{w�L�@�)���ٿ�t��w�@��w���3@!�0��!?D{w�L�@�Z��g�ٿAc���@������3@����!?~�Mi͹�@�����ٿ�?&��@q!�Z�3@����.�!?��T����@�����ٿ�?&��@q!�Z�3@����.�!?��T����@�����ٿ�?&��@q!�Z�3@����.�!?��T����@H����ٿ���a�@�|1n]�3@1����!?҇!?��@H����ٿ���a�@�|1n]�3@1����!?҇!?��@H����ٿ���a�@�|1n]�3@1����!?҇!?��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@[@�F��ٿk��t��@P���z�3@h�:�!?�kE�
��@	aj*�ٿA��o@>�@�`I�3@�ml���!?��Ѯt��@��T�p�ٿL(X��@��>���3@���yz�!?���0���@��T�p�ٿL(X��@��>���3@���yz�!?���0���@�L�!C�ٿS�N����@T���3@ڢh�q�!?��6����@�L�!C�ٿS�N����@T���3@ڢh�q�!?��6����@�L�!C�ٿS�N����@T���3@ڢh�q�!?��6����@�4�ۡٿ�,���@e�;T��3@������!?���� �@�4�ۡٿ�,���@e�;T��3@������!?���� �@A��Y��ٿ7��TVd�@����^�3@s�.��!?9QPD���@A��Y��ٿ7��TVd�@����^�3@s�.��!?9QPD���@��'(�ٿ"��!��@*]���3@�^޿�!?����%�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@XP)�ٿ���7�@R$g�3@���j��!?GگF2�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@��D�ٿ�!D�,��@Ԩ>���3@R�y�!??��=ND�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@T��I��ٿ�E����@�@���3@��ǎ�!?5�{�f�@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@��5��ٿ�$���@N�G#�3@)�!?��ɶ#��@3j��ٿU���xf�@/�>|�3@Ĉ/A��!?��o����@3j��ٿU���xf�@/�>|�3@Ĉ/A��!?��o����@3j��ٿU���xf�@/�>|�3@Ĉ/A��!?��o����@3j��ٿU���xf�@/�>|�3@Ĉ/A��!?��o����@�j}o��ٿ^��#�@tk����3@��5D��!?��y0�
�@�*�B �ٿ��%l�R�@$�Zs��3@=h���!?v�e���@�*�B �ٿ��%l�R�@$�Zs��3@=h���!?v�e���@�*�B �ٿ��%l�R�@$�Zs��3@=h���!?v�e���@�*�B �ٿ��%l�R�@$�Zs��3@=h���!?v�e���@�*�B �ٿ��%l�R�@$�Zs��3@=h���!?v�e���@�@�
�ٿz�p	�%�@I�"T\�3@��s���!?U����@ "��V�ٿN*�l���@������3@L/�ʐ!?����@ "��V�ٿN*�l���@������3@L/�ʐ!?����@ "��V�ٿN*�l���@������3@L/�ʐ!?����@ "��V�ٿN*�l���@������3@L/�ʐ!?����@ "��V�ٿN*�l���@������3@L/�ʐ!?����@lx�E�ٿB�JD�k�@�Ԯ��3@on���!?:7���@lx�E�ٿB�JD�k�@�Ԯ��3@on���!?:7���@�$k%�ٿ��]>zz�@�Ū���3@�&� ��!?=�Yz��@�$k%�ٿ��]>zz�@�Ū���3@�&� ��!?=�Yz��@�$k%�ٿ��]>zz�@�Ū���3@�&� ��!?=�Yz��@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@��w�ٿ��yQ�O�@��Y��3@h�r�!?b��6���@�o5ݠٿ�o2ö7�@Q�W��3@ke�m�!?��C�S�@�o5ݠٿ�o2ö7�@Q�W��3@ke�m�!?��C�S�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@�GF`�ٿ��ѧ�@������3@�&p|�!?���6�@s�^_��ٿ���[��@E��L	�3@;#z��!?�~���@s�^_��ٿ���[��@E��L	�3@;#z��!?�~���@s�^_��ٿ���[��@E��L	�3@;#z��!?�~���@s�^_��ٿ���[��@E��L	�3@;#z��!?�~���@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@k-�+�ٿB%CD2�@� �m��3@��U�n�!?9���__�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@���W�ٿ������@�#�v�3@t����!?��0�Ӕ�@ ^:��ٿ)IUئ	�@Lg��Y�3@��8�"�!?�ղQ��@ ^:��ٿ)IUئ	�@Lg��Y�3@��8�"�!?�ղQ��@ ^:��ٿ)IUئ	�@Lg��Y�3@��8�"�!?�ղQ��@ ^:��ٿ)IUئ	�@Lg��Y�3@��8�"�!?�ղQ��@y6��"�ٿ%e�˜;�@ɧt,��3@�<[�*�!?ݩj�ù�@y6��"�ٿ%e�˜;�@ɧt,��3@�<[�*�!?ݩj�ù�@y6��"�ٿ%e�˜;�@ɧt,��3@�<[�*�!?ݩj�ù�@y6��"�ٿ%e�˜;�@ɧt,��3@�<[�*�!?ݩj�ù�@Ug�w�ٿN�_�3�@D�hՆ�3@���2ِ!?^h����@Ug�w�ٿN�_�3�@D�hՆ�3@���2ِ!?^h����@
���ٿq����@m]G1��3@��W��!?>�/;|�@=����ٿdg�l��@�ݚ�[�3@H�hӐ!?x:ɣ���@=����ٿdg�l��@�ݚ�[�3@H�hӐ!?x:ɣ���@=����ٿdg�l��@�ݚ�[�3@H�hӐ!?x:ɣ���@=����ٿdg�l��@�ݚ�[�3@H�hӐ!?x:ɣ���@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@ܤs��ٿH����@��WTW�3@����!?����@�]�ϟٿ	s��g2�@�^��i�3@��`���!?�<��-��@�]�ϟٿ	s��g2�@�^��i�3@��`���!?�<��-��@�]�ϟٿ	s��g2�@�^��i�3@��`���!?�<��-��@]�`��ٿ~��^�@�13B�3@�I` �!?c���@]�`��ٿ~��^�@�13B�3@�I` �!?c���@]�`��ٿ~��^�@�13B�3@�I` �!?c���@&ݓ�/�ٿ
$~�6�@�:E�3@z9�ΐ!?�rCB��@���7�ٿ�"@��Y�@4���0�3@.q�ؐ!?�d�COL�@u���ٿ�,�LI��@��5�3@���Pk�!?���&�@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@*��-��ٿ�l)O��@F�ܵ�3@�#F�!?�������@�N���ٿ��$P���@�[�*��3@�M����!?��04,�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@�$N�ٿØ�����@������3@�P� ��!?��i)�:�@����ٿ�X�sN��@BwdB�3@�}�t�!?�i߹��@����ٿ�X�sN��@BwdB�3@�}�t�!?�i߹��@�A#�ٿ���R�@�`4�3@|�<��!?��%L��@OV)Q��ٿ��!�͈�@� �a�3@<�,w��!?�ݜ�=��@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@������ٿ(Q�3���@�pu�.�3@��c*ѐ!?�,���@�布Y�ٿn�0�@�@����3@�b����!?ͧ��\�@�布Y�ٿn�0�@�@����3@�b����!?ͧ��\�@�布Y�ٿn�0�@�@����3@�b����!?ͧ��\�@�布Y�ٿn�0�@�@����3@�b����!?ͧ��\�@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@n�?N��ٿX
�z/�@�(Y��3@gvԴ��!?�_˷���@��%�ٿ���Y���@��Z�3@I�qP��!?�������@��%�ٿ���Y���@��Z�3@I�qP��!?�������@�7�0�ٿأ�����@�N�C��3@5��˴�!?o� ��@�1�V�ٿ��;�A��@�qd�3@ j��z�!?�t����@�A�ܦٿ�5����@bm����3@�R�Ȓ�!?��_�F��@�A�ܦٿ�5����@bm����3@�R�Ȓ�!?��_�F��@�A�ܦٿ�5����@bm����3@�R�Ȓ�!?��_�F��@�A�ܦٿ�5����@bm����3@�R�Ȓ�!?��_�F��@D��bW�ٿ���Z��@W��54�3@tpa{�!?}U�O�@�Gn�D�ٿ�E����@�L���3@����!?�:r?�X�@~P��ٿ������@X³|.�3@����!?�
$���@�֙�d�ٿ�M��@y�@�!����3@W��!?P�Lz^��@�֙�d�ٿ�M��@y�@�!����3@W��!?P�Lz^��@�֙�d�ٿ�M��@y�@�!����3@W��!?P�Lz^��@,���ٿ�.��e�@8����3@��{��!?��{�Jd�@��S�Ԝٿ$����@ �U���3@H���!?�c�[�@��S�Ԝٿ$����@ �U���3@H���!?�c�[�@��S�Ԝٿ$����@ �U���3@H���!?�c�[�@�R�k�ٿa+6���@�c�A��3@�(�y�!?�:�@�R�k�ٿa+6���@�c�A��3@�(�y�!?�:�@=,$��ٿ�Zr�S�@/##7�3@?M���!?NH=��@8v�孠ٿ�3�G�@%�k���3@�_p��!?;�lds=�@��
��ٿ��e��)�@_�[���3@G��yߐ!?�o�g�q�@��
��ٿ��e��)�@_�[���3@G��yߐ!?�o�g�q�@��
��ٿ��e��)�@_�[���3@G��yߐ!?�o�g�q�@��
��ٿ��e��)�@_�[���3@G��yߐ!?�o�g�q�@
iN�ٿ zj�I��@:L�n�3@/9�zΐ!?B}�zj�@o��䖛ٿ��٫��@����3@e�pn��!?��e!��@(c��ٿ�q��i&�@�;z��3@�Ց��!?�~�ݩ�@�G�✣ٿ6cl1��@ð1;��3@$��Kِ!?%�	WM��@�G�✣ٿ6cl1��@ð1;��3@$��Kِ!?%�	WM��@)��ٿ��V��>�@5���?�3@�.����!?0���K��@)��ٿ��V��>�@5���?�3@�.����!?0���K��@)��ٿ��V��>�@5���?�3@�.����!?0���K��@�3���ٿ�7�5�@�O_�z�3@�׷)͐!?'J	�@��q�ٿ\4���F�@�/|��3@9Ye��!?��И���@��q�ٿ\4���F�@�/|��3@9Ye��!?��И���@��Ь[�ٿ�?�n�@X�J�3@�^�x��!?�D{�G��@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@8�n�u�ٿC5vM���@��W)u�3@�iB<z�!?9ȿ���@�}~�k�ٿ����@�@fm_�3@���ƈ�!?wA9�@�}~�k�ٿ����@�@fm_�3@���ƈ�!?wA9�@�}~�k�ٿ����@�@fm_�3@���ƈ�!?wA9�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@��b�,�ٿh�8Q�<�@�גk�3@�s1��!?=X���,�@�=��ٿ�8�����@ �, ��3@xKʐ!?E\rJ���@؁�t��ٿ)I�����@\���w�3@c�Q;ؐ!?�%y�y3�@؁�t��ٿ)I�����@\���w�3@c�Q;ؐ!?�%y�y3�@؁�t��ٿ)I�����@\���w�3@c�Q;ؐ!?�%y�y3�@�ޛu��ٿ�6�����@[o?p��3@C�J��!?{�玡��@�ޛu��ٿ�6�����@[o?p��3@C�J��!?{�玡��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@yʌ�U�ٿMS���i�@���j�3@��W;��!?����r��@�Q78�ٿvQ�;�y�@�
�ղ�3@t��t��!?��� 3�@�F�I�ٿ�|��@�J�Ӌ�3@�u*���!?]�˹��@���L�ٿ�TݓI��@4���E�3@T^G�~�!?�-�f��@���L�ٿ�TݓI��@4���E�3@T^G�~�!?�-�f��@��y\إٿ���� �@����3@���~Đ!?���7	�@��y\إٿ���� �@����3@���~Đ!?���7	�@��y\إٿ���� �@����3@���~Đ!?���7	�@'0W�~�ٿU�\���@ۭ�5N�3@��JN[�!?F�5���@'0W�~�ٿU�\���@ۭ�5N�3@��JN[�!?F�5���@'0W�~�ٿU�\���@ۭ�5N�3@��JN[�!?F�5���@H��xJ�ٿk�Ak�@�p�x&�3@��YȐ!?�{�%L�@H��xJ�ٿk�Ak�@�p�x&�3@��YȐ!?�{�%L�@H��xJ�ٿk�Ak�@�p�x&�3@��YȐ!?�{�%L�@��x�^�ٿ{��Xa�@�pL.�3@d��!?􈀪 e�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@���O��ٿ��W� �@������3@��V/��!?z#�N�a�@�[bE�ٿ��u�2�@��*Z�3@��0 (�!?cK����@�[bE�ٿ��u�2�@��*Z�3@��0 (�!?cK����@#V��ݛٿ<<����@k��Q�3@�ks��!?S�7ˠ��@��l�{�ٿ4ѯ���@q���3@$��C��!?iPq�'��@�X�-��ٿ
�,�]�@�B-��3@�Ŕ"�!?�(�Q��@�X�-��ٿ
�,�]�@�B-��3@�Ŕ"�!?�(�Q��@�5�ٿ9l�n`�@�ݤ��3@����!?H�hi���@�5�ٿ9l�n`�@�ݤ��3@����!?H�hi���@4�@�ץٿ��NW�=�@R!�M��3@T��Œ�!?%���I��@4�@�ץٿ��NW�=�@R!�M��3@T��Œ�!?%���I��@4�@�ץٿ��NW�=�@R!�M��3@T��Œ�!?%���I��@4�@�ץٿ��NW�=�@R!�M��3@T��Œ�!?%���I��@�ölh�ٿ������@�n2��3@��A��!?L ����@�ölh�ٿ������@�n2��3@��A��!?L ����@�ölh�ٿ������@�n2��3@��A��!?L ����@�ölh�ٿ������@�n2��3@��A��!?L ����@�ölh�ٿ������@�n2��3@��A��!?L ����@&�H�w�ٿ�*��@���'��3@����ِ!?v�i����@&�H�w�ٿ�*��@���'��3@����ِ!?v�i����@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@��mS�ٿ,qd��X�@?<�/��3@ʕ����!?��j��@Dh/�ٿ,Y�m��@SE�3@K��I�!?-pR?�(�@���N�ٿ�2��@��l���3@���F|�!?=���j��@���N�ٿ�2��@��l���3@���F|�!?=���j��@�`�^�ٿ5���@���y�3@v)�ӻ�!?գ2���@�`�^�ٿ5���@���y�3@v)�ӻ�!?գ2���@�`�^�ٿ5���@���y�3@v)�ӻ�!?գ2���@�`�^�ٿ5���@���y�3@v)�ӻ�!?գ2���@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@������ٿ     ��@      4@�t><K�!?��|3)��@�9����ٿ̵����@��(k��3@��l*�!?��)��@�9����ٿ̵����@��(k��3@��l*�!?��)��@�9����ٿ̵����@��(k��3@��l*�!?��)��@�I��ٿ�$J����@W���3@��v�ؐ!?w��(��@�I��ٿ�$J����@W���3@��v�ؐ!?w��(��@�I��ٿ�$J����@W���3@��v�ؐ!?w��(��@�I��ٿ�$J����@W���3@��v�ؐ!?w��(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@�b�ٿ�G���@�K&��3@�����!?�a*�(��@��R��ٿ�q@���@԰y�  4@\��̧�!?8��(��@��R��ٿ�q@���@԰y�  4@\��̧�!?8��(��@��R��ٿ�q@���@԰y�  4@\��̧�!?8��(��@��R��ٿ�q@���@԰y�  4@\��̧�!?8��(��@��R��ٿ�q@���@԰y�  4@\��̧�!?8��(��@m����ٿm6Mx���@�alF 4@�H�M�!?Gm�(��@m����ٿm6Mx���@�alF 4@�H�M�!?Gm�(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@��E	��ٿ������@kF�m��3@)�-ʐ!?�.��(��@[YS��ٿuR"����@�s�!��3@�ryِ!?=�%�(��@[YS��ٿuR"����@�s�!��3@�ryِ!?=�%�(��@[YS��ٿuR"����@�s�!��3@�ryِ!?=�%�(��@���~��ٿvS����@!����3@D�@�Ԑ!?.���(��@���~��ٿvS����@!����3@D�@�Ԑ!?.���(��@���~��ٿvS����@!����3@D�@�Ԑ!?.���(��@���~��ٿvS����@!����3@D�@�Ԑ!?.���(��@'��ٿ�G~����@}�� ��3@L����!?ˢ��(��@'��ٿ�G~����@}�� ��3@L����!?ˢ��(��@'��ٿ�G~����@}�� ��3@L����!?ˢ��(��@'��ٿ�G~����@}�� ��3@L����!?ˢ��(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�悜��ٿ������@<h�  4@}r|�Ɛ!?5�\�(��@�T��ٿ�\�����@�ڄ:  4@���Yf�!?�u�(��@�T��ٿ�\�����@�ڄ:  4@���Yf�!?�u�(��@�T��ٿ�\�����@�ڄ:  4@���Yf�!?�u�(��@�T��ٿ�\�����@�ڄ:  4@���Yf�!?�u�(��@(�=U��ٿ Iw����@7l���3@��O#�!?%��(��@(�=U��ٿ Iw����@7l���3@��O#�!?%��(��@�Hܾ�ٿ�I����@�댒  4@ۭ�0~�!?���(��@�Hܾ�ٿ�I����@�댒  4@ۭ�0~�!?���(��@�Hܾ�ٿ�I����@�댒  4@ۭ�0~�!?���(��@�Hܾ�ٿ�I����@�댒  4@ۭ�0~�!?���(��@�+����ٿ������@2�WU  4@�p��x�!?	��(��@�+����ٿ������@2�WU  4@�p��x�!?	��(��@�o}?��ٿ��b����@Bf����3@0%hN��!?HQ�(��@�����ٿ������@�W\}��3@��q�e�!?���(��@O�UL��ٿL�#����@7�g��3@�G�ѐ!?i㢵(��@O�UL��ٿL�#����@7�g��3@�G�ѐ!?i㢵(��@O�UL��ٿL�#����@7�g��3@�G�ѐ!?i㢵(��@�2�y��ٿ�|W����@�����3@g���!?X�L�(��@�2�y��ٿ�|W����@�����3@g���!?X�L�(��@�2�y��ٿ�|W����@�����3@g���!?X�L�(��@�ނC��ٿo�'����@oB����3@M��ʨ�!?��Ӵ(��@^��嵙ٿ�x����@�����3@����Ɛ!?�Ga�(��@"�����ٿzv�����@���S��3@�����!?�1��(��@"�����ٿzv�����@���S��3@�����!?�1��(��@"�����ٿzv�����@���S��3@�����!?�1��(��@"�����ٿzv�����@���S��3@�����!?�1��(��@0>�Ю�ٿ5W݋���@^^g���3@h��ݐ!?3���(��@�w~@��ٿw�����@ ����3@x�ͳ�!? ]i�(��@�w~@��ٿw�����@ ����3@x�ͳ�!? ]i�(��@eTaG��ٿ�w�����@�_LM��3@7��*�!?�=�(��@x�0��ٿ}21����@軉��3@8T{RC�!?1��(��@'�<O��ٿJ ����@CvN���3@]}fY�!?���(��@'�<O��ٿJ ����@CvN���3@]}fY�!?���(��@'�<O��ٿJ ����@CvN���3@]}fY�!?���(��@z��襙ٿKJ5����@|�9��3@��6ِ!?W)+�(��@z��襙ٿKJ5����@|�9��3@��6ِ!?W)+�(��@�]J���ٿ�����@,1M���3@DO���!?&z׹(��@�]J���ٿ�����@,1M���3@DO���!?&z׹(��@�]J���ٿ�����@,1M���3@DO���!?&z׹(��@�]J���ٿ�����@,1M���3@DO���!?&z׹(��@��q��ٿ�4�����@�^����3@�yF�!?���(��@��q��ٿ�4�����@�^����3@�yF�!?���(��@�e���ٿ4	G����@p�����3@Ֆ���!?�Eܰ(��@/�V��ٿi)����@��5���3@�Ǽ���!?9��(��@/�V��ٿi)����@��5���3@�Ǽ���!?9��(��@/�V��ٿi)����@��5���3@�Ǽ���!?9��(��@�i�6��ٿ���~���@^h�G��3@�XR�!?L?*�(��@�i�6��ٿ���~���@^h�G��3@�XR�!?L?*�(��@ЩIU��ٿ~�t|���@�yW��3@ Fپ�!?b:�(��@�Gd��ٿ�fz���@�E)��3@� 5Đ!?�':�(��@,"����ٿ�?�u���@=jI���3@�l��!?Z�z�(��@!��E��ٿ��{���@ƞ>���3@3�sL��!?����(��@!��E��ٿ��{���@ƞ>���3@3�sL��!?����(��@!��E��ٿ��{���@ƞ>���3@3�sL��!?����(��@!��E��ٿ��{���@ƞ>���3@3�sL��!?����(��@_����ٿ�L�v���@Ɋv���3@�����!?��,�(��@_����ٿ�L�v���@Ɋv���3@�����!?��,�(��@⾦Ě�ٿ|dwo���@���d��3@�'�q��!?nR��(��@⾦Ě�ٿ|dwo���@���d��3@�'�q��!?nR��(��@�Q�ە�ٿ��r���@�i��3@�^ׁ��!?�c�(��@0m4���ٿ�Vrw���@0��0��3@�l�
��!?Tt��(��@0m4���ٿ�Vrw���@0��0��3@�l�
��!?Tt��(��@0m4���ٿ�Vrw���@0��0��3@�l�
��!?Tt��(��@m����ٿ=�u���@W�u��3@�CH�!?�f�~(��@m����ٿ=�u���@W�u��3@�CH�!?�f�~(��@% Г�ٿb��u���@{�����3@�nx���!?;W(��@Z�a��ٿ�*�w���@Bc����3@R׸Ӑ!?�<�(��@_�c4��ٿ���q���@�^<��3@)�rqِ!?c��y(��@_�c4��ٿ���q���@�^<��3@)�rqِ!?c��y(��@̡]Ő�ٿowDo���@�����3@,��<��!?:�w(��@2�����ٿQ@as���@�����3@��\E�!?�A~w(��@|�j�ٿ�� p���@٨Ϝ��3@h6�!?qIx(��@|�j�ٿ�� p���@٨Ϝ��3@h6�!?qIx(��@��'��ٿWOnj���@�-�W��3@���W�!?��,j(��@-�'V��ٿ�Lkq���@�
AK��3@I��!��!?*&_m(��@���'��ٿ	\d���@�I/��3@b�6�"�!?�e�`(��@���'��ٿ	\d���@�I/��3@b�6�"�!?�e�`(��@���'��ٿ	\d���@�I/��3@b�6�"�!?�e�`(��@A�:;��ٿ��h���@@+L	��3@��G��!?i��m(��@m��8��ٿN�?e���@�J ��3@&:�߼�!?Ec�i(��@�e��ٿ6c���@�����3@i��.�!?��'f(��@��Ј��ٿ���m���@��V��3@%NP,��!?V@�k(��@��Ј��ٿ���m���@��V��3@%NP,��!?V@�k(��@��Ј��ٿ���m���@��V��3@%NP,��!?V@�k(��@g�D��ٿ?q)b���@ڄW���3@i�b&Ɛ!?L�M](��@g�D��ٿ?q)b���@ڄW���3@i�b&Ɛ!?L�M](��@������ٿ�6�d���@OP����3@V�k��!?O�[(��@������ٿ�6�d���@OP����3@V�k��!?O�[(��@�X�A��ٿ��j���@�ަ8��3@MC桐!?�M3_(��@EW����ٿ)��r���@�
���3@\L��Ɛ!?�F9r(��@rT��ٿfy���@Il���3@��b��!?Kn��(��@I�L��ٿ�BRw���@���c��3@8��PՐ!?��x(��@I�L��ٿ�BRw���@���c��3@8��PՐ!?��x(��@�\��ٿ�"����@���;��3@�H&���!?RT}�(��@�Rғ�ٿ��z���@�F(���3@�r��ڐ!?W�f�(��@��v���ٿ¦\u���@�$���3@�S�V��!?�30(��@?א�ٿi��s���@�����3@������!?<ă(��@��Bc��ٿ7g�{���@��#P��3@�R���!?����(��@�!Ǫ��ٿF��|���@�1��3@	w�l��!?��K�(��@�qku��ٿ��}|���@7���3@���氐!?_�(��@r!�瘙ٿ�:ك���@������3@�Q�+��!?i��(��@�3-ӗ�ٿ:��}���@�q���3@�5�&��!?�X �(��@7�J���ٿQ!�{���@�����3@e���!?��v�(��@�8����ٿ�O|���@Wn���3@u/���!?�5�(��@X����ٿO8�{���@T����3@LUP�Đ!?�oͯ(��@�`�d��ٿ�����@������3@�Z���!?+���(��@O�s��ٿ��s����@�q�=��3@�xp��!?+���(��@u���ٿI*ۀ���@�����3@#��
�!?D{��(��@��9��ٿԽ�w���@�9���3@TWӪ8�!?�w��(��@��9��ٿԽ�w���@�9���3@TWӪ8�!?�w��(��@��9��ٿԽ�w���@�9���3@TWӪ8�!?�w��(��@��9��ٿԽ�w���@�9���3@TWӪ8�!?�w��(��@��9��ٿԽ�w���@�9���3@TWӪ8�!?�w��(��@�e����ٿ%�p{���@��3���3@�e�9�!?��(��@KQJ3��ٿ64����@�Yq��3@�� wD�!?k�	�(��@R⋞�ٿ-��~���@�����3@�<�� �!?�)�(��@R⋞�ٿ-��~���@�����3@�<�� �!?�)�(��@���(��ٿ��{���@[�`���3@rT�� �!?]���(��@���(��ٿ��{���@[�`���3@rT�� �!?]���(��@=�c���ٿi��y���@R�����3@&�S7�!?�M��(��@Wl|���ٿ�lwr���@��}���3@wD�s��!?���(��@�Z��ٿD+�k���@����3@I�._�!?H��(��@�Ue���ٿ�jm���@���C��3@�E��!?"B��(��@��ٿ���l���@��2z��3@B�E�ې!?�JX�(��@�crƇ�ٿ�.�b���@Qh��3@�����!?���(��@_����ٿ���g���@�	��3@�= ��!?�Ѯ(��@x�C��ٿEa���@�;xd��3@�.'�Z�!?qKx�(��@x�C��ٿEa���@�;xd��3@�.'�Z�!?qKx�(��@^�;�}�ٿ+O�`���@;���3@�Гk�!?=�"�(��@�(�l{�ٿN��]���@"���3@�F;d��!?A�I�(��@�u�*}�ٿ�i]���@Շ����3@1.+M͐!?zO�(��@�T2�|�ٿ��[���@1W���3@������!?FV��(��@��v�w�ٿ���X���@�pM���3@������!?WU��(��@��v�w�ٿ���X���@�pM���3@������!?WU��(��@�C&�m�ٿ��M���@�=y#��3@�= ��!?�)h�(��@�x
�c�ٿe�!C���@+�u��3@�*.ߐ!?[R�(��@��^j�ٿ	hRK���@3=����3@�N�x�!?)! �(��@ *��k�ٿ�G���@���3@>�ݙ�!?wt��(��@0 �m�ٿvg�E���@
��T��3@��3���!?���(��@0 �m�ٿvg�E���@
��T��3@��3���!?���(��@0 �m�ٿvg�E���@
��T��3@��3���!?���(��@z#��y�ٿ�T���@,���3@]VSc.�!?�5��(��@�H^m��ٿ��Hc���@�P����3@�rO1 �!?.�=�(��@�H^m��ٿ��Hc���@�P����3@�rO1 �!?.�=�(��@S:C9��ٿRL�[���@����3@PO�z�!?����(��@�y,�~�ٿ�G�V���@.����3@ؿmJސ!?���(��@�y,�~�ٿ�G�V���@.����3@ؿmJސ!?���(��@j�:ri�ٿ�\�@���@[kQ:��3@bA��!?��y�(��@j�:ri�ٿ�\�@���@[kQ:��3@bA��!?��y�(��@j�:ri�ٿ�\�@���@[kQ:��3@bA��!?��y�(��@j�:ri�ٿ�\�@���@[kQ:��3@bA��!?��y�(��@j�:ri�ٿ�\�@���@[kQ:��3@bA��!?��y�(��@�e�h�ٿ��y=���@(�����3@aˌ0�!?�c��(��@Iគi�ٿGo?���@�1��3@t���!?��f�(��@Iគi�ٿGo?���@�1��3@t���!?��f�(��@�d��l�ٿ�"E���@������3@��«
�!?� Y�(��@�s�_i�ٿJ�EF���@-�q���3@*v#��!?D�?�(��@g���r�ٿ|�4Q���@[����3@�^!?!U�(��@ݬ�||�ٿy��a���@/�E��3@ʻ߀��!?�
�(��@Z��腙ٿ%(�m���@�Z����3@X*qI}�!?o^(��@�h�늙ٿfln���@��Y��3@��!�ǐ!?��N�(��@9|:��ٿ�ʈl���@B[u��3@�����!?�f��(��@�ڈ�u�ٿwՓY���@�l8m��3@��TJ��!?�2٬(��@�ڈ�u�ٿwՓY���@�l8m��3@��TJ��!?�2٬(��@�ڈ�u�ٿwՓY���@�l8m��3@��TJ��!?�2٬(��@���n�ٿ*��O���@��u��3@p:���!?��ٺ(��@��n�ٿ�FO���@ �
r��3@���!?����(��@C�_�ٿq:���@́����3@���!?��)��@���u�ٿ���T���@n����3@�Ds��!?_r��(��@���u�ٿ���T���@n����3@�Ds��!?_r��(��@�铖��ٿ�{�`���@�+:5��3@O�����!?(��(��@���j�ٿ	�F���@W�����3@�j���!?�w�)��@D��\i�ٿ�a J���@A���3@�G\�Ɛ!?e�G�(��@)��k�ٿ=o>N���@����3@�%=�ǐ!?��P�(��@�q�\�ٿ�|�?���@d�����3@`7@ѯ�!?Vn�(��@�q�\�ٿ�|�?���@d�����3@`7@ѯ�!?Vn�(��@I��Z�ٿ�[B���@�9����3@uo�j�!?r3X�(��@�Y0vU�ٿ��B���@�����3@�4�t�!?:J��(��@E�sV�ٿI��?���@S�����3@�Kઐ!?���(��@E�sV�ٿI��?���@S�����3@�Kઐ!?���(��@�%L�J�ٿ��R:���@#����3@<���!?�M��(��@�%L�J�ٿ��R:���@#����3@<���!?�M��(��@K�^�R�ٿ�?���@8�lI��3@Þg^��!?IΆ�(��@K�^�R�ٿ�?���@8�lI��3@Þg^��!?IΆ�(��@K�^�R�ٿ�?���@8�lI��3@Þg^��!?IΆ�(��@K�^�R�ٿ�?���@8�lI��3@Þg^��!?IΆ�(��@`
1>�ٿt�/+���@�����3@l�4���!?�Eb�(��@��w�G�ٿ��a4���@��L��3@"��Up�!?�!�(��@j ?�ٿӶp*���@�~����3@k�
'n�!?a9�(��@j ?�ٿӶp*���@�~����3@k�
'n�!?a9�(��@�O�W�ٿǀ�:���@ t,��3@WgwR��!?C1h�(��@�dDGX�ٿ�ǩ/���@Aԑ���3@N�|6ʐ!?��$)��@L��D�ٿjŊ���@���K��3@���Ŵ�!?1��/)��@L��D�ٿjŊ���@���K��3@���Ŵ�!?1��/)��@�6�N�ٿ�m,���@���s��3@�Pw���!?�C	�(��@�6�N�ٿ�m,���@���s��3@�Pw���!?�C	�(��@h+4�?�ٿ�u���@�A���3@�Hű֐!?wU�
)��@u\_�*�ٿ.�����@�����3@�2^��!?�\�()��@l��E�ٿ������@�sU}��3@Os���!?ߪ�')��@l��E�ٿ������@�sU}��3@Os���!?ߪ�')��@�oQ��ٿ\s����@8�c��3@VU��!?���1)��@�z�՘ٿ{V�����@��v���3@SE6D��!?�}�8)��@�
g�ܘٿ�PO����@ȣ�r��3@�_1D�!?O�/)��@X�b�ٿ ������@������3@��!4�!?.�')��@R��8H�ٿB���@2�����3@�����!?����(��@R��8H�ٿB���@2�����3@�����!?����(��@R��8H�ٿB���@2�����3@�����!?����(��@���i0�ٿ��A
���@�o���3@Uй�ڐ!?���(��@��Z5�ٿ�����@�����3@Դ��!?�VD�(��@-�2�ٿ��}���@	&+���3@Z��	�!?q$1)��@-�2�ٿ��}���@	&+���3@Z��	�!?q$1)��@-�2�ٿ��}���@	&+���3@Z��	�!?q$1)��@A�w�/�ٿ�e����@��J��3@�B9�!?����(��@�?90@�ٿ�u##���@.9����3@�y���!?y�;
)��@�?90@�ٿ�u##���@.9����3@�y���!?y�;
)��@�?90@�ٿ�u##���@.9����3@�y���!?y�;
)��@�?90@�ٿ�u##���@.9����3@�y���!?y�;
)��@�?90@�ٿ�u##���@.9����3@�y���!?y�;
)��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@#eͰ.�ٿ
����@,[����3@K�ԅ��!?�l�))��@Ө ��ٿ�E����@�?����3@9����!?t$\)��@��=B�ٿ�i�����@���i��3@�:�D��!?�1|r)��@Id���ٿWa\����@V�%���3@8�N�ߐ!?{zm�)��@G*ژٿq�s����@�v="��3@;L|�!?�L��)��@W���ٿO�j����@}���3@�X�8�!?9�:�)��@W���ٿO�j����@}���3@�X�8�!?9�:�)��@���ޘٿ6�&����@�4x���3@&��/�!?�S�)��@� k�јٿ������@��{���3@T�K�9�!?�s��)��@�N�"��ٿST�����@<M����3@3��!?�AD�)��@@?��Řٿ�t����@�Y����3@%��y��!?�i��)��@U��|�ٿx��d���@�#���3@m=/��!?QW�*��@U��|�ٿx��d���@�#���3@m=/��!?QW�*��@�<��+�ٿ���@�k"��3@}g����!?�7}*��@�ik��ٿ������@��a��3@_Ʋ���!?@�h +��@�ik��ٿ������@��a��3@_Ʋ���!?@�h +��@�~��ٿ O_����@������3@2�O���!?ر��*��@��Q�(�ٿ�>]���@oa&��3@4y�=�!?��_*��@��Q�(�ٿ�>]���@oa&��3@4y�=�!?��_*��@��Q�(�ٿ�>]���@oa&��3@4y�=�!?��_*��@�����ٿ�t����@)1!��3@!	Q:�!?mO�*��@�����ٿ�t����@)1!��3@!	Q:�!?mO�*��@��ͳ�ٿw�����@=�HL��3@�~q|'�!?��ȶ*��@��ͳ�ٿw�����@=�HL��3@�~q|'�!?��ȶ*��@�l�:6�ٿ������@�q1���3@&��3�!?J`�H*��@@6T85�ٿ�Vt!���@F6O��3@��@��!?�1�5*��@@6T85�ٿ�Vt!���@F6O��3@��@��!?�1�5*��@@6T85�ٿ�Vt!���@F6O��3@��@��!?�1�5*��@@6T85�ٿ�Vt!���@F6O��3@��@��!?�1�5*��@?�kV��ٿ`��r���@M����3@�EZ&��!?��*��@?�kV��ٿ`��r���@M����3@�EZ&��!?��*��@�����ٿ��s����@>�6
��3@�8�mb�!?Z��)��@�����ٿ��s����@>�6
��3@�8�mb�!?Z��)��@�ihn�ٿP�Q���@P3��3@�DI`��!?�6�H*��@� +ޤ�ٿ������@�`�>��3@+�nr��!?�v�.+��@�<S�ٿj�N����@������3@��!?K��*��@���g�ٿ"�\C���@-7���3@H[^�?�!?)�!*��@	�Pz&�ٿ�{����@�>����3@�oErn�!?��#Q*��@	�Pz&�ٿ�{����@�>����3@�oErn�!?��#Q*��@	�Pz&�ٿ�{����@�>����3@�oErn�!?��#Q*��@��+�ٿR�����@��5}��3@���7��!?Ӽ7*��@��+�ٿR�����@��5}��3@���7��!?Ӽ7*��@���}g�ٿI=$C���@XW����3@�����!?�~ۿ)��@��+?�ٿ�u3����@�y��3@��Ա��!?I�|*��@
cj��ٿ��q���@�� ���3@ ��
�!?��d�*��@Y� ��ٿ��7����@@����3@����I�!?�e��*��@Y� ��ٿ��7����@@����3@����I�!?�e��*��@Y� ��ٿ��7����@@����3@����I�!?�e��*��@w�@P�ٿ¯�����@�z	���3@�Cg�ɐ!?��|�*��@S:�a�ٿ�j(Z���@�����3@��]3�!?A�R�)��@ i�ٿ������@�����3@C6|�!?i�Ea*��@�;%˘ٿWx����@J����3@l�BА!?�^�)��@�;%˘ٿWx����@J����3@l�BА!?�^�)��@�d��-�ٿm=T���@ޕ���3@��'��!?i���(��@�wrӘٿTW����@�����3@�O�ǐ!?Cb-)��@�wrӘٿTW����@�����3@�O�ǐ!?Cb-)��@�wrӘٿTW����@�����3@�O�ǐ!?Cb-)��@v�ۗٿ�������@�g����3@��]А!?���*��@vR.X˗ٿ{�����@�l���3@���˕�!?OV�0*��@� ���ٿ܉{����@�s*���3@L��B��!?����)��@Z�iHٿ������@e�<��3@%��g��!?�d��(��@4RjaS�ٿ�o�7���@�-���3@�c�C��!?0%�)��@"3����ٿ��}���@����3@�k���!?���(��@�0gX��ٿ��T����@|l����3@�	W���!?Z�}(��@�0gX��ٿ��T����@|l����3@�	W���!?Z�}(��@� h��ٿآ����@�
����3@�##Ր!?�%��'��@�𻟘ٿ�ɋ|���@,,mU��3@�`�O��!?FPSl'��@1V�s�ٿ3Y�F���@��
 4@��w��!?J��}&��@�Z�+�ٿ�� ��@�^�? 4@�yG��!?.Da&��@�Z�+�ٿ�� ��@�^�? 4@�yG��!?.Da&��@bD����ٿ�{����@oS� 4@�V.���!?���&��@bD����ٿ�{����@oS� 4@�V.���!?���&��@bD����ٿ�{����@oS� 4@�V.���!?���&��@bD����ٿ�{����@oS� 4@�V.���!?���&��@���X�ٿ#J�?���@�	�	 4@e��y�!?jX�(��@��b̷�ٿ�h����@l���	 4@�]2ٯ�!?b�+'��@��b̷�ٿ�h����@l���	 4@�]2ٯ�!?b�+'��@ҭ\Иٿ������@�����3@��HÐ!?{'�@)��@v�3�ڗٿ3�@����@������3@���c�!?Bv�)��@v�3�ڗٿ3�@����@������3@���c�!?Bv�)��@v�3�ڗٿ3�@����@������3@���c�!?Bv�)��@�`��z�ٿ%�0a���@�
�= 4@�?^v�!?|p9-'��@�`��z�ٿ%�0a���@�
�= 4@�?^v�!?|p9-'��@�� �ٿ������@��� 4@8�y���!?�K�&��@�� �ٿ������@��� 4@8�y���!?�K�&��@��A��ٿx�{���@3_���3@\��!?.L'�(��@�̬a{�ٿzm?`���@�d���3@�L*qɐ!?\M�(��@�̬a{�ٿzm?`���@�d���3@�L*qɐ!?\M�(��@u��J�ٿ	�����@З���3@0Ó���!?K�q*��@u��J�ٿ	�����@З���3@0Ó���!?K�q*��@u��J�ٿ	�����@З���3@0Ó���!?K�q*��@u��J�ٿ	�����@З���3@0Ó���!?K�q*��@�e-���ٿKgk����@[U$��3@p�_���!?���+(��@��햘ٿC2|w���@�����3@ϡ���!?��)��@ӛ��ٿ9������@�r<���3@=>JKߐ!?�p��+��@͡����ٿ�������@�K���3@�����!?#���,��@.`��f�ٿ7S�����@�m\��3@R���!?�0��@$mY��ٿMc�����@)'���3@JP3�!?��c�*��@$mY��ٿMc�����@)'���3@JP3�!?��c�*��@�>GY�ٿp��,���@e/�W��3@ ��ː!?�cB.��@[��c��ٿ�F� ��@!����3@�t���!?p�Ԩ0��@��M�@�ٿ*��j���@ 1�n��3@�����!?.���1��@:����ٿ��~8��@rj�T��3@��Kh�!?@��u0��@:����ٿ��~8��@rj�T��3@��Kh�!?@��u0��@:����ٿ��~8��@rj�T��3@��Kh�!?@��u0��@:����ٿ��~8��@rj�T��3@��Kh�!?@��u0��@�V`��ٿ+0���@2~Q��3@��Iх�!?��?1��@h>���ٿ�]�p��@�aQ< 4@ ŋgo�!?����(��@'� t�ٿ��6���@OJ$��3@dvXԒ�!?Ř��-��@�;şٿU'ߺ��@���� 4@�����!?���)��@����a�ٿ���;��@^5� 4@h�����!?[U�x'��@����a�ٿ���;��@^5� 4@h�����!?[U�x'��@p� �ٿRM]���@��j" 4@Q�WYܐ!?�72))��@=}����ٿ����@��� 4@��u��!?��)��@=}����ٿ����@��� 4@��u��!?��)��@?��o{�ٿ�v�*��@?��2 4@h0H��!?\�\%��@%��
�ٿ&d��	��@Z�, 4@,&Đ!?:GD�(��@Ө���ٿ��"��@��n�( 4@���!?�h�+��@Ө���ٿ��"��@��n�( 4@���!?�h�+��@Ө���ٿ��"��@��n�( 4@���!?�h�+��@Ө���ٿ��"��@��n�( 4@���!?�h�+��@Ө���ٿ��"��@��n�( 4@���!?�h�+��@c-�F�ٿ�vKB��@o��� 4@�;�䖐!?"i$�)��@c-�F�ٿ�vKB��@o��� 4@�;�䖐!?"i$�)��@b�w��ٿ�=>���@��� 4@����!?��LE(��@b�w��ٿ�=>���@��� 4@����!?��LE(��@L�}"�ٿ<����@�^f� 4@��q��!?�@*��@L�}"�ٿ<����@�^f� 4@��q��!?�@*��@L�}"�ٿ<����@�^f� 4@��q��!?�@*��@L�}"�ٿ<����@�^f� 4@��q��!?�@*��@L�}"�ٿ<����@�^f� 4@��q��!?�@*��@�M��m�ٿ�A`g��@�2 4@M���Ȑ!?�)�i+��@�M��m�ٿ�A`g��@�2 4@M���Ȑ!?�)�i+��@�M��m�ٿ�A`g��@�2 4@M���Ȑ!?�)�i+��@�M��m�ٿ�A`g��@�2 4@M���Ȑ!?�)�i+��@�̫Io�ٿB��H��@
V�� 4@YvY��!?e�&��@��x�0�ٿ7�`
��@y��� 4@v��{�!?��m�/��@a���0�ٿg23W	��@-i�� 4@>%ío�!?6Du/��@�>w�ٿ��o���@� ���3@�/o���!?#���-��@�>w�ٿ��o���@� ���3@�/o���!?#���-��@�>w�ٿ��o���@� ���3@�/o���!?#���-��@�>w�ٿ��o���@� ���3@�/o���!?#���-��@��ߏ�ٿ�=��
��@X�̷��3@|G����!?Y��Z4��@����ٿ|�$��@9�pq��3@��|Ɛ!?	\�0��@����ٿ|�$��@9�pq��3@��|Ɛ!?	\�0��@����ٿ|�$��@9�pq��3@��|Ɛ!?	\�0��@����ٿ|�$��@9�pq��3@��|Ɛ!?	\�0��@����ٿ|�$��@9�pq��3@��|Ɛ!?	\�0��@ ��ׯ�ٿA�ļ��@V����3@�ӡp�!?J�!-��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@� ޘٿh�ۣ���@)�[`��3@%&o�!?OTr�'��@n�w*��ٿ|I2��@���4��3@��.\ɐ!?�]�z4��@� ��ٿ反.���@=�����3@��5!?y��7.��@� ��ٿ反.���@=�����3@��5!?y��7.��@d%y�3�ٿRT����@<�e���3@����f�!?YD��4��@d%y�3�ٿRT����@<�e���3@����f�!?YD��4��@d��)�ٿ�gm��@'l����3@I���l�!?'.z�2��@d��)�ٿ�gm��@'l����3@I���l�!?'.z�2��@d��)�ٿ�gm��@'l����3@I���l�!?'.z�2��@d��)�ٿ�gm��@'l����3@I���l�!?'.z�2��@d��)�ٿ�gm��@'l����3@I���l�!?'.z�2��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@<�#/��ٿ�E��	��@P�����3@4"8T�!?�!�6��@h����ٿ�����@ﮕ���3@D�)ӥ�!?�-�6��@h����ٿ�����@ﮕ���3@D�)ӥ�!?�-�6��@O;�hp�ٿ�j���@0M��3@# ��!?=z�f7��@O;�hp�ٿ�j���@0M��3@# ��!?=z�f7��@O;�hp�ٿ�j���@0M��3@# ��!?=z�f7��@O;�hp�ٿ�j���@0M��3@# ��!?=z�f7��@.�����ٿ Sˠ ��@U�/�4 4@Jt�m�!?���i"��@.�����ٿ Sˠ ��@U�/�4 4@Jt�m�!?���i"��@.�����ٿ Sˠ ��@U�/�4 4@Jt�m�!?���i"��@.�����ٿ Sˠ ��@U�/�4 4@Jt�m�!?���i"��@�ʧ]I�ٿ�Ĕ����@	���/ 4@�9�H��!?�� ��@9F�!�ٿm�C��@���L��3@�Xħ�!?�Ҥ4��@9F�!�ٿm�C��@���L��3@�Xħ�!?�Ҥ4��@�v9J��ٿ���'��@���v�3@x�8���!?��=��@�u�ٿ�J���@�����3@�6�7�!?��'�L��@zԵ��ٿjh/���@[����3@T	���!?��$�Y��@Ľ'�ٿG�b%��@O�&�e�3@ڈo�m�!?<uvi��@F�����ٿ6��)��@QN��3@EJ��B�!?�xG�t��@F�����ٿ6��)��@QN��3@EJ��B�!?�xG�t��@����ٿ�Ŝ��@g���3@5�+�ؐ!?��/�s��@����ٿ�Ŝ��@g���3@5�+�ؐ!?��/�s��@����ٿ�Ŝ��@g���3@5�+�ؐ!?��/�s��@u��wK�ٿ�uP
��@�ʾ�3@)��X�!?�*�Q[��@u��wK�ٿ�uP
��@�ʾ�3@)��X�!?�*�Q[��@�\�nƛٿX�T���@?�����3@��)��!?��E3��@	��wM�ٿr�g���@�}~F�3@�rM�c�!?ɚHfE��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@����O�ٿ��M��@�� 4@�rM��!?p�|�(��@�M9]�ٿԥh,��@���g��3@-P����!?=d�X��@~RE�P�ٿ�T�	��@�>��$�3@�c��!?��(O��@~RE�P�ٿ�T�	��@�>��$�3@�c��!?��(O��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@��HR�ٿkAZ���@���]D�3@�gyא!?�c�L��@�ꨢٿm�����@�bܜ�3@�#�ؐ!?.f��A��@�ꨢٿm�����@�bܜ�3@�#�ؐ!?.f��A��@�ꨢٿm�����@�bܜ�3@�#�ؐ!?.f��A��@�ꨢٿm�����@�bܜ�3@�#�ؐ!?.f��A��@�ꨢٿm�����@�bܜ�3@�#�ؐ!?.f��A��@ѽ�;��ٿ*����@��P�3@ԙ��*�!?���Q��@ѽ�;��ٿ*����@��P�3@ԙ��*�!?���Q��@ѽ�;��ٿ*����@��P�3@ԙ��*�!?���Q��@�x!/�ٿ� �4 ��@H�r��3@�a46ސ!?:���H��@�x!/�ٿ� �4 ��@H�r��3@�a46ސ!?:���H��@�x!/�ٿ� �4 ��@H�r��3@�a46ސ!?:���H��@�gbΞ�ٿW��	��@���(��3@t�xNp�!? ��u��@�gbΞ�ٿW��	��@���(��3@t�xNp�!? ��u��@�gbΞ�ٿW��	��@���(��3@t�xNp�!? ��u��@�gbΞ�ٿW��	��@���(��3@t�xNp�!? ��u��@�8%NA�ٿ'h���@SRU�
�3@��*!�!?���gk��@�8%NA�ٿ'h���@SRU�
�3@��*!�!?���gk��@�8%NA�ٿ'h���@SRU�
�3@��*!�!?���gk��@�8%NA�ٿ'h���@SRU�
�3@��*!�!?���gk��@�*�F�ٿ$��f��@J�ŭ;�3@�+���!?+�	?��@_O�j�ٿ������@yZ���3@��vܐ!?�.8/��@_O�j�ٿ������@yZ���3@��vܐ!?�.8/��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@���f�ٿDi����@$�ʓp�3@w��
�!?�q{�]��@�)��e�ٿ]+���@. ��3@�α��!?���HW��@����ٿ�!���@c��3@�D2	�!?e�r.���@����ٿ�!���@c��3@�D2	�!?e�r.���@����ٿ�!���@c��3@�D2	�!?e�r.���@����ٿ�!���@c��3@�D2	�!?e�r.���@����ٿ�!���@c��3@�D2	�!?e�r.���@q��ٿ!>9���@��C��3@="ы��!?���?��@q��ٿ!>9���@��C��3@="ы��!?���?��@q��ٿ!>9���@��C��3@="ы��!?���?��@q��ٿ!>9���@��C��3@="ы��!?���?��@v]�ٿҺ���@?Kd��3@�8�쐐!?�;H��@���L�ٿ�����@c�wN�3@G_��!?�Qh����@R�4l(�ٿQ�q���@?A�K��3@��=�ǐ!?ͳ����@gN��G�ٿ�oM���@�E�A�3@P���!?[+����@gN��G�ٿ�oM���@�E�A�3@P���!?[+����@gN��G�ٿ�oM���@�E�A�3@P���!?[+����@h��eӡٿ�p�D
��@�J�3@_s��!?�Ѣf���@j�s�2�ٿM(���@%BsZ��3@�mz}�!?l:f���@j�s�2�ٿM(���@%BsZ��3@�mz}�!?l:f���@j�s�2�ٿM(���@%BsZ��3@�mz}�!?l:f���@j�s�2�ٿM(���@%BsZ��3@�mz}�!?l:f���@�.>�@�ٿC,J4��@)k����3@uT"`�!?�>f<���@�.>�@�ٿC,J4��@)k����3@uT"`�!?�>f<���@�.>�@�ٿC,J4��@)k����3@uT"`�!?�>f<���@$_0I��ٿ;����@4���3@�DL���!?�n����@$_0I��ٿ;����@4���3@�DL���!?�n����@$_0I��ٿ;����@4���3@�DL���!?�n����@$_0I��ٿ;����@4���3@�DL���!?�n����@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@Oj{�ٿ�y��@�ڡ�<�3@X��E�!?��>i3��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@:�n�+�ٿ#U��@�dM�{�3@ۜ����!?�9�:��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@�*�Ӡ�ٿ�B�-��@x-�3@S�gА!?uoH0��@ደW�ٿ~�o&��@��?�3@����+�!?�0�����@/���ٿ�#A���@�E(wx�3@^<s�q�!?\�?����@@B[�Y�ٿo�:���@c�R5Z�3@��~Ð!?�'D%��@@B[�Y�ٿo�:���@c�R5Z�3@��~Ð!?�'D%��@@B[�Y�ٿo�:���@c�R5Z�3@��~Ð!?�'D%��@@B[�Y�ٿo�:���@c�R5Z�3@��~Ð!?�'D%��@@B[�Y�ٿo�:���@c�R5Z�3@��~Ð!?�'D%��@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@{�:?�ٿ�ءV��@�lM'��3@�PD`��!?98z���@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@d{�-��ٿ9�
��@G[�~��3@n�{���!?s@3�^��@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@��Z|��ٿsU���@|��?&�3@=W�
ې!?�sQ����@A�sw��ٿ�"3�
��@����3@6T�zk�!?t	/Z���@A�sw��ٿ�"3�
��@����3@6T�zk�!?t	/Z���@A�sw��ٿ�"3�
��@����3@6T�zk�!?t	/Z���@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@!�#�ٿ��w���@1s���3@���Z�!?�	t��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@���ܞٿ%\����@�ݨ�W�3@c�MG�!?Y���V��@����ٿ�[����@��Ћ��3@޵�A�!?&�V����@�3�UR�ٿ'�?���@�u(b�3@�*���!?_,Z���@�3�UR�ٿ'�?���@�u(b�3@�*���!?_,Z���@�3�UR�ٿ'�?���@�u(b�3@�*���!?_,Z���@Ur��ٿ.�����@� e��3@2�$}֐!?����+��@Ur��ٿ.�����@� e��3@2�$}֐!?����+��@�&���ٿ��G���@ ����3@y|>��!?V�_���@�&���ٿ��G���@ ����3@y|>��!?V�_���@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@�Ϋ(�ٿ�����@jqY��3@B^��ݐ!?��&Rs��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@��E�ٿR�G���@�Rl��3@Q�O��!?�13��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@�%�Y�ٿ���.��@�r;�3@v@���!?���y��@~��|�ٿ_p�>��@:�"�3@���!?b�����@~��|�ٿ_p�>��@:�"�3@���!?b�����@~��|�ٿ_p�>��@:�"�3@���!?b�����@��ٿ�d�}��@��*��3@{�Ĥ�!?֝_t���@��JM�ٿ���Q��@\i�m��3@��D$�!?���v��@��JM�ٿ���Q��@\i�m��3@��D$�!?���v��@S����ٿ.9
��@��{��3@�L���!?L�hq��@�T:��ٿ��j�
��@�i,��3@�3qؐ!?������@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@��)�ٿ]R�D��@o��by�3@X�M�!?���Y��@5��eԢٿA����@���PW�3@���f�!?+��Z��@5��eԢٿA����@���PW�3@���f�!?+��Z��@5��eԢٿA����@���PW�3@���f�!?+��Z��@5��eԢٿA����@���PW�3@���f�!?+��Z��@5��eԢٿA����@���PW�3@���f�!?+��Z��@5��eԢٿA����@���PW�3@���f�!?+��Z��@�Z�sI�ٿ�%8���@I�q$�3@+x��!?dm�D ��@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@�|j��ٿD����@M��o��3@���Ӑ!?�	*���@o`�ҷ�ٿ������@\�c��3@�����!?A�����@o`�ҷ�ٿ������@\�c��3@�����!?A�����@VPb&��ٿˈAz��@ �D_K�3@��Ff�!?L`?	��@VPb&��ٿˈAz��@ �D_K�3@��Ff�!?L`?	��@VPb&��ٿˈAz��@ �D_K�3@��Ff�!?L`?	��@VPb&��ٿˈAz��@ �D_K�3@��Ff�!?L`?	��@VPb&��ٿˈAz��@ �D_K�3@��Ff�!?L`?	��@���ՓٿW����@�j�M��3@�f��o�!?J1�����@���ՓٿW����@�j�M��3@�f��o�!?J1�����@���ՓٿW����@�j�M��3@�f��o�!?J1�����@���ՓٿW����@�j�M��3@�f��o�!?J1�����@z6��ٿ�P>��@��{��3@�[ ��!?������@z6��ٿ�P>��@��{��3@�[ ��!?������@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@�r�5��ٿ�g�����@����3@��&I	�!?�"�s��@F_x�Ĝٿ�� ��@̠���3@[�񑿐!?9���]��@F_x�Ĝٿ�� ��@̠���3@[�񑿐!?9���]��@F_x�Ĝٿ�� ��@̠���3@[�񑿐!?9���]��@�l�F{�ٿ$�j��@CW\-�3@���=��!?+,,���@�l�F{�ٿ$�j��@CW\-�3@���=��!?+,,���@�l�F{�ٿ$�j��@CW\-�3@���=��!?+,,���@�l�F{�ٿ$�j��@CW\-�3@���=��!?+,,���@�l�F{�ٿ$�j��@CW\-�3@���=��!?+,,���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@���|�ٿ,r�@��@ٷ�s�3@� )S��!?+E���@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@�/5j�ٿ5w}��@?!�+��3@KzǗ�!?��Iay��@��1�ٿ�s���@�]5b�3@�ڣ���!?\�0"���@IQ�r�ٿh����@��S5�3@띤dg�!?���x��@IQ�r�ٿh����@��S5�3@띤dg�!?���x��@IQ�r�ٿh����@��S5�3@띤dg�!?���x��@IQ�r�ٿh����@��S5�3@띤dg�!?���x��@IQ�r�ٿh����@��S5�3@띤dg�!?���x��@�6��؜ٿFnv���@P��Y�3@��=\��!?b� ���@�A���ٿ�u����@д��1�3@�EWOҐ!?q�t����@�A���ٿ�u����@д��1�3@�EWOҐ!?q�t����@�A���ٿ�u����@д��1�3@�EWOҐ!?q�t����@4���ٿeaު	��@1����3@_{�!��!?������@4���ٿeaު	��@1����3@_{�!��!?������@4���ٿeaު	��@1����3@_{�!��!?������@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@���S�ٿ��!K��@��3@u���!?��zTh��@³�Z�ٿ&c@>��@*a��3@ޢ�گ�!?M���o��@³�Z�ٿ&c@>��@*a��3@ޢ�گ�!?M���o��@³�Z�ٿ&c@>��@*a��3@ޢ�گ�!?M���o��@³�Z�ٿ&c@>��@*a��3@ޢ�گ�!?M���o��@�A�T�ٿBcb���@a��K_�3@vb��!?!��8���@���1Ѣٿ�>���@+N���3@��ȏ�!?�rj|���@��m���ٿ"����@'�3F�3@k��`��!?<e8���@��m���ٿ"����@'�3F�3@k��`��!?<e8���@��m���ٿ"����@'�3F�3@k��`��!?<e8���@��m���ٿ"����@'�3F�3@k��`��!?<e8���@��m���ٿ"����@'�3F�3@k��`��!?<e8���@�g�ٿ|���@۞�X��3@���0ِ!?8ӝ���@�g�ٿ|���@۞�X��3@���0ِ!?8ӝ���@��c��ٿ (y���@x����3@�gi�ې!?`��5���@��c��ٿ (y���@x����3@�gi�ې!?`��5���@��c��ٿ (y���@x����3@�gi�ې!?`��5���@��c��ٿ (y���@x����3@�gi�ې!?`��5���@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@U����ٿ*����@����3@]sqՐ!?�-�n0��@7]��8�ٿ�F����@#O�N��3@8�Vgڐ!?[�˽���@7]��8�ٿ�F����@#O�N��3@8�Vgڐ!?[�˽���@7]��8�ٿ�F����@#O�N��3@8�Vgڐ!?[�˽���@����a�ٿ�3����@S ��u�3@�\Hˊ�!?	:�G��@����a�ٿ�3����@S ��u�3@�\Hˊ�!?	:�G��@����a�ٿ�3����@S ��u�3@�\Hˊ�!?	:�G��@����a�ٿ�3����@S ��u�3@�\Hˊ�!?	:�G��@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@�a�x�ٿ�ȼ�	��@�[Wz�3@iHa���!?��P���@ީ�cٜٿw�����@��8}�3@R}����!?�{����@a�!u͙ٿu)���@(��Sb�3@FͰ/�!?����@a�!u͙ٿu)���@(��Sb�3@FͰ/�!?����@a�!u͙ٿu)���@(��Sb�3@FͰ/�!?����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@����]�ٿ������@�qN��3@:�Q�C�!?�G����@��&e�ٿ���=��@:�����3@�{;�!?�7ͼ(��@��&e�ٿ���=��@:�����3@�{;�!?�7ͼ(��@��&e�ٿ���=��@:�����3@�{;�!?�7ͼ(��@��&e�ٿ���=��@:�����3@�{;�!?�7ͼ(��@��P2�ٿd7�}��@O����3@Eގ3�!?ы�a��@��P2�ٿd7�}��@O����3@Eގ3�!?ы�a��@��P2�ٿd7�}��@O����3@Eގ3�!?ы�a��@y�i�,�ٿ(�5��@qJ��3@��c���!?�P���@Rg��ٿM��L���@��� M�3@E���!?N�U���@Rg��ٿM��L���@��� M�3@E���!?N�U���@~U�(K�ٿ<z���@y�%[S�3@[b]d8�!?������@~U�(K�ٿ<z���@y�%[S�3@[b]d8�!?������@~U�(K�ٿ<z���@y�%[S�3@[b]d8�!?������@~U�(K�ٿ<z���@y�%[S�3@[b]d8�!?������@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@�y
�ٿ�v9��@l��U��3@{B�ݐ!?�N�Ш��@��<��ٿOa�1��@�"f���3@���Ґ!?�SXp���@��<��ٿOa�1��@�"f���3@���Ґ!?�SXp���@��<��ٿOa�1��@�"f���3@���Ґ!?�SXp���@��<��ٿOa�1��@�"f���3@���Ґ!?�SXp���@��<��ٿOa�1��@�"f���3@���Ґ!?�SXp���@Y��a�ٿX��x��@�<����3@�LY�!?w_����@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@�t�m��ٿ$`����@I�'4>�3@���U��!?2�ؔ{��@���c!�ٿK����@R��{��3@�@!��!?�p�ڛ��@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@i?$ܢٿL���@�����3@R��!?�@�)���@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@����B�ٿ'�����@J�;�V�3@v�Zx}�!?�}E����@�ay���ٿr�aI��@�#���3@xp0�l�!?W�r���@�ay���ٿr�aI��@�#���3@xp0�l�!?W�r���@�ay���ٿr�aI��@�#���3@xp0�l�!?W�r���@�t�H�ٿ�}��	��@J����3@�ç&�!?/��	��@�t�H�ٿ�}��	��@J����3@�ç&�!?/��	��@U�fR��ٿ�PS���@���3@b�Nܴ�!?)�&���@�M��ٿlQn���@�Km��3@��Æ��!?�U�A��@�M��ٿlQn���@�Km��3@��Æ��!?�U�A��@|Cޜٿ�x'd���@����1�3@9yE鿐!?�	ΐn��@|Cޜٿ�x'd���@����1�3@9yE鿐!?�	ΐn��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@SЮ|��ٿ�Fb���@Kq�"�3@�[6��!?.�UH��@ U�?�ٿ��@ ��@%����3@��� �!?Y������@S��L�ٿ�m[���@�C�M4�3@�H���!?��<���@S��L�ٿ�m[���@�C�M4�3@�H���!?��<���@S��L�ٿ�m[���@�C�M4�3@�H���!?��<���@ͱ�j�ٿچ̨���@{�f~%�3@w�ug�!?��f�V��@Xκ=��ٿ�d��@�\��3@I���ɐ!?��pk��@Xκ=��ٿ�d��@�\��3@I���ɐ!?��pk��@Xκ=��ٿ�d��@�\��3@I���ɐ!?��pk��@Xκ=��ٿ�d��@�\��3@I���ɐ!?��pk��@Xκ=��ٿ�d��@�\��3@I���ɐ!?��pk��@Y���ٿ�]����@ó�r��3@�y��!?�]ӎ���@Y���ٿ�]����@ó�r��3@�y��!?�]ӎ���@Y���ٿ�]����@ó�r��3@�y��!?�]ӎ���@���̟ٿ�3���@���i�3@�L���!?4�����@��yO��ٿ����@�T�@h�3@)��Đ!?�#����@�B0,˚ٿ�Ȅ���@�S55]�3@K=��ʐ!??j
%o��@�B0,˚ٿ�Ȅ���@�S55]�3@K=��ʐ!??j
%o��@�B0,˚ٿ�Ȅ���@�S55]�3@K=��ʐ!??j
%o��@�B0,˚ٿ�Ȅ���@�S55]�3@K=��ʐ!??j
%o��@:�e���ٿT1�c��@)�#*s�3@J�ħ��!?�\ �@��@:�e���ٿT1�c��@)�#*s�3@J�ħ��!?�\ �@��@:�e���ٿT1�c��@)�#*s�3@J�ħ��!?�\ �@��@����ٿs�6���@��}�3@&�uw,�!?�B��]��@��ꎣٿB����@�B���3@��
~�!?�_� ���@��ꎣٿB����@�B���3@��
~�!?�_� ���@��ꎣٿB����@�B���3@��
~�!?�_� ���@��UƜٿ ݄[���@��v�q�3@����&�!?U�m��@W��֜ٿ�����@��M�*�3@���̐!?���(���@W��֜ٿ�����@��M�*�3@���̐!?���(���@W��֜ٿ�����@��M�*�3@���̐!?���(���@��(v�ٿ�������@���u�3@��S���!?=n>���@��(v�ٿ�������@���u�3@��S���!?=n>���@��(v�ٿ�������@���u�3@��S���!?=n>���@��(v�ٿ�������@���u�3@��S���!?=n>���@��(v�ٿ�������@���u�3@��S���!?=n>���@�ݐ��ٿ���@h����3@���Ȑ!?Z%1����@�ݐ��ٿ���@h����3@���Ȑ!?Z%1����@�ݐ��ٿ���@h����3@���Ȑ!?Z%1����@�ݐ��ٿ���@h����3@���Ȑ!?Z%1����@�ݐ��ٿ���@h����3@���Ȑ!?Z%1����@�}��ٿN�����@���h�3@��(���!?(3ο��@�}��ٿN�����@���h�3@��(���!?(3ο��@�}��ٿN�����@���h�3@��(���!?(3ο��@�}��ٿN�����@���h�3@��(���!?(3ο��@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@�ԟ���ٿ!�6���@�����3@��C|�!?^�����@B�Oo�ٿ^y���@���Hb�3@U�ϫ��!?q?����@R���B�ٿI�G���@�UЕ��3@<�l�x�!?���v��@R���B�ٿI�G���@�UЕ��3@<�l�x�!?���v��@R���B�ٿI�G���@�UЕ��3@<�l�x�!?���v��@�V�Ӝٿ?������@:�J���3@��	��!?fQ6cF��@�V�Ӝٿ?������@:�J���3@��	��!?fQ6cF��@�V�Ӝٿ?������@:�J���3@��	��!?fQ6cF��@�V�Ӝٿ?������@:�J���3@��	��!?fQ6cF��@m�>r��ٿXdr���@�X'���3@�􎢦�!?��&ߏ��@P�>աٿI����@@-`V��3@ D��!?�+����@P�>աٿI����@@-`V��3@ D��!?�+����@P�>աٿI����@@-`V��3@ D��!?�+����@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�ٙ�ٿ\�JJ$��@^!�ID�3@G����!?\���[��@�O6�a�ٿ^l����@/��L�3@N���M�!?��6{��@�O6�a�ٿ^l����@/��L�3@N���M�!?��6{��@�O6�a�ٿ^l����@/��L�3@N���M�!?��6{��@q��$�ٿ���
��@�.���3@�8c�L�!?�7Ν���@q��$�ٿ���
��@�.���3@�8c�L�!?�7Ν���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�@�\��ٿ����J��@���j�3@�`�U��!?�& v���@�Q }�ٿ	������@�V��3@u�ϐ!?�������@�Q }�ٿ	������@�V��3@u�ϐ!?�������@&��ٿ�����@�����3@�H>W��!?%�&���@&��ٿ�����@�����3@�H>W��!?%�&���@B	��x�ٿh��χ�@x����3@�Z�YE�!?w�-`���@B	��x�ٿh��χ�@x����3@�Z�YE�!?w�-`���@�Zi�ٿ�ѽ���@˗D�7�3@����!?��dd��@�Zi�ٿ�ѽ���@˗D�7�3@����!?��dd��@j���ٿ)����@��fG��3@>?�c�!?z�A ���@���>��ٿ��	eL��@�V���3@Iѓyސ!?����a��@���>��ٿ��	eL��@�V���3@Iѓyސ!?����a��@���>��ٿ��	eL��@�V���3@Iѓyސ!?����a��@���>��ٿ��	eL��@�V���3@Iѓyސ!?����a��@�x�ٿ���n��@I9���3@����:�!?�s�5���@�x�ٿ���n��@I9���3@����:�!?�s�5���@�x�ٿ���n��@I9���3@����:�!?�s�5���@�n��ؠٿ��`-(��@w}[���3@ݩ�	�!?W�os��@�n��ؠٿ��`-(��@w}[���3@ݩ�	�!?W�os��@�n��ؠٿ��`-(��@w}[���3@ݩ�	�!?W�os��@BV�Z��ٿK���@�q�A��3@��ky�!?~:V����@�<Y(Şٿ��L���@L/��;�3@��?��!? `Ț3��@�<Y(Şٿ��L���@L/��;�3@��?��!? `Ț3��@�<Y(Şٿ��L���@L/��;�3@��?��!? `Ț3��@�<Y(Şٿ��L���@L/��;�3@��?��!? `Ț3��@�Z��ٿ����w��@܀���3@Ы |�!?�y�h��@�Z��ٿ����w��@܀���3@Ы |�!?�y�h��@�Z��ٿ����w��@܀���3@Ы |�!?�y�h��@�Z��ٿ����w��@܀���3@Ы |�!?�y�h��@�>�-�ٿ���/x��@��a�M�3@tK[�!?q\�O��@�>�-�ٿ���/x��@��a�M�3@tK[�!?q\�O��@�>�-�ٿ���/x��@��a�M�3@tK[�!?q\�O��@ix�L͝ٿ'p�bE��@�f�2�3@[m���!? ����@ix�L͝ٿ'p�bE��@�f�2�3@[m���!? ����@ix�L͝ٿ'p�bE��@�f�2�3@[m���!? ����@�(&�˙ٿ�`s֤��@�G�A�3@,�F|��!?'����@�(&�˙ٿ�`s֤��@�G�A�3@,�F|��!?'����@�(&�˙ٿ�`s֤��@�G�A�3@,�F|��!?'����@�(&�˙ٿ�`s֤��@�G�A�3@,�F|��!?'����@�(&�˙ٿ�`s֤��@�G�A�3@,�F|��!?'����@��Ź�ٿV�lIĈ�@Ԩ����3@][�4��!?6��n�	�@��Ź�ٿV�lIĈ�@Ԩ����3@][�4��!?6��n�	�@p����ٿ�3a���@ f���3@v���*�!?Nę����@�
�ךٿFQ�1}��@����3@����X�!?]�v��@�
�ךٿFQ�1}��@����3@����X�!?]�v��@z5�ٿ��c����@y���7�3@��a��!?n+*�@z5�ٿ��c����@y���7�3@��a��!?n+*�@��3Ԥٿ\�t�B��@h�����3@�Z�!?]�6��@��3Ԥٿ\�t�B��@h�����3@�Z�!?]�6��@��3Ԥٿ\�t�B��@h�����3@�Z�!?]�6��@��3Ԥٿ\�t�B��@h�����3@�Z�!?]�6��@��3Ԥٿ\�t�B��@h�����3@�Z�!?]�6��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@�f͂��ٿ�J3���@1���3@���+��!?�N&��@N���՚ٿ�=%����@?���A�3@-��NQ�!?|*Ji��@N���՚ٿ�=%����@?���A�3@-��NQ�!?|*Ji��@N���՚ٿ�=%����@?���A�3@-��NQ�!?|*Ji��@.�r�ٿXj@���@��7#�3@��B9��!? B��k��@.�r�ٿXj@���@��7#�3@��B9��!? B��k��@.�r�ٿXj@���@��7#�3@��B9��!? B��k��@.�r�ٿXj@���@��7#�3@��B9��!? B��k��@.�r�ٿXj@���@��7#�3@��B9��!? B��k��@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@c���ٿk:�V��@i�z�j�3@ξ��Ӑ!?8��r���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@��kq�ٿ�l.]��@F%L(b�3@��=��!?�8)v���@6?6b
�ٿCc,>P��@@{T��3@����7�!?`+�J��@6?6b
�ٿCc,>P��@@{T��3@����7�!?`+�J��@gI�Ӈ�ٿ��Ȃ��@��ɔ��3@E(�y֐!?������@gI�Ӈ�ٿ��Ȃ��@��ɔ��3@E(�y֐!?������@�b]�
�ٿN'�Db��@e�K�3@o�1�!?th�U}
�@�b]�
�ٿN'�Db��@e�K�3@o�1�!?th�U}
�@�b]�
�ٿN'�Db��@e�K�3@o�1�!?th�U}
�@��V���ٿ��b^���@8���3@?�s��!?�7�%��@��V���ٿ��b^���@8���3@?�s��!?�7�%��@��V���ٿ��b^���@8���3@?�s��!?�7�%��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@7Ž֦�ٿ:�@����@�g7��3@O��!?Am��@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@BI�t�ٿ"�6����@��'���3@��@��!?|���
�@<8��x�ٿ��&��@<ӟ9�3@P���!?�'��@<8��x�ٿ��&��@<ӟ9�3@P���!?�'��@��7 ��ٿ��3z��@��{b!�3@�!*��!?�i�h �@���'�ٿ���!��@q{����3@}Ϻ��!?�=�J��@���'�ٿ���!��@q{����3@}Ϻ��!?�=�J��@V_4���ٿ@�,���@��60�3@h[%��!?���{���@oBPzP�ٿ�ŭ%Æ�@�^�3@c� Ґ!?,S��?��@oBPzP�ٿ�ŭ%Æ�@�^�3@c� Ґ!?,S��?��@oBPzP�ٿ�ŭ%Æ�@�^�3@c� Ґ!?,S��?��@ൻ�ʜٿ�5��͇�@�@���3@��û*�!?�c]����@ൻ�ʜٿ�5��͇�@�@���3@��û*�!?�c]����@ൻ�ʜٿ�5��͇�@�@���3@��û*�!?�c]����@ൻ�ʜٿ�5��͇�@�@���3@��û*�!?�c]����@ൻ�ʜٿ�5��͇�@�@���3@��û*�!?�c]����@t�8�m�ٿ�@4N:��@&��_�3@����ǐ!?�T�ީ��@���_}�ٿ�^����@�d���3@��7r�!?oeZx�@���_}�ٿ�^����@�d���3@��7r�!?oeZx�@���_}�ٿ�^����@�d���3@��7r�!?oeZx�@���_}�ٿ�^����@�d���3@��7r�!?oeZx�@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@��8:p�ٿ������@��9{��3@���O�!?��T	��@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�_��ǡٿ�����@��KW{�3@8��]�!?v6�-���@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@�n/���ٿJ('����@�#e&�3@�!��!?[�9��@(���˟ٿX��@��@���q�3@!�����!?��Z$��@(���˟ٿX��@��@���q�3@!�����!?��Z$��@(���˟ٿX��@��@���q�3@!�����!?��Z$��@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@�fp�P�ٿ�V��W��@m.�� �3@_��6ʐ!?��[����@���)�ٿ�궿3��@e��+�3@�W���!?�BvԠ�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@��q�`�ٿh�W˃�@K�w���3@�>�|�!?f>�4i�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@�2�ٿh��B��@���3@��G�_�!?ssC�@^�@M}>#ޤٿv7Y�|��@H�CKW�3@,�\�:�!?�
�M�4�@M}>#ޤٿv7Y�|��@H�CKW�3@,�\�:�!?�
�M�4�@M}>#ޤٿv7Y�|��@H�CKW�3@,�\�:�!?�
�M�4�@M}>#ޤٿv7Y�|��@H�CKW�3@,�\�:�!?�
�M�4�@��آٿ��cQ���@�#�,�3@a?l敖!?�!����@��آٿ��cQ���@�#�,�3@a?l敖!?�!����@��آٿ��cQ���@�#�,�3@a?l敖!?�!����@��آٿ��cQ���@�#�,�3@a?l敖!?�!����@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@��+:�ٿh�>�+��@���Ba�3@��MÐ!?��ߜ�@�����ٿ������@b�e<7�3@^ѲZ��!?lz)O}��@�����ٿ������@b�e<7�3@^ѲZ��!?lz)O}��@G�zT7�ٿ�fk)��@쟺l�3@��f�>�!?I�Zo�@���K��ٿ��$���@�v&��3@�0���!?r��Nӛ�@�aW')�ٿ'�����@VN��R�3@���(��!?9A=;t��@�aW')�ٿ'�����@VN��R�3@���(��!?9A=;t��@�aW')�ٿ'�����@VN��R�3@���(��!?9A=;t��@�aW')�ٿ'�����@VN��R�3@���(��!?9A=;t��@���,ڦٿ�����@��٦Q�3@c�l5��!?{K����@���,ڦٿ�����@��٦Q�3@c�l5��!?{K����@���,ڦٿ�����@��٦Q�3@c�l5��!?{K����@���,ڦٿ�����@��٦Q�3@c�l5��!?{K����@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@�L��ٿ����1��@���K��3@�`&���!?�k�fb�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@Wa�w)�ٿFq����@W$a��3@J��!?�+��U�@2��%d�ٿ�>H���@<ѡ[��3@���!?^�*G�;�@2��%d�ٿ�>H���@<ѡ[��3@���!?^�*G�;�@2��%d�ٿ�>H���@<ѡ[��3@���!?^�*G�;�@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@�6��ٿZ�7��@��`;��3@B��[��!?��߭H��@0��RE�ٿB��	��@;�&���3@�j �!?!�TA��@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@��o�ٿ.K�~���@������3@�����!?�=��U�@
��Ԛٿ��"}Ԉ�@�<���3@�˳غ�!?�P<4L�@
��Ԛٿ��"}Ԉ�@�<���3@�˳غ�!?�P<4L�@
��Ԛٿ��"}Ԉ�@�<���3@�˳غ�!?�P<4L�@
��Ԛٿ��"}Ԉ�@�<���3@�˳غ�!?�P<4L�@K����ٿ2��@je���3@�����!?��]��a�@K����ٿ2��@je���3@�����!?��]��a�@K����ٿ2��@je���3@�����!?��]��a�@K����ٿ2��@je���3@�����!?��]��a�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@>T���ٿՂ�XS��@��b�3@zR����!?�p��v�@�"�.�ٿG�-lj��@�֮Y��3@u-*�{�!?b�<���@�"�.�ٿG�-lj��@�֮Y��3@u-*�{�!?b�<���@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@�"�ٿ�>����@]�C=e�3@��Ɛ!?�V�29��@W��	��ٿH������@��$3��3@$p�Έ�!?uz���@W��	��ٿH������@��$3��3@$p�Έ�!?uz���@W��	��ٿH������@��$3��3@$p�Έ�!?uz���@W��	��ٿH������@��$3��3@$p�Έ�!?uz���@��[w�ٿS��#���@fL:0�3@qav���!?�,p����@��[w�ٿS��#���@fL:0�3@qav���!?�,p����@��[w�ٿS��#���@fL:0�3@qav���!?�,p����@��[w�ٿS��#���@fL:0�3@qav���!?�,p����@��[w�ٿS��#���@fL:0�3@qav���!?�,p����@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@� �5�ٿ$��옆�@u���3@�'�A��!?���L��@Z��b�ٿ�M9M���@.���H�3@�U����!?-h*��1�@Z��b�ٿ�M9M���@.���H�3@�U����!?-h*��1�@�����ٿ��',}�@�YLb{�3@>T���!?��d���@�����ٿ��',}�@�YLb{�3@>T���!?��d���@�u��2�ٿ����j��@,��(��3@d/�ʐ!?@�L2�T�@�u��2�ٿ����j��@,��(��3@d/�ʐ!?@�L2�T�@�u��2�ٿ����j��@,��(��3@d/�ʐ!?@�L2�T�@O?]��ٿ�./+���@��Ҕ�3@ъ�ِ!?tF!B���@O?]��ٿ�./+���@��Ҕ�3@ъ�ِ!?tF!B���@O?]��ٿ�./+���@��Ҕ�3@ъ�ِ!?tF!B���@O?]��ٿ�./+���@��Ҕ�3@ъ�ِ!?tF!B���@O?]��ٿ�./+���@��Ҕ�3@ъ�ِ!?tF!B���@��b'�ٿ��~˓�@����3@�"�9ސ!?O��۰��@��b'�ٿ��~˓�@����3@�"�9ސ!?O��۰��@���f�ٿ�����@~�Ę7�3@��*G�!?���Ip�@���f�ٿ�����@~�Ę7�3@��*G�!?���Ip�@R�.S>�ٿ�p��@��`�p�3@��&l��!?$iѧ��@�yޛٿ �.��@�Cɦ�3@Q��ߐ!?�%�v��@�yޛٿ �.��@�Cɦ�3@Q��ߐ!?�%�v��@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@)YM4��ٿ�6ލ5��@��� u�3@�]	?�!?��h�4�@���暥ٿ6g��=��@���<��3@��+��!?��z���@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@}_ƍ��ٿ�C�P��@?�8���3@7M(��!?e�UL�D�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@t��V�ٿ���a���@Ƃm4�3@��xT�!?y���.�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@q����ٿD5�0X��@��`��3@�����!?KT�19P�@z���šٿ��jS���@,|��\�3@�1���!?0r��l�@z���šٿ��jS���@,|��\�3@�1���!?0r��l�@��s�ٿ�V�|�@*�b2�3@�99w�!?k��o6�@��s�ٿ�V�|�@*�b2�3@�99w�!?k��o6�@��s�ٿ�V�|�@*�b2�3@�99w�!?k��o6�@��s�ٿ�V�|�@*�b2�3@�99w�!?k��o6�@��s�ٿ�V�|�@*�b2�3@�99w�!?k��o6�@_���ٿ��#o��@���T�3@|u0E}�!?̑���@b���ßٿg*��Ԁ�@Z<�u�3@�N~b��!?l�ah��@b���ßٿg*��Ԁ�@Z<�u�3@�N~b��!?l�ah��@�ihn��ٿg���5��@k�ǐ�3@�2�.��!?��H����@�ihn��ٿg���5��@k�ǐ�3@�2�.��!?��H����@��)�ٿ_?W|�@tmN7G�3@jǢ<��!?SQ�#q�@��)�ٿ_?W|�@tmN7G�3@jǢ<��!?SQ�#q�@O'��ٿ�?V��@�Z���3@�G!?�H&����@O'��ٿ�?V��@�Z���3@�G!?�H&����@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�T�B�ٿ���|�@��#sW�3@�( �<�!?���'G�@�Rˬ2�ٿ;�h���@����t�3@9��O�!?w콍���@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@��y�ؠٿ���'��@��6�� 4@<�́ΐ!?W��^H!�@�l�l�ٿ-L��o��@%�H���3@��ք�!?�*O�~�@�l�l�ٿ-L��o��@%�H���3@��ք�!?�*O�~�@$y�I�ٿ<�aٓ�@'7en��3@�MN_�!?hS����@$y�I�ٿ<�aٓ�@'7en��3@�MN_�!?hS����@$y�I�ٿ<�aٓ�@'7en��3@�MN_�!?hS����@$y�I�ٿ<�aٓ�@'7en��3@�MN_�!?hS����@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�5��ٿL�ܡ��@��^�3@���e �!?%�i%Q��@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�����ٿ7�"��@M���3@�F�|��!?ϧ�^���@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�u܊�ٿ�$��ŕ�@�k���3@	��`͐!?b�>m�@�����ٿ+�J��@��zG�3@�~�W��!?����k�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@���U�ٿ��e��@�����3@�~�oܐ!?k�MeH�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@l���4�ٿ�<u.@��@z`����3@�n�K��!?e۩��C�@9�u��ٿ�g v'��@�*i��3@[��F��!?pr��E��@V^t�ٿ@�:����@��Ă��3@�3��!?�sB}"�@V^t�ٿ@�:����@��Ă��3@�3��!?�sB}"�@V^t�ٿ@�:����@��Ă��3@�3��!?�sB}"�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@�}�/��ٿ�'���@�Z�%�3@��	)�!?-���m�@F���ٿXm��)��@���u��3@f����!?��VA�+�@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��$�ٿ�,�n���@:A�C�3@��K�ϐ!?X�����@��!��ٿ�h�se��@����3@�-{ǐ!?�j��Q�@��!��ٿ�h�se��@����3@�-{ǐ!?�j��Q�@��!��ٿ�h�se��@����3@�-{ǐ!?�j��Q�@'��6ӡٿV�v"}�@_O^Ub�3@�����!?�8̈2��@'��6ӡٿV�v"}�@_O^Ub�3@�����!?�8̈2��@'��6ӡٿV�v"}�@_O^Ub�3@�����!?�8̈2��@'��6ӡٿV�v"}�@_O^Ub�3@�����!?�8̈2��@��>{�ٿ�]�� z�@�zb��3@|�f�!?�+�q{��@��>{�ٿ�]�� z�@�zb��3@|�f�!?�+�q{��@��>{�ٿ�]�� z�@�zb��3@|�f�!?�+�q{��@��>{�ٿ�]�� z�@�zb��3@|�f�!?�+�q{��@��>{�ٿ�]�� z�@�zb��3@|�f�!?�+�q{��@��*~�ٿ,K:t�q�@�o��1�3@�د�!?�{<ـ��@��*~�ٿ,K:t�q�@�o��1�3@�د�!?�{<ـ��@��*~�ٿ,K:t�q�@�o��1�3@�د�!?�{<ـ��@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@��6�c�ٿ]4٘Iv�@���(�3@D�ِ!?����|�@u�<V�ٿc���|�@c��.��3@����!?��8�z�@u�<V�ٿc���|�@c��.��3@����!?��8�z�@u�<V�ٿc���|�@c��.��3@����!?��8�z�@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@��J�ٿU1~����@���K�3@�4R��!?��o�d��@#Mޱ[�ٿ>�-��@������3@%ț�ʐ!?�V�h0�@!S�x$�ٿ���gx��@q�և��3@�z��!?�ѿ=��@��L�ٿei�xr�@Dd��P�3@������!?.]AQ���@��L�ٿei�xr�@Dd��P�3@������!?.]AQ���@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@BՎ�ٿXSV���@U�[R�3@)��Ɛ!?�I$Ms2�@f��6��ٿ����"z�@�-۵�3@3��!?\��+"R�@f��6��ٿ����"z�@�-۵�3@3��!?\��+"R�@f��6��ٿ����"z�@�-۵�3@3��!?\��+"R�@f��6��ٿ����"z�@�-۵�3@3��!?\��+"R�@f��6��ٿ����"z�@�-۵�3@3��!?\��+"R�@
$�ٿ��}�L��@s�!@+�3@v����!?~Յ�`*�@
$�ٿ��}�L��@s�!@+�3@v����!?~Յ�`*�@
$�ٿ��}�L��@s�!@+�3@v����!?~Յ�`*�@
$�ٿ��}�L��@s�!@+�3@v����!?~Յ�`*�@�L/��ٿ6Q:5��@'�d�J�3@�E��l�!?L�+I���@�L/��ٿ6Q:5��@'�d�J�3@�E��l�!?L�+I���@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��}�Ϛٿ��lK��@�����3@D����!?������@��ݭ�ٿ�҂�z�@��@�3@�~���!?C�*iT��@hk��ٿ�p�����@,)���3@�"J��!?d���@hk��ٿ�p�����@,)���3@�"J��!?d���@hk��ٿ�p�����@,)���3@�"J��!?d���@hk��ٿ�p�����@,)���3@�"J��!?d���@hk��ٿ�p�����@,)���3@�"J��!?d���@�-{n�ٿ�P��I��@�:�Q{�3@����!?�u�R��@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@���p�ٿL�0Yd��@�=J��3@�����!?�x�p���@-ֵc�ٿ������@xd�C�3@��Bސ!?&�{G��@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@���U��ٿ�)���@�w�3@cߩ��!?G���Y�@�M��ٿ���x��@t�j&�3@���ڐ!?'���ż�@�M��ٿ���x��@t�j&�3@���ڐ!?'���ż�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��5ý�ٿy&���@x�w��3@�JjS��!?,<I�+�@��N�2�ٿ��">0��@�K���3@:��K�!? ��v�@!�n���ٿ)�5$Ϧ�@�n �3@�&��ϐ!?��6���@!�n���ٿ)�5$Ϧ�@�n �3@�&��ϐ!?��6���@��@ԃ�ٿ��)���@�B���3@Ư����!?�߯lE��@%��$�ٿ$k\?\��@�2(h�3@��+��!?��TOR��@,]�ٿ��^�Έ�@'���3@�N/���!?����:��@����ٿ�c/�2i�@'9�I��3@}�3	��!?;ٹyY0�@����ٿ�c/�2i�@'9�I��3@}�3	��!?;ٹyY0�@�4���ٿ�tE��^�@һP"�3@�H2��!?�������@�	
��ٿ.;
K�u�@�L�pU�3@�މ4�!?�Hxz�,�@O-��ٿ��i;ca�@JZF��3@ɀ�>��!?�0lyB��@O-��ٿ��i;ca�@JZF��3@ɀ�>��!?�0lyB��@O-��ٿ��i;ca�@JZF��3@ɀ�>��!?�0lyB��@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�/��ٿU��@�n�@ό�"��3@
\꣐!?�8�ږ�@�g�p�ٿpI	����@�]�O��3@�F����!?�����z�@�g�p�ٿpI	����@�]�O��3@�F����!?�����z�@�g�p�ٿpI	����@�]�O��3@�F����!?�����z�@Z��(I�ٿ������@r����3@r�i��!?����8��@Z��(I�ٿ������@r����3@r�i��!?����8��@Z��(I�ٿ������@r����3@r�i��!?����8��@��~P�ٿ��M`�@Un
��3@��Ð!???Ɓp�@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@k*���ٿ �d��b�@B��^-�3@^X�]Ր!?֘�����@Р"#t�ٿ0������@`�|k�3@	���!?u�i�.��@Р"#t�ٿ0������@`�|k�3@	���!?u�i�.��@Р"#t�ٿ0������@`�|k�3@	���!?u�i�.��@Р"#t�ٿ0������@`�|k�3@	���!?u�i�.��@�����ٿ�Bt��@�"lV�3@��U[��!?S��ˠ�@�����ٿ�Bt��@�"lV�3@��U[��!?S��ˠ�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@پ���ٿ� ����@�&�i�3@a��埐!?�hɖl\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@]p�ٿ��	1���@R�HQ�3@Ԕ�!?	[M�\�@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@�uG*i�ٿN�H���@��AR�3@&rÐ!?^R�E��@D�2���ٿ�|#\��@gr����3@-�e�Ґ!?���@��@D�2���ٿ�|#\��@gr����3@-�e�Ґ!?���@��@D�2���ٿ�|#\��@gr����3@-�e�Ґ!?���@��@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@�.�=�ٿ�)���@GL6l�3@<�$��!?�-,W���@Mgߚٿ��tﻩ�@
�Ki��3@K��z�!?(�H�C�@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@���L�ٿ�����@�(���3@Pw(~��!?D)�j��@]{AGz�ٿ,��sƊ�@�͛��3@����!?�w"(�@]{AGz�ٿ,��sƊ�@�͛��3@����!?�w"(�@]{AGz�ٿ,��sƊ�@�͛��3@����!?�w"(�@]{AGz�ٿ,��sƊ�@�͛��3@����!?�w"(�@`<�b�ٿ]uV��@Ǯ���3@ x҄Ԑ!?K)�}P�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@8k�p �ٿJ:۹4��@�3h���3@?�Gּ�!?��1�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@��S��ٿ�V ���@^ջ�x�3@�.�"��!?2M�G�e�@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@8,�o��ٿ�/
�q��@�$q��3@�#�.��!?ܛ&%��@)Jw��ٿ_-�8���@{_��3@���T�!?��8�=c�@w�\��ٿ�n���@�J7R�3@��Vx�!?�m,)���@jP��d�ٿ������@b��Y��3@�"o=a�!?9}��@jP��d�ٿ������@b��Y��3@�"o=a�!?9}��@jP��d�ٿ������@b��Y��3@�"o=a�!?9}��@����ӟٿg��ٕ�@\SՌ�3@B[ᨫ�!?�sXD�@����ӟٿg��ٕ�@\SՌ�3@B[ᨫ�!?�sXD�@����ӟٿg��ٕ�@\SՌ�3@B[ᨫ�!?�sXD�@!+�w��ٿ�)�D��@o�D��3@G�А!?���@!+�w��ٿ�)�D��@o�D��3@G�А!?���@!+�w��ٿ�)�D��@o�D��3@G�А!?���@!+�w��ٿ�)�D��@o�D��3@G�А!?���@!+�w��ٿ�)�D��@o�D��3@G�А!?���@!+�w��ٿ�)�D��@o�D��3@G�А!?���@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@*��ğٿ��F����@�-�9O�3@Xs'��!?b{� `��@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�?N�ٿ\�[���@2��U+�3@��=Px�!?�{�ܗ^�@�.ڧ<�ٿ��G+��@Yk1��3@�=��!?��/eF�@�.ڧ<�ٿ��G+��@Yk1��3@�=��!?��/eF�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@2�y��ٿ���bB��@.l����3@��ل&�!?�ZWt!
�@��Ӝx�ٿ��-8��@���w�3@X�5�]�!?d��a��@2\�x�ٿ��Լ4��@�"&n�3@lk�*K�!?�T����@2\�x�ٿ��Լ4��@�"&n�3@lk�*K�!?�T����@2\�x�ٿ��Լ4��@�"&n�3@lk�*K�!?�T����@�G�I͠ٿ�ڲ�R��@kQ��3@�Zx���!?��m�Z�@�G�I͠ٿ�ڲ�R��@kQ��3@�Zx���!?��m�Z�@�FҮ�ٿ�C����@EJ�A{�3@^�:��!?t�g}��@;\;w��ٿ�I�oL��@ ���3@���.��!?�I6��z�@;\;w��ٿ�I�oL��@ ���3@���.��!?�I6��z�@;\;w��ٿ�I�oL��@ ���3@���.��!?�I6��z�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@q���ٿ4:�Z���@ ��U<�3@��>���!?m�c̎�@2%�~�ٿ���xc�@}<���3@l�6XƐ!?vH�L�@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@�g�8�ٿc��p�x�@	J��a�3@����3�!?�����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@*)���ٿ�膵���@��U��3@�G�� �!?�%]����@��ד�ٿ����@!�WQ�3@}#���!?�9��B�@��ד�ٿ����@!�WQ�3@}#���!?�9��B�@��ד�ٿ����@!�WQ�3@}#���!?�9��B�@��ד�ٿ����@!�WQ�3@}#���!?�9��B�@n���ٿ2z�����@�vK���3@�:H��!?Ѥp
��@n���ٿ2z�����@�vK���3@�:H��!?Ѥp
��@n���ٿ2z�����@�vK���3@�:H��!?Ѥp
��@n���ٿ2z�����@�vK���3@�:H��!?Ѥp
��@�ϵ��ٿoTn�@�@Efc,��3@e�˙�!?\�Ł~�@�ϵ��ٿoTn�@�@Efc,��3@e�˙�!?\�Ł~�@�ϵ��ٿoTn�@�@Efc,��3@e�˙�!?\�Ł~�@�ϵ��ٿoTn�@�@Efc,��3@e�˙�!?\�Ł~�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@�[kaƜٿ;8u�X3�@@�K��3@tu�ސ!?�ݓ��@�@/�3�ٿ'��5�M�@�V\��3@����!?Oe���@/�3�ٿ'��5�M�@�V\��3@����!?Oe���@�l��L�ٿ�,KwS�@�]��P�3@�W����!?�Laޭ�@���Ġ�ٿ��G�=�@�!c���3@XJ@�v�!?���/�@���Ġ�ٿ��G�=�@�!c���3@XJ@�v�!?���/�@���Ġ�ٿ��G�=�@�!c���3@XJ@�v�!?���/�@��͚ٿ�oD!?�@������3@On�h��!?|+Խ��@��͚ٿ�oD!?�@������3@On�h��!?|+Խ��@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@�D/��ٿ��~��@�J�n�3@1&;�ِ!?Y|���@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@ �v���ٿI,�S���@ ��M�3@��	�ߐ!?	�֧c��@����(�ٿ�6H��@�W꺣�3@�~�0�!?�t��b�@K#�h��ٿ�H�>��@��U~n�3@��g �!?͙��:�@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@P�c�3�ٿ6��F�@4Z�3@�vI9�!?���e^��@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@yaM��ٿ#`�B�:�@ uZ1M�3@���lÐ!?��d;���@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@�HBZ�ٿFL ��#�@3T)���3@='	ΐ!?�.�=�@옶��ٿ��`���@��xf�3@���cȐ!?���JZ��@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@�I��#�ٿ�3t���@��^':�3@/܋��!?���Cb�@>���ٿ����_�@u��ǳ�3@(N���!?���HYp�@>���ٿ����_�@u��ǳ�3@(N���!?���HYp�@>���ٿ����_�@u��ǳ�3@(N���!?���HYp�@>���ٿ����_�@u��ǳ�3@(N���!?���HYp�@>���ٿ����_�@u��ǳ�3@(N���!?���HYp�@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@��c��ٿ��w���@�w��3@�P�!?ը!dw��@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@Zo[�ܢٿw(�1���@��,��3@ۨa� �!?�������@�ؕ˖�ٿ7��[`�@�����3@ȧH�!?�<����@�=���ٿ��;EeX�@jE��,�3@7�jŐ!?e��^��@�=���ٿ��;EeX�@jE��,�3@7�jŐ!?e��^��@�=���ٿ��;EeX�@jE��,�3@7�jŐ!?e��^��@�=���ٿ��;EeX�@jE��,�3@7�jŐ!?e��^��@�ʈm�ٿC��`��@�ʼ��3@k�Y��!?��  �r�@�ʈm�ٿC��`��@�ʼ��3@k�Y��!?��  �r�@�ʈm�ٿC��`��@�ʼ��3@k�Y��!?��  �r�@�ʈm�ٿC��`��@�ʼ��3@k�Y��!?��  �r�@�ʈm�ٿC��`��@�ʼ��3@k�Y��!?��  �r�@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@��pMܢٿ�#jD��@f����3@�� ��!?=q {9��@�����ٿ�����@��yM��3@���M�!?�����&�@�����ٿ�����@��yM��3@���M�!?�����&�@�ළ�ٿ�R�+ J�@��|��3@��,5�!?u	r�H��@�ළ�ٿ�R�+ J�@��|��3@��,5�!?u	r�H��@�ළ�ٿ�R�+ J�@��|��3@��,5�!?u	r�H��@�kH��ٿ*
����@���S�3@�Ux4�!?M�
E�f�@����d�ٿ�gvL�@!P�-a�3@4�O���!?�݂b�!�@����d�ٿ�gvL�@!P�-a�3@4�O���!?�݂b�!�@����d�ٿ�gvL�@!P�-a�3@4�O���!?�݂b�!�@����d�ٿ�gvL�@!P�-a�3@4�O���!?�݂b�!�@��R���ٿ�Il�C�@e��k�3@'�k(O�!?���9��@��R���ٿ�Il�C�@e��k�3@'�k(O�!?���9��@� N�ٿ��+~�:�@�2����3@�I���!?�/0���@� N�ٿ��+~�:�@�2����3@�I���!?�/0���@���p�ٿ,�Y�m�@!�	��3@�9���!?�<$���@X�ߤ�ٿ��5)�5�@�"���3@~�G�ʐ!?}�̐��@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@��.��ٿ�����@��n��3@�Wz)��!?�S��>]�@%&C\�ٿ���ݤt�@s�Q���3@#nM䁐!?����٪�@%&C\�ٿ���ݤt�@s�Q���3@#nM䁐!?����٪�@%&C\�ٿ���ݤt�@s�Q���3@#nM䁐!?����٪�@%&C\�ٿ���ݤt�@s�Q���3@#nM䁐!?����٪�@���_�ٿ2nw�C��@����3@
UV-�!?��Uܧ��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@���01�ٿpV2:@�@�LϽ�3@�Z��i�!?X��xH��@Nj'BN�ٿY�lvg�@��Z�M�3@㸼�n�!?$�]���@Nj'BN�ٿY�lvg�@��Z�M�3@㸼�n�!?$�]���@����ٿP.���@�D0t�3@�Y�(��!?���
���@����ٿP.���@�D0t�3@�Y�(��!?���
���@����ٿP.���@�D0t�3@�Y�(��!?���
���@����ٿP.���@�D0t�3@�Y�(��!?���
���@%Q+�ٿ��i����@n��h��3@Kw(<�!?��ѩ&�@%Q+�ٿ��i����@n��h��3@Kw(<�!?��ѩ&�@ܟ��ٿ.6�z|�@q!��4@��J8��!?��r�&5�@ܟ��ٿ.6�z|�@q!��4@��J8��!?��r�&5�@��!��ٿ�`�P��@nmz�4@�1���!?y�ڌ���@��!��ٿ�`�P��@nmz�4@�1���!?y�ڌ���@C��5X�ٿ!��{w��@�I��3@j�Տ��!?�|cGz@�@?q��ٿ�g6��@�zu_�3@�Ssﳐ!?�)�w��@?q��ٿ�g6��@�zu_�3@�Ssﳐ!?�)�w��@?q��ٿ�g6��@�zu_�3@�Ssﳐ!?�)�w��@?q��ٿ�g6��@�zu_�3@�Ssﳐ!?�)�w��@?q��ٿ�g6��@�zu_�3@�Ssﳐ!?�)�w��@�ܐ�ٿ���]_�@��]|�3@��Ґ!?qP��{�@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@���}	�ٿ~�D`~�@F�OJ�3@]	�z{�!?E���+��@b����ٿ��O����@�[^,�3@�ś��!?��<%d��@b����ٿ��O����@�[^,�3@�ś��!?��<%d��@b����ٿ��O����@�[^,�3@�ś��!?��<%d��@b����ٿ��O����@�[^,�3@�ś��!?��<%d��@b����ٿ��O����@�[^,�3@�ś��!?��<%d��@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@�֢3�ٿ��G�|�@0D�i��3@ѐ�f��!?p��[?z�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@���5��ٿ2&�I���@pg��3@�~�y�!?��_a̹�@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@!�S�,�ٿE��I��@fC��(�3@���P�!?-d��v��@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@/����ٿ�}+>���@�t�)�3@�=�ސ!?�j�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@0}��۠ٿ�-V�@Vg%�Q�3@��s��!?����J�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@�i��W�ٿ���S<�@6�_�3@�Un]ܐ!?p�O�9�@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@)3Gi��ٿ�m�����@3H�$�3@5}��Ӑ!?S-����@�	�+��ٿ�d{g��@��2-�3@a���!?�!��G9�@�	�+��ٿ�d{g��@��2-�3@a���!?�!��G9�@Ɯ)��ٿ�:pl���@n�tf��3@lm��!?}�^e�@�MvܟٿJi�*�[�@��!��3@��Q���!?KZ,
J�@�[���ٿ4c�[Ą�@��ۥ�3@m�hz��!?���Ƞ7�@�W;Ś�ٿE���/y�@dK���3@[��ߐ!?�(�!�u�@�e	�ٿ��v��$�@~����3@O�<�!?��y�2��@�e	�ٿ��v��$�@~����3@O�<�!?��y�2��@�l�c>�ٿV[*�ɓ�@znDN��3@��)ѭ�!?�|K�@�l�c>�ٿV[*�ɓ�@znDN��3@��)ѭ�!?�|K�@��֑N�ٿ��"�r��@R����3@�p�!?��
���@��֑N�ٿ��"�r��@R����3@�p�!?��
���@��֑N�ٿ��"�r��@R����3@�p�!?��
���@�"Y>�ٿ��0yd��@qb��3@V���!?�R�R!�@�"Y>�ٿ��0yd��@qb��3@V���!?�R�R!�@]_z���ٿ e�L��@�8��3@�Q,ِ!?��Q���@]_z���ٿ e�L��@�8��3@�Q,ِ!?��Q���@LJ)��ٿ�h���%�@AS���4@	0����!?pڭ�%��@�� �ٿށE��@EB)���3@��M�!?5�s��o�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@O�m�W�ٿ�O�����@�0&�(�3@He]��!?���ԷZ�@�1��8�ٿ ZY�z��@k����3@3|�D��!?I-�j��@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@2���ٿ�7(���@p�(���3@�m!��!?^��5�	�@u=��ٿǕ�}o�@�4@%�3@������!?�_"��@u=��ٿǕ�}o�@�4@%�3@������!?�_"��@u=��ٿǕ�}o�@�4@%�3@������!?�_"��@^]eem�ٿ�������@&'��3@);r��!?*��`���@�A�P=�ٿ��Ucx�@h�5k-�3@̈́���!?�uƫ��@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��7$��ٿ ��X7�@����3@�&Μ!?���Su�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@��ٿ��</�@&8��L�3@���>�!?�%�}�@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@3X��ٿ�s:>{U�@�l��S�3@�hDݐ!?�t�Q���@����ٿ�������@��l���3@�׿��!?[U	��@����ٿ�������@��l���3@�׿��!?[U	��@����ٿ�������@��l���3@�׿��!?[U	��@����ٿ�������@��l���3@�׿��!?[U	��@����ٿ�������@��l���3@�׿��!?[U	��@Hrϧٿ16w�G��@�����3@r��ϐ!?"ҡ"�@Hrϧٿ16w�G��@�����3@r��ϐ!?"ҡ"�@Hrϧٿ16w�G��@�����3@r��ϐ!?"ҡ"�@q���%�ٿiQsE�@��(���3@6-=a��!?M���]�@q���%�ٿiQsE�@��(���3@6-=a��!?M���]�@q���%�ٿiQsE�@��(���3@6-=a��!?M���]�@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@��P�ٿ˼��Z��@��ю�3@��Պא!??��>]��@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@"��ŝٿ'��c��@O�L��3@���!?�D�Ue�@ b}�7�ٿ��+'jp�@L�ފ�3@��ȭ�!?�E�Kz�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@��W���ٿ�P�u�@�'ez�3@e�ΐ!?�A�n�@~��Kٿ�7J62�@ !?�3@�W�̐!?����@~��Kٿ�7J62�@ !?�3@�W�̐!?����@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@4��S��ٿK{�Z6�@I="���3@R0�Y��!?�ǦJ_w�@����ٿӾ��F�@N�Eeh�3@�(O�!?8J��x��@����ٿӾ��F�@N�Eeh�3@�(O�!?8J��x��@����ٿӾ��F�@N�Eeh�3@�(O�!?8J��x��@����ٿӾ��F�@N�Eeh�3@�(O�!?8J��x��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@p��gJ�ٿ���j	�@w�v;��3@�	�\ϐ!?��A=��@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@7۵\�ٿ�����@*�}0��3@��˧�!?H:�����@g����ٿ1�|?5�@¼A&��3@Z߲�Ր!?�'G$��@g����ٿ1�|?5�@¼A&��3@Z߲�Ր!?�'G$��@����i�ٿV[�	�F�@i��W��3@��Ԑ!?Ql1*
�@����i�ٿV[�	�F�@i��W��3@��Ԑ!?Ql1*
�@����i�ٿV[�	�F�@i��W��3@��Ԑ!?Ql1*
�@�ɶ���ٿ�j/d�h�@�e�O�3@�=��!?���jO�@�2�ٿ$V�%��@M�y+r�3@� �^�!?����{V�@�2�ٿ$V�%��@M�y+r�3@� �^�!?����{V�@�'S֟ٿ���b��@�;h͓�3@�P䔐!?��u��@�'S֟ٿ���b��@�;h͓�3@�P䔐!?��u��@�'S֟ٿ���b��@�;h͓�3@�P䔐!?��u��@����ٿ��GI�@^��Y��3@f	��ѐ!?�@B[��@����ٿ��GI�@^��Y��3@f	��ѐ!?�@B[��@����ٿ��GI�@^��Y��3@f	��ѐ!?�@B[��@ݏ@)�ٿcX�K�2�@�h�e�3@[�3HĐ!?Ð����@e�AS�ٿ�9QvR�@,k��U�3@ ���!?��\���@e�AS�ٿ�9QvR�@,k��U�3@ ���!?��\���@e�AS�ٿ�9QvR�@,k��U�3@ ���!?��\���@e�AS�ٿ�9QvR�@,k��U�3@ ���!?��\���@.�Y�U�ٿk�]�@+zfg��3@�͚P��!?є�J���@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@�d˯Z�ٿv����d�@��#p�3@3���!?Q]�Q~�@���n�ٿ-����@&����3@�HĽϐ!?=��C��@���n�ٿ-����@&����3@�HĽϐ!?=��C��@�z(��ٿ�&E���@���)��3@�ϐ!?�<͞��@e�G��ٿ�@M�0~�@:�(u��3@����!?�R�Y1�@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@eɭg�ٿ�o=��x�@"�H���3@�ꐈ��!?��Z��@ȫ����ٿ�m��I�@�SI��3@T��!?�Γ(��@ȫ����ٿ�m��I�@�SI��3@T��!?�Γ(��@ȫ����ٿ�m��I�@�SI��3@T��!?�Γ(��@l����ٿ������@tv;�3@C,͐!?5R]/�@��N_�ٿ^��1�@Ց^\�3@�_��ϐ!?A��w:-�@��N_�ٿ^��1�@Ց^\�3@�_��ϐ!?A��w:-�@��N_�ٿ^��1�@Ց^\�3@�_��ϐ!?A��w:-�@��N_�ٿ^��1�@Ց^\�3@�_��ϐ!?A��w:-�@u�@e�ٿ�{�A8�@����3@Ϻ�5��!?�A�,3��@u�@e�ٿ�{�A8�@����3@Ϻ�5��!?�A�,3��@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�N>e�ٿ&L�'�N�@3�0���3@/�?Z��!?F*�����@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�uU���ٿ�L�!J�@�Z����3@��(��!?Eh7*�u�@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�o,t�ٿ������@%]F��3@������!?ao�y��@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�H�)�ٿ�|����@������3@A�X���!?��1��>�@�SX�M�ٿt��2���@�}����3@`^R<ې!?��]qu�@�SX�M�ٿt��2���@�}����3@`^R<ې!?��]qu�@�3����ٿ{S��m�@B~z���3@1�^ε�!?�[�k��@�3����ٿ{S��m�@B~z���3@1�^ε�!?�[�k��@�3����ٿ{S��m�@B~z���3@1�^ε�!?�[�k��@�3����ٿ{S��m�@B~z���3@1�^ε�!?�[�k��@à��ٿ�VE���@�RW��3@q?]���!?� ��9�@à��ٿ�VE���@�RW��3@q?]���!?� ��9�@F��ب�ٿ1w�a��@�^�V!�3@F^�0��!?�F,5�@F��ب�ٿ1w�a��@�^�V!�3@F^�0��!?�F,5�@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@.�L��ٿQ�V�X�@OC2� �3@碟��!?�����@�^�"��ٿ�GF����@���Y��3@��PH��!?I蜓��@�>��ٿ�6"��%�@9c�=�3@C�QM��!?���YD]�@�>��ٿ�6"��%�@9c�=�3@C�QM��!?���YD]�@�>��ٿ�6"��%�@9c�=�3@C�QM��!?���YD]�@���KR�ٿ�k���,�@��i�3@��u΄�!?�,{n h�@.��oh�ٿ)W'0
�@J2��}�3@��e�!?�I�8�,�@غ��ٿ`W�'e�@�U�M�3@:a��t�!?�B��x�@غ��ٿ`W�'e�@�U�M�3@:a��t�!?�B��x�@غ��ٿ`W�'e�@�U�M�3@:a��t�!?�B��x�@غ��ٿ`W�'e�@�U�M�3@:a��t�!?�B��x�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@���ٿ �F���@�2f��3@i:擪�!?@�n$�N�@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@�����ٿ�=���@=����3@寒cҐ!?"_P��@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@���ٿNz*ƻ�@����3@��4R��!?( &Nʚ�@ �fp֡ٿU@�5�r�@�*�h��3@�ΦĐ!?�:i@4k�@ �fp֡ٿU@�5�r�@�*�h��3@�ΦĐ!?�:i@4k�@��S�ڣٿ Vhf7��@�����3@����!?ͮs����@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@��<�W�ٿz��Gxm�@����1�3@�ݨU�!?��	���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@dO��:�ٿ�x����@kuki��3@��5=֐!?��%D���@'rhx�ٿ(��D��@,�dJ)�3@6��!?wbol&�@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@��97��ٿ���B�@�����3@Ҵ�$�!?�t����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@;�j�ٿZ�;�fI�@�t���3@��K�'�!?����@��]�ٿ����`�@�[j��3@�:i�4�!?�>��=�@f�AR�ٿ%���ۅ�@4�����3@i�}�!?�'9��@�˥��ٿ��Kn���@�`���3@��,Ŵ�!?j�94�J�@�˥��ٿ��Kn���@�`���3@��,Ŵ�!?j�94�J�@�˥��ٿ��Kn���@�`���3@��,Ŵ�!?j�94�J�@�˥��ٿ��Kn���@�`���3@��,Ŵ�!?j�94�J�@�˥��ٿ��Kn���@�`���3@��,Ŵ�!?j�94�J�@>����ٿ���z@�@�A��3@��CҐ!?s����@>����ٿ���z@�@�A��3@��CҐ!?s����@>����ٿ���z@�@�A��3@��CҐ!?s����@�y���ٿs�!![~�@�ڢ���3@E-����!?�;�9�y�@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�y�!�ٿ�3�6_�@��>H�3@B��:��!?�Έl��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@�9虧�ٿ�,u@��@.�y7�3@�@ЯҐ!?���JT��@��w���ٿ}=yYV��@VZ<\H�3@P�d���!?h�at��@��͡ٿ\�"l!��@ᠬǸ�3@*�A�f�!?��@���@��͡ٿ\�"l!��@ᠬǸ�3@*�A�f�!?��@���@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@K^�S�ٿ"n�R���@}�.��3@��:H�!?��^�z�@nz��ٿW��'���@��SU��3@���1�!? tr��@nz��ٿW��'���@��SU��3@���1�!? tr��@nz��ٿW��'���@��SU��3@���1�!? tr��@nz��ٿW��'���@��SU��3@���1�!? tr��@nz��ٿW��'���@��SU��3@���1�!? tr��@H�v�ϟٿ+$�T1�@<;����3@~��P�!?�7����@H�v�ϟٿ+$�T1�@<;����3@~��P�!?�7����@H�v�ϟٿ+$�T1�@<;����3@~��P�!?�7����@H�v�ϟٿ+$�T1�@<;����3@~��P�!?�7����@ܶ	{��ٿ��`���@Sc�9�3@[���v�!?�;�� �@ܶ	{��ٿ��`���@Sc�9�3@[���v�!?�;�� �@�tE�N�ٿ�
�����@*�3Ia�3@1��q�!?Oi0
���@�tE�N�ٿ�
�����@*�3Ia�3@1��q�!?Oi0
���@�tE�N�ٿ�
�����@*�3Ia�3@1��q�!?Oi0
���@��KŜٿ�Yr6:Q�@���X��3@˓�"Ԑ!?�k�~��@��KŜٿ�Yr6:Q�@���X��3@˓�"Ԑ!?�k�~��@��KŜٿ�Yr6:Q�@���X��3@˓�"Ԑ!?�k�~��@��KŜٿ�Yr6:Q�@���X��3@˓�"Ԑ!?�k�~��@��KŜٿ�Yr6:Q�@���X��3@˓�"Ԑ!?�k�~��@�+T��ٿ��)f��@��)74@�e=ϐ!?]�z]T�@�+T��ٿ��)f��@��)74@�e=ϐ!?]�z]T�@�+T��ٿ��)f��@��)74@�e=ϐ!?]�z]T�@�+T��ٿ��)f��@��)74@�e=ϐ!?]�z]T�@�+T��ٿ��)f��@��)74@�e=ϐ!?]�z]T�@\�M�ߕٿ�wlYQ��@�G&b��3@�W��!?�Å+���@jڪ�ٿ�	eq�@1Cj���3@�����!?��U���@�,+T�ٿ���v�@f�8�l�3@x�M� �!?��S99�@�,+T�ٿ���v�@f�8�l�3@x�M� �!?��S99�@�,+T�ٿ���v�@f�8�l�3@x�M� �!?��S99�@�h2��ٿ��$vtz�@�5P�H�3@��D���!?DG&�I��@�h2��ٿ��$vtz�@�5P�H�3@��D���!?DG&�I��@�臩:�ٿ]�q-��@��7��3@4�T�!? ɫ'��@�臩:�ٿ]�q-��@��7��3@4�T�!? ɫ'��@�臩:�ٿ]�q-��@��7��3@4�T�!? ɫ'��@�臩:�ٿ]�q-��@��7��3@4�T�!? ɫ'��@4	ӓM�ٿ�����@�+��,�3@V����!?x�f�<��@4	ӓM�ٿ�����@�+��,�3@V����!?x�f�<��@4	ӓM�ٿ�����@�+��,�3@V����!?x�f�<��@4	ӓM�ٿ�����@�+��,�3@V����!?x�f�<��@���K@�ٿ�Z^���@nr����3@�S0WĐ!?����p�@���K@�ٿ�Z^���@nr����3@�S0WĐ!?����p�@���K@�ٿ�Z^���@nr����3@�S0WĐ!?����p�@���K@�ٿ�Z^���@nr����3@�S0WĐ!?����p�@�࡟�ٿ�OU��@�.���3@�ܼ���!?���K��@�࡟�ٿ�OU��@�.���3@�ܼ���!?���K��@�࡟�ٿ�OU��@�.���3@�ܼ���!?���K��@ ���~�ٿ/�qw�f�@�&I��3@��$F��!?��a(�@ ���~�ٿ/�qw�f�@�&I��3@��$F��!?��a(�@ ���~�ٿ/�qw�f�@�&I��3@��$F��!?��a(�@ ���~�ٿ/�qw�f�@�&I��3@��$F��!?��a(�@ ���~�ٿ/�qw�f�@�&I��3@��$F��!?��a(�@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@@p^'1�ٿ�YO*��@�	�?n�3@>��!?f�}�w��@�r,�ٿ�/�b��@�\���3@M�����!?���� �@J��k��ٿ��06!�@n��s��3@1Ov,�!?��ȱ��@s�&��ٿ�~�@�_�@t*����3@.-]ܝ�!?�l�r�8�@s�&��ٿ�~�@�_�@t*����3@.-]ܝ�!?�l�r�8�@^Q�(�ٿ��˱q��@�*U��3@�a��̐!?@��P!��@^Q�(�ٿ��˱q��@�*U��3@�a��̐!?@��P!��@9.{�ٿ`�����@��	~�3@�9]�k�!?D4չ+�@9.{�ٿ`�����@��	~�3@�9]�k�!?D4չ+�@9.{�ٿ`�����@��	~�3@�9]�k�!?D4չ+�@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@���M�ٿ�/�:�@.ѧ8�3@+���q�!?+������@��8��ٿ�jХ�8�@ �0b��3@�4�J�!?0�hMP�@��8��ٿ�jХ�8�@ �0b��3@�4�J�!?0�hMP�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@x L��ٿYK�U�@~"d3��3@��%7\�!?B�J�Ĉ�@�F���ٿ�'���h�@����3@)�[Z��!?������@�F���ٿ�'���h�@����3@)�[Z��!?������@�F���ٿ�'���h�@����3@)�[Z��!?������@�F���ٿ�'���h�@����3@)�[Z��!?������@�F���ٿ�'���h�@����3@)�[Z��!?������@�F���ٿ�'���h�@����3@)�[Z��!?������@6�w�ٿ�+��g��@������3@�%!?}�����@6�w�ٿ�+��g��@������3@�%!?}�����@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@DJ*F�ٿ!�����@�(�X�3@X&�I��!?n��&���@�'�Y۩ٿ��=�/�@eN��,�3@�z9U��!?�$S�H�@�'�Y۩ٿ��=�/�@eN��,�3@�z9U��!?�$S�H�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@FhA콣ٿɏ�K{�@�˹ٟ�3@Yї���!?��/f�h�@�R���ٿ��*�b��@z��@��3@��-R��!?_q����@�R���ٿ��*�b��@z��@��3@��-R��!?_q����@�R���ٿ��*�b��@z��@��3@��-R��!?_q����@�R���ٿ��*�b��@z��@��3@��-R��!?_q����@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@����%�ٿ��r\��@{��[��3@۰$nא!?a5Y�$�@<t􎱥ٿZT����@*�ע��3@l#�ɐ!?��&�@<t􎱥ٿZT����@*�ע��3@l#�ɐ!?��&�@<t􎱥ٿZT����@*�ע��3@l#�ɐ!?��&�@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@�s��ٿ=�p`t�@3�0��3@�B8��!?q�R��@<f'�w�ٿ�,���Q�@!����3@y+�酐!?)>&(��@G}�b��ٿ���3W�@�q6#c�3@�1@��!?]E�߾�@G}�b��ٿ���3W�@�q6#c�3@�1@��!?]E�߾�@G}�b��ٿ���3W�@�q6#c�3@�1@��!?]E�߾�@G}�b��ٿ���3W�@�q6#c�3@�1@��!?]E�߾�@G}�b��ٿ���3W�@�q6#c�3@�1@��!?]E�߾�@�sB��ٿ��ι!��@�*I��3@�R%�!?�l0*�@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@~�ᶝٿD	*%G��@sy�߹�3@�&�]��!?�6���@� �j�ٿteE����@�E"��3@������!?�g�=���@w0���ٿ�W�u`�@��I��3@�c1B�!?b�N��@w0���ٿ�W�u`�@��I��3@�c1B�!?b�N��@w0���ٿ�W�u`�@��I��3@�c1B�!?b�N��@��=/��ٿ2�9|>�@��s�r�3@�&vq	�!?�y�����@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@��JɜٿV�����@ ���\�3@�Ƈ���!?x��2��@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@`?=Ťٿ������@��2��3@`DBڐ!?ܞa���@7�|�A�ٿ,�NŤ!�@�T���3@aU��!?[�P4��@7�|�A�ٿ,�NŤ!�@�T���3@aU��!?[�P4��@7�|�A�ٿ,�NŤ!�@�T���3@aU��!?[�P4��@7�|�A�ٿ,�NŤ!�@�T���3@aU��!?[�P4��@7�|�A�ٿ,�NŤ!�@�T���3@aU��!?[�P4��@�3�&�ٿ�Y�\>��@f]�v��3@�e�ݐ!?�-��%o�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@� �Ҡٿ�7����@B�k���3@�����!?��҆�@��7I�ٿx{;�Ӓ�@�_v�]�3@~�)�!?��h��@��7I�ٿx{;�Ӓ�@�_v�]�3@~�)�!?��h��@��7I�ٿx{;�Ӓ�@�_v�]�3@~�)�!?��h��@��7I�ٿx{;�Ӓ�@�_v�]�3@~�)�!?��h��@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@���סٿ�����@YL�a�3@�v���!?!���@�I���ٿE�_?���@-�G��3@Q��0��!?�dLl�@�I���ٿE�_?���@-�G��3@Q��0��!?�dLl�@�I���ٿE�_?���@-�G��3@Q��0��!?�dLl�@�I���ٿE�_?���@-�G��3@Q��0��!?�dLl�@�VU'�ٿY���'�@[�v��3@�|�;ܐ!?t0B.�B�@CN:�}�ٿ��u�5��@+o��3@�ݯVo�!?�}���@CN:�}�ٿ��u�5��@+o��3@�ݯVo�!?�}���@CN:�}�ٿ��u�5��@+o��3@�ݯVo�!?�}���@Qf��ڜٿ��h�ҿ�@A���z�3@i�وz�!?E�o�>�@Qf��ڜٿ��h�ҿ�@A���z�3@i�وz�!?E�o�>�@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@�)��ٿ���c�@\T4N2�3@�,�Oڐ!?3��"/��@� b!עٿ�#��\��@��)M�3@Q}J£�!?$��p��@A�r{��ٿ5u�ɖ�@u��	��3@u
k��!?�rHsO��@A�r{��ٿ5u�ɖ�@u��	��3@u
k��!?�rHsO��@A�r{��ٿ5u�ɖ�@u��	��3@u
k��!?�rHsO��@A�r{��ٿ5u�ɖ�@u��	��3@u
k��!?�rHsO��@�ט��ٿ_o��	�@� 7o=�3@��YLϐ!?� ����@\�`��ٿ&��tj�@�0��3@O�G�!?+�]Z���@\�`��ٿ&��tj�@�0��3@O�G�!?+�]Z���@\�`��ٿ&��tj�@�0��3@O�G�!?+�]Z���@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@�m�a�ٿ��z���@�%��S�3@�A5��!?S���*��@��@��ٿS��7(�@�j�w��3@���dv�!?bT�+ j�@��@��ٿS��7(�@�j�w��3@���dv�!?bT�+ j�@��@��ٿS��7(�@�j�w��3@���dv�!?bT�+ j�@�YHh�ٿZ5�b��@�_�.�3@} ��ɐ!?�=̽���@U��H��ٿ?Z�(���@Հ��s�3@t��I��!?+������@U��H��ٿ?Z�(���@Հ��s�3@t��I��!?+������@U��H��ٿ?Z�(���@Հ��s�3@t��I��!?+������@U��H��ٿ?Z�(���@Հ��s�3@t��I��!?+������@L���ٿ뇆r>��@'y�TT�3@�(Mv�!?�*�4P�@qe�l��ٿ	����@�*��=�3@&qE��!?�k���@qe�l��ٿ	����@�*��=�3@&qE��!?�k���@qe�l��ٿ	����@�*��=�3@&qE��!?�k���@qe�l��ٿ	����@�*��=�3@&qE��!?�k���@qe�l��ٿ	����@�*��=�3@&qE��!?�k���@�xn�P�ٿu;(v��@c�k���3@�ݹ�y�!?k��T��@�xn�P�ٿu;(v��@c�k���3@�ݹ�y�!?k��T��@#�З�ٿ�ci�3�@�0����3@j~�p͐!?J�Na��@#�З�ٿ�ci�3�@�0����3@j~�p͐!?J�Na��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@E��~j�ٿ~���@d� �p�3@��+&�!?�Ž� ��@�x�n��ٿu1o�l��@������3@fs^א!?ͳV!��@���<�ٿ���k�@?fGi'�3@�C?��!?&�҅y��@���<�ٿ���k�@?fGi'�3@�C?��!?&�҅y��@ǔ�>�ٿ!�����@���,E�3@vd[��!?#���9��@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@J�	��ٿ^���@�-<�e�3@Y�ސ!?�C��*^�@4���ٿ�4>X��@�����3@I�/�!?�[�� �@4���ٿ�4>X��@�����3@I�/�!?�[�� �@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@�]GC��ٿ��m*���@�N3��3@$J��!?(�J嘽�@��'šٿ��|��K�@�v�
S�3@��S���!?�;SiL��@��'šٿ��|��K�@�v�
S�3@��S���!?�;SiL��@��'šٿ��|��K�@�v�
S�3@��S���!?�;SiL��@��'šٿ��|��K�@�v�
S�3@��S���!?�;SiL��@}�繛ٿh��_ײ�@d|MQ�3@�2T��!?0!�t�@}�繛ٿh��_ײ�@d|MQ�3@�2T��!?0!�t�@}�繛ٿh��_ײ�@d|MQ�3@�2T��!?0!�t�@Eኩ�ٿ���T���@�ܕ��3@�	\t��!?�#ۢ޻�@E��[�ٿ�-�����@ȎW�3@�!��Ԑ!?���`2��@E��[�ٿ�-�����@ȎW�3@�!��Ԑ!?���`2��@'?&�U�ٿ�����@��b
�3@�YƳ�!?ǣ,(�5�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@���H��ٿk���E�@���'T�3@�:{-�!?�S&�rQ�@�Bz�ٿ��ϐI6�@S����3@�IX���!?�Aɾ;�@H���ܤٿji�/�@i=�"�3@�lH��!?ɳO�?V�@ŏ��ٿ=� �3�@t$��?�3@f6��א!?m�Sd��@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@���`��ٿ񧥂���@7!����3@�pfEސ!?Kf�(V�@bz��ۣٿ-� �B�@,�y=��3@�G靐!?�ET���@bz��ۣٿ-� �B�@,�y=��3@�G靐!?�ET���@bz��ۣٿ-� �B�@,�y=��3@�G靐!?�ET���@�ݏ�B�ٿt$�8y�@� ���3@�d�㷐!?��Ɍ�6�@�ݏ�B�ٿt$�8y�@� ���3@�d�㷐!?��Ɍ�6�@��y��ٿ���x�@p�Y�3@~m�p�!?J)��9�@Z���7�ٿ��|^��@p~���3@/���!?sҡZ�Y�@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@=�âߤٿj5j����@���3@��^�ؐ!?������@:Y�ɥٿ,���1��@"�ǲ�3@`�>��!?�����@:Y�ɥٿ,���1��@"�ǲ�3@`�>��!?�����@:Y�ɥٿ,���1��@"�ǲ�3@`�>��!?�����@�&i4��ٿ�"*Q�@O�!	*�3@�R�j�!?�ɕE��@�&i4��ٿ�"*Q�@O�!	*�3@�R�j�!?�ɕE��@��AU��ٿ��A�h�@��]^0�3@	4a̐!?\ճ�ű�@��AU��ٿ��A�h�@��]^0�3@	4a̐!?\ճ�ű�@��AU��ٿ��A�h�@��]^0�3@	4a̐!?\ճ�ű�@��AU��ٿ��A�h�@��]^0�3@	4a̐!?\ճ�ű�@vz&KP�ٿ�C�H�y�@lޭ,��3@_�#�!?	��P�@$�|�ٿ����M�@8�;���3@�3��!?��J��@$�|�ٿ����M�@8�;���3@�3��!?��J��@�K�狘ٿc3c���@���y��3@0NJ��!?^=t�,�@I����ٿԐ���@τ�)!�3@�YKޤ�!?j\����@k��V�ٿm�F�@��X��3@Z��)F�!?��gR�"�@k��V�ٿm�F�@��X��3@Z��)F�!?��gR�"�@k��V�ٿm�F�@��X��3@Z��)F�!?��gR�"�@k��V�ٿm�F�@��X��3@Z��)F�!?��gR�"�@�2Y�ٿ�RDJ�|�@�֓���3@>�s��!?t�aş�@�q'\�ٿ}�H��4�@ت����3@ܛ����!?m
7#���@�q'\�ٿ}�H��4�@ت����3@ܛ����!?m
7#���@�q'\�ٿ}�H��4�@ت����3@ܛ����!?m
7#���@�q'\�ٿ}�H��4�@ت����3@ܛ����!?m
7#���@�q'\�ٿ}�H��4�@ت����3@ܛ����!?m
7#���@E�L�ٿm
#"��@4�m���3@9�1֐!?����l�@E�L�ٿm
#"��@4�m���3@9�1֐!?����l�@#h3I@�ٿe�w��@P`�d�3@пs��!?O�#����@#h3I@�ٿe�w��@P`�d�3@пs��!?O�#����@zvJ���ٿ����@F`K��3@��8��!?1$.�z�@zvJ���ٿ����@F`K��3@��8��!?1$.�z�@zvJ���ٿ����@F`K��3@��8��!?1$.�z�@zvJ���ٿ����@F`K��3@��8��!?1$.�z�@�&�݋�ٿ��CN.'�@�]�d�3@~:/�!?��q�,��@�&�݋�ٿ��CN.'�@�]�d�3@~:/�!?��q�,��@%/��נٿ6_����@--�3@z��ݐ!?�h�QK�@��yg�ٿ��yjc��@���p��3@,ֿ���!?g[��@��yg�ٿ��yjc��@���p��3@,ֿ���!?g[��@���B�ٿk,�'���@2F=��3@B�d��!?(�
�4�@؎ �ٿ*�5r \�@�(�3@��OW��!?	^�L�@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@�Ъٿ�����@��l��3@I���{�!?R��i��@S���֥ٿBDktM��@�W橽�3@z=Mn�!?R�ʲ���@S���֥ٿBDktM��@�W橽�3@z=Mn�!?R�ʲ���@S���֥ٿBDktM��@�W橽�3@z=Mn�!?R�ʲ���@S���֥ٿBDktM��@�W橽�3@z=Mn�!?R�ʲ���@S���֥ٿBDktM��@�W橽�3@z=Mn�!?R�ʲ���@;g�x�ٿ�V�����@!7x�`�3@�3���!?N��C�9�@;g�x�ٿ�V�����@!7x�`�3@�3���!?N��C�9�@;g�x�ٿ�V�����@!7x�`�3@�3���!?N��C�9�@;g�x�ٿ�V�����@!7x�`�3@�3���!?N��C�9�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��&s�ٿ�G���@H�
^��3@���ex�!?�s�j�@��^��ٿ�s����@�0��y�3@-����!?[�в���@��^��ٿ�s����@�0��y�3@-����!?[�в���@��^��ٿ�s����@�0��y�3@-����!?[�в���@��^��ٿ�s����@�0��y�3@-����!?[�в���@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@���=Z�ٿ�X4s��@����3@����А!?h=Y�Y�@��8_�ٿn��o�@�le	�3@^��Ð!?r!�C �@��8_�ٿn��o�@�le	�3@^��Ð!?r!�C �@��8_�ٿn��o�@�le	�3@^��Ð!?r!�C �@��8_�ٿn��o�@�le	�3@^��Ð!?r!�C �@��8_�ٿn��o�@�le	�3@^��Ð!?r!�C �@u�hQK�ٿ�5�`���@}�Y2B�3@B�B��!?�#e=ߋ�@u�hQK�ٿ�5�`���@}�Y2B�3@B�B��!?�#e=ߋ�@D�3dT�ٿ,�&��@���v��3@�Q�ݐ!?��I��b�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@͕���ٿb�~�8z�@<�p`��3@܄0Ր!?�A��?�@�^"���ٿ���\��@��hB�3@�'��!?�F�^��@�^"���ٿ���\��@��hB�3@�'��!?�F�^��@�^"���ٿ���\��@��hB�3@�'��!?�F�^��@_:<8�ٿ���^�J�@#�Z���3@���A��!?� ���@_:<8�ٿ���^�J�@#�Z���3@���A��!?� ���@_:<8�ٿ���^�J�@#�Z���3@���A��!?� ���@ݦg� �ٿJ�����@���1�3@��]K��!?�A@�Kv�@ݦg� �ٿJ�����@���1�3@��]K��!?�A@�Kv�@ݦg� �ٿJ�����@���1�3@��]K��!?�A@�Kv�@ݦg� �ٿJ�����@���1�3@��]K��!?�A@�Kv�@���, �ٿX���@ң7
w�3@��]�!?�X�l�u�@�}@�ٿ���H�@�1���3@G��!?�'��@�g�&�ٿ܂�R�8�@QA����3@�e��/�!?��M����@�Q�I��ٿ���k`�@V�-�3@`����!?ھv�>�@�Q�I��ٿ���k`�@V�-�3@`����!?ھv�>�@�QG �ٿ렇|���@#V���3@J_���!?�����a�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@T�÷�ٿ��n ��@��I��3@���Z�!?�{��1�@����ٿz��F��@rzG%�3@��<���!?��s�q�@����ٿz��F��@rzG%�3@��<���!?��s�q�@�{���ٿ�lh����@K�j�k�3@J!H.�!?>�;��@�[�tL�ٿ΅�YA]�@(��2��3@(pM�!?>�4"ՠ�@�[�tL�ٿ΅�YA]�@(��2��3@(pM�!?>�4"ՠ�@�[�tL�ٿ΅�YA]�@(��2��3@(pM�!?>�4"ՠ�@�[�tL�ٿ΅�YA]�@(��2��3@(pM�!?>�4"ՠ�@Y�FԚ�ٿzO���@>�+�3@��p)�!?S�PA��@Y�FԚ�ٿzO���@>�+�3@��p)�!?S�PA��@M�*ߥٿ7��3�@Z�����3@��k��!?�o���@M�*ߥٿ7��3�@Z�����3@��k��!?�o���@M�*ߥٿ7��3�@Z�����3@��k��!?�o���@M�*ߥٿ7��3�@Z�����3@��k��!?�o���@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@Uy��	�ٿX�����@�L ��3@�c�Ɛ!?K�7����@�t]i�ٿ���_N*�@�.���3@a�͐!?>9�,> �@�t]i�ٿ���_N*�@�.���3@a�͐!?>9�,> �@��e��ٿ���^�@-�ͳy�3@
i�x��!?���:��@��e��ٿ���^�@-�ͳy�3@
i�x��!?���:��@��e��ٿ���^�@-�ͳy�3@
i�x��!?���:��@��e��ٿ���^�@-�ͳy�3@
i�x��!?���:��@FT����ٿ�������@lőR��3@���3��!?;�D���@FT����ٿ�������@lőR��3@���3��!?;�D���@FT����ٿ�������@lőR��3@���3��!?;�D���@FT����ٿ�������@lőR��3@���3��!?;�D���@FT����ٿ�������@lőR��3@���3��!?;�D���@���W�ٿ2s~7���@,)���3@~�����!?�5!=��@���W�ٿ2s~7���@,)���3@~�����!?�5!=��@���W�ٿ2s~7���@,)���3@~�����!?�5!=��@���W�ٿ2s~7���@,)���3@~�����!?�5!=��@���W�ٿ2s~7���@,)���3@~�����!?�5!=��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@� K0�ٿDHv�'��@�/M��3@��Q��!?��VgB��@���6��ٿ	�=Z���@�\��L�3@R/N�ې!?w4J���@��٠�ٿ2���@k^��w�3@3���!?�]�ӗ��@��٠�ٿ2���@k^��w�3@3���!?�]�ӗ��@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@�CE�ؘٿ`����@���jN�3@�KN��!?�B�r˅�@[΄�x�ٿB�~6�w�@���^�3@+�y��!?��'x9��@[΄�x�ٿB�~6�w�@���^�3@+�y��!?��'x9��@�fn^�ٿ#����M�@'��U�3@�K����!?R3��\��@�v���ٿa%�k�T�@�}�[U�3@o[�{��!?�Vq�T��@�v���ٿa%�k�T�@�}�[U�3@o[�{��!?�Vq�T��@�v���ٿa%�k�T�@�}�[U�3@o[�{��!?�Vq�T��@i��,��ٿ�w+U��@�!�;�3@v�ݖZ�!?P��)b�@i��,��ٿ�w+U��@�!�;�3@v�ݖZ�!?P��)b�@i��,��ٿ�w+U��@�!�;�3@v�ݖZ�!?P��)b�@i��,��ٿ�w+U��@�!�;�3@v�ݖZ�!?P��)b�@�ކS�ٿ���x�E�@`�4���3@ٖd�!?��Mg�@�ކS�ٿ���x�E�@`�4���3@ٖd�!?��Mg�@�ކS�ٿ���x�E�@`�4���3@ٖd�!?��Mg�@�ކS�ٿ���x�E�@`�4���3@ٖd�!?��Mg�@�ކS�ٿ���x�E�@`�4���3@ٖd�!?��Mg�@��%iR�ٿ}��ی��@�̺~�3@����ɐ!?g�XՍ�@��%iR�ٿ}��ی��@�̺~�3@����ɐ!?g�XՍ�@axA�ߙٿ�&т�f�@��S��3@����!?��[�0��@axA�ߙٿ�&т�f�@��S��3@����!?��[�0��@axA�ߙٿ�&т�f�@��S��3@����!?��[�0��@axA�ߙٿ�&т�f�@��S��3@����!?��[�0��@axA�ߙٿ�&т�f�@��S��3@����!?��[�0��@�B?��ٿ=;\�s��@vYB��3@���Z��!?PR(�l�@�B?��ٿ=;\�s��@vYB��3@���Z��!?PR(�l�@�B?��ٿ=;\�s��@vYB��3@���Z��!?PR(�l�@�B?��ٿ=;\�s��@vYB��3@���Z��!?PR(�l�@Q��I�ٿ9���c�@���3@5 ؐ!?�q^��@Q��I�ٿ9���c�@���3@5 ؐ!?�q^��@�b
b�ٿp��;��@C]G�(�3@��sai�!?W+��~�@�b
b�ٿp��;��@C]G�(�3@��sai�!?W+��~�@�x��ٿ�_�^��@�!p�W�3@�\�̇�!?G*>��@�*K۩ٿ��D�#�@1���3@��I��!?TT���I�@�*K۩ٿ��D�#�@1���3@��I��!?TT���I�@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@Jv�:�ٿ��,[h��@%��x��3@�<J��!?�hRxD��@�����ٿ�5����@J��,)�3@w,�X��!?��r6�5�@�px�ٿ���On��@Qxз��3@kԁ'��!?:wI��e�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@\����ٿr"f���@G>_�1�3@�p���!?`�e�l�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���l�ٿ�.��]�@�t��3@Q��ݠ�!?NB��~�@���Rڛٿ��Db��@�	��3@�D%�!?�������@���Rڛٿ��Db��@�	��3@�D%�!?�������@���Rڛٿ��Db��@�	��3@�D%�!?�������@���Rڛٿ��Db��@�	��3@�D%�!?�������@���Rڛٿ��Db��@�	��3@�D%�!?�������@7��'�ٿF*���@aNK��3@�T�ː!?��S�đ�@7��'�ٿF*���@aNK��3@�T�ː!?��S�đ�@7��'�ٿF*���@aNK��3@�T�ː!?��S�đ�@7��'�ٿF*���@aNK��3@�T�ː!?��S�đ�@7��'�ٿF*���@aNK��3@�T�ː!?��S�đ�@���y��ٿ�=�����@�l�;��3@'}��q�!?�*��u��@���y��ٿ�=�����@�l�;��3@'}��q�!?�*��u��@w��� �ٿO����Z�@d�D���3@75���!?�6.g��@w��� �ٿO����Z�@d�D���3@75���!?�6.g��@w��� �ٿO����Z�@d�D���3@75���!?�6.g��@�듞n�ٿ����$�@���3@+@Ry��!?.�\"�@�듞n�ٿ����$�@���3@+@Ry��!?.�\"�@��pc.�ٿ�IoH�@BnPA��3@Pq^��!?T���
��@��pc.�ٿ�IoH�@BnPA��3@Pq^��!?T���
��@��pc.�ٿ�IoH�@BnPA��3@Pq^��!?T���
��@��pc.�ٿ�IoH�@BnPA��3@Pq^��!?T���
��@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@^���v�ٿzgbz��@M A���3@�;E��!?#���r�@�`�
ěٿ����xp�@W�����3@ � ��!?���,N~�@�`�
ěٿ����xp�@W�����3@ � ��!?���,N~�@�`�
ěٿ����xp�@W�����3@ � ��!?���,N~�@�`�
ěٿ����xp�@W�����3@ � ��!?���,N~�@ϧ�śٿo�N��@�0���3@�k���!?OQ�"�u�@ϧ�śٿo�N��@�0���3@�k���!?OQ�"�u�@ϧ�śٿo�N��@�0���3@�k���!?OQ�"�u�@ϧ�śٿo�N��@�0���3@�k���!?OQ�"�u�@F�T�ٿ�5P]-z�@t+�a��3@ w�!?�� 'A��@F�T�ٿ�5P]-z�@t+�a��3@ w�!?�� 'A��@F�T�ٿ�5P]-z�@t+�a��3@ w�!?�� 'A��@F�T�ٿ�5P]-z�@t+�a��3@ w�!?�� 'A��@F�T�ٿ�5P]-z�@t+�a��3@ w�!?�� 'A��@#.f�V�ٿ� �"l�@��$�3@$m4v��!?|�5��@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�p`8�ٿj���`�@約"�3@x铗Ő!?�bB_�@�y�i�ٿs"H�F�@S@�s�3@�5�ސ!?��ͦ�N�@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@tNݡٿ������@O�7�C�3@v1)'̐!?�_���@���P�ٿk�#�m��@�Y
��3@�4r�!?�!���!�@�@�h�ٿ�P���@�����3@¨���!?�݈6� �@�@�h�ٿ�P���@�����3@¨���!?�݈6� �@�@�h�ٿ�P���@�����3@¨���!?�݈6� �@�n5Řٿ���>�V�@�����3@�X���!?��7�
�@�n5Řٿ���>�V�@�����3@�X���!?��7�
�@�n5Řٿ���>�V�@�����3@�X���!?��7�
�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@����u�ٿe�N�|�@���8��3@"Q���!?��P-�l�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@)F����ٿ�� �[�@H�6C�3@��d9�!?)��)�7�@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@������ٿ��9x�@$��d�3@9Jc��!?��O���@�s��s�ٿ�%��+��@qdb�a�3@a�`�)�!?:�jƦ[�@�s��s�ٿ�%��+��@qdb�a�3@a�`�)�!?:�jƦ[�@�s��s�ٿ�%��+��@qdb�a�3@a�`�)�!?:�jƦ[�@�s��s�ٿ�%��+��@qdb�a�3@a�`�)�!?:�jƦ[�@�s��s�ٿ�%��+��@qdb�a�3@a�`�)�!?:�jƦ[�@���r?�ٿ��ǳEg�@#b���3@[L�]�!?��r�t��@4��[��ٿ��"�v?�@`
����3@q##�!?K�U���@4��[��ٿ��"�v?�@`
����3@q##�!?K�U���@4��[��ٿ��"�v?�@`
����3@q##�!?K�U���@4��[��ٿ��"�v?�@`
����3@q##�!?K�U���@ϯ,F�ٿt�p@��@H���3@��{T�!?/�${|j�@��f�(�ٿ���<��@a��P}�3@� ��!?�t%s�X�@��f�(�ٿ���<��@a��P}�3@� ��!?�t%s�X�@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@�X�B�ٿ��cj�&�@�j����3@�^��ِ!?�^p����@���o��ٿx[R~�4�@N�0"�3@��� ��!?kT�߉�@���o��ٿx[R~�4�@N�0"�3@��� ��!?kT�߉�@���o��ٿx[R~�4�@N�0"�3@��� ��!?kT�߉�@�z���ٿ1;h���@"o�}�3@C����!?e��ѭ�@�?�5�ٿ���¹�@�<�J�3@��
�!?�sN�:��@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��1	e�ٿ����j�@or0D�3@E�M"�!?�tه�@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@��q��ٿ��ۺ�]�@��E�3@~��$��!?2}`��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@���=�ٿ[��j�@U�7��3@����c�!?�遅��@��6`�ٿ��M%U�@~�HM8�3@&%�qW�!?E�ɾ�@��6`�ٿ��M%U�@~�HM8�3@&%�qW�!?E�ɾ�@��6`�ٿ��M%U�@~�HM8�3@&%�qW�!?E�ɾ�@��6`�ٿ��M%U�@~�HM8�3@&%�qW�!?E�ɾ�@��6`�ٿ��M%U�@~�HM8�3@&%�qW�!?E�ɾ�@y��z��ٿ��?0��@�hؿ-�3@�nH�!?VK#%��@y��z��ٿ��?0��@�hؿ-�3@�nH�!?VK#%��@"IQ���ٿ���o���@��s�	�3@X|���!?���U�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@*�\���ٿ�~��@Ao�N�3@����!?b�ǈGU�@�g�!��ٿy?�����@�'=8��3@�Hʧ:�!?��P��u�@�;+(�ٿ���3@��@dp¸��3@��	D�!??�b���@�;+(�ٿ���3@��@dp¸��3@��	D�!??�b���@�;+(�ٿ���3@��@dp¸��3@��	D�!??�b���@�q��^�ٿ~��q��@`��j��3@o�C��!?$3�v{�@t�Q��ٿ3�ܒE�@X��L��3@��]8u�!?��jR���@t�Q��ٿ3�ܒE�@X��L��3@��]8u�!?��jR���@t�Q��ٿ3�ܒE�@X��L��3@��]8u�!?��jR���@t�Q��ٿ3�ܒE�@X��L��3@��]8u�!?��jR���@��Oq�ٿ^�WF%��@$��%�3@���?��!?�W�|j�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@"�4a�ٿ���s2�@�9x��3@��2��!?�F���B�@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@��LKX�ٿ>H�	�=�@OS*���3@g�\��!?�U�9��@����ٿ3q�.tZ�@��&���3@�.+�!?�o��b��@�`Ҟ��ٿ�#/�c?�@G̰d�3@�Pf���!?Y��?���@�`Ҟ��ٿ�#/�c?�@G̰d�3@�Pf���!?Y��?���@�`Ҟ��ٿ�#/�c?�@G̰d�3@�Pf���!?Y��?���@�r5�4�ٿ�&���K�@�KY(��3@ ��&�!?�ش�L�@�r5�4�ٿ�&���K�@�KY(��3@ ��&�!?�ش�L�@�r5�4�ٿ�&���K�@�KY(��3@ ��&�!?�ش�L�@���鄠ٿ$�]Ly��@f�5���3@��Ĺb�!?n��@ח�@���鄠ٿ$�]Ly��@f�5���3@��Ĺb�!?n��@ח�@���鄠ٿ$�]Ly��@f�5���3@��Ĺb�!?n��@ח�@���鄠ٿ$�]Ly��@f�5���3@��Ĺb�!?n��@ח�@�0�I�ٿZ`�%}��@B' �9�3@�B���!?� ��c�@�0�I�ٿZ`�%}��@B' �9�3@�B���!?� ��c�@�0�I�ٿZ`�%}��@B' �9�3@�B���!?� ��c�@�0�I�ٿZ`�%}��@B' �9�3@�B���!?� ��c�@X��}Ťٿ���5��@]�C��3@���n�!?SH�vK��@X��}Ťٿ���5��@]�C��3@���n�!?SH�vK��@X��}Ťٿ���5��@]�C��3@���n�!?SH�vK��@X��}Ťٿ���5��@]�C��3@���n�!?SH�vK��@D��*8�ٿ��T�g��@Q��v(�3@I�>`��!?��~��@D��*8�ٿ��T�g��@Q��v(�3@I�>`��!?��~��@D��*8�ٿ��T�g��@Q��v(�3@I�>`��!?��~��@D��*8�ٿ��T�g��@Q��v(�3@I�>`��!?��~��@D��*8�ٿ��T�g��@Q��v(�3@I�>`��!?��~��@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��J#�ٿ���( �@�����3@+��z�!?|c��f�@��?�ٿ.��y~��@v5��3@t@/��!?��,��h�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@P���ٿL�>��`�@<�����3@<��ϐ!?ˮ܀�#�@��&Ո�ٿQ7�J�&�@ߔ"�~�3@*6�ɛ�!?�tl#���@��&Ո�ٿQ7�J�&�@ߔ"�~�3@*6�ɛ�!?�tl#���@�0���ٿ�����@n�����3@
��c��!?�6����@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��_�r�ٿ�tT�%|�@�d����3@u��q�!?t0٤���@��L�]�ٿ���z��@�"l���3@��p��!?�D��2u�@��L�]�ٿ���z��@�"l���3@��p��!?�D��2u�@��L�]�ٿ���z��@�"l���3@��p��!?�D��2u�@��L�]�ٿ���z��@�"l���3@��p��!?�D��2u�@��t�ٿW�W�7��@Ȥ<�'�3@�0�Đ!?O�=�-^�@��.~�ٿ*^���@����y�3@�ËQ��!?��mO}�@��.~�ٿ*^���@����y�3@�ËQ��!?��mO}�@��.~�ٿ*^���@����y�3@�ËQ��!?��mO}�@l"4�ٿ������@-�~s�3@��ِ!?r8�-���@l"4�ٿ������@-�~s�3@��ِ!?r8�-���@�l�(2�ٿW7u����@'lf��3@PArߐ!?�ɷ�DW�@�l�(2�ٿW7u����@'lf��3@PArߐ!?�ɷ�DW�@81u�j�ٿN�u��@�/�3@w����!?M�w�d��@.����ٿ8h78�O�@��E��3@�
�ɐ!?�خ�h�@.����ٿ8h78�O�@��E��3@�
�ɐ!?�خ�h�@.����ٿ8h78�O�@��E��3@�
�ɐ!?�خ�h�@.����ٿ8h78�O�@��E��3@�
�ɐ!?�خ�h�@S9'-��ٿ�N����@'U~c�3@g��Ɛ!?r�y��@S9'-��ٿ�N����@'U~c�3@g��Ɛ!?r�y��@S9'-��ٿ�N����@'U~c�3@g��Ɛ!?r�y��@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@9���ٿ��_�(H�@RK�W�3@���!?|��~�=�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@��$�)�ٿ���71��@��&���3@QH���!?�DiU�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@�JIR�ٿ�ɿf�p�@�kLo��3@�b��!?���ߘ�@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@��@`g�ٿ�Jox:�@d��Z�3@T�V��!?���{���@:A����ٿ	�Y��@n.����3@�kv�!?��Y>�@:A����ٿ	�Y��@n.����3@�kv�!?��Y>�@:A����ٿ	�Y��@n.����3@�kv�!?��Y>�@:A����ٿ	�Y��@n.����3@�kv�!?��Y>�@:A����ٿ	�Y��@n.����3@�kv�!?��Y>�@;*�B�ٿ�dZH��@4�����3@�s�=��!?��F����@;*�B�ٿ�dZH��@4�����3@�s�=��!?��F����@���r��ٿ	*�]?��@���D��3@�>�!?P�?\{(�@)d3A�ٿ62-ŧ��@[����3@��ϋڐ!?���<*	�@)d3A�ٿ62-ŧ��@[����3@��ϋڐ!?���<*	�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@��xa�ٿhbR/�@_��h�3@b{`א!?��f�^#�@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@����ٿ�_�~,��@
+�3@���ސ!?ڟ�V��@�+؝�ٿk�2x�@�N&���3@��qdƐ!?�b@�+�@�+؝�ٿk�2x�@�N&���3@��qdƐ!?�b@�+�@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@�K��ٿ�;��V�@;��e�3@
����!?J���H��@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@<���]�ٿ��73�@4��j�3@LC���!?+ÚE�m�@�]��Ϙٿ�����h�@�s�p��3@7�����!?v	��u�@�]��Ϙٿ�����h�@�s�p��3@7�����!?v	��u�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@���=�ٿv_��.�@}�OR�3@�����!?�ԕ��d�@G��%�ٿV��/�R�@�gJ���3@��ؐ!?2����@���.&�ٿ)w��C�@���c�3@����!?��o`v��@���.&�ٿ)w��C�@���c�3@����!?��o`v��@���.&�ٿ)w��C�@���c�3@����!?��o`v��@��H�-�ٿ}�7k��@��q�3@1�p�!�!?�(J"��@���Ē�ٿDw���@	a!��3@�k�
�!?��a�c�@���Ē�ٿDw���@	a!��3@�k�
�!?��a�c�@���Ē�ٿDw���@	a!��3@�k�
�!?��a�c�@�����ٿT�;�)�@ʔ A�3@vX%�ؐ!?/���S#�@C�K��ٿ!k�f8�@Za�C�3@��^�j�!?��䎯�@�d�Cˤٿ�n��.��@N�f!��3@�Zj
��!?����
�@�d�Cˤٿ�n��.��@N�f!��3@�Zj
��!?����
�@�d�Cˤٿ�n��.��@N�f!��3@�Zj
��!?����
�@�d�Cˤٿ�n��.��@N�f!��3@�Zj
��!?����
�@�vbӧٿ�|p�$��@��ӻ��3@���!?�T�����@�vbӧٿ�|p�$��@��ӻ��3@���!?�T�����@�vbӧٿ�|p�$��@��ӻ��3@���!?�T�����@�vbӧٿ�|p�$��@��ӻ��3@���!?�T�����@:��}�ٿ��=bP��@�ƞ���3@e��Ȑ!?��!�@�@:��}�ٿ��=bP��@�ƞ���3@e��Ȑ!?��!�@�@:��}�ٿ��=bP��@�ƞ���3@e��Ȑ!?��!�@�@:��}�ٿ��=bP��@�ƞ���3@e��Ȑ!?��!�@�@:��}�ٿ��=bP��@�ƞ���3@e��Ȑ!?��!�@�@Z@�P�ٿ:(z/[s�@� �IG�3@��x��!?���{p�@Z@�P�ٿ:(z/[s�@� �IG�3@��x��!?���{p�@�P��B�ٿ�S5MG�@��v��3@���!?oV���@�P��B�ٿ�S5MG�@��v��3@���!?oV���@�P��B�ٿ�S5MG�@��v��3@���!?oV���@�P��B�ٿ�S5MG�@��v��3@���!?oV���@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@P�Aˡٿ���'�@�WF���3@�5����!? ������@��F���ٿ������@.�����3@8���ǐ!?�U(��@��F���ٿ������@.�����3@8���ǐ!?�U(��@��F���ٿ������@.�����3@8���ǐ!?�U(��@����f�ٿו����@�)l���3@|��!?� �1��@� :��ٿ��d�O�@���/��3@��)�!?�u[��@� :��ٿ��d�O�@���/��3@��)�!?�u[��@� :��ٿ��d�O�@���/��3@��)�!?�u[��@� :��ٿ��d�O�@���/��3@��)�!?�u[��@� :��ٿ��d�O�@���/��3@��)�!?�u[��@�K{�V�ٿ�tΙk�@@n��3@U�U%ϐ!?6Y4[���@�K{�V�ٿ�tΙk�@@n��3@U�U%ϐ!?6Y4[���@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@ʳ6D%�ٿ��O{ �@�4]��3@��O3��!?DvG����@�M��ٿɍ�\1�@����3@�I4P��!?U}9����@\f�N#�ٿ���d|��@���v��3@v,&�s�!?a��﯐�@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@�+N�|�ٿ��#_�@*>[ˍ�3@�0�ː!?ٺA���@#����ٿ�O��rh�@IhO��3@	$[�!?���`�	�@#����ٿ�O��rh�@IhO��3@	$[�!?���`�	�@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@]EN�h�ٿ�Y���@�;���3@J��Ȑ!?�����@eE��d�ٿ.��f��@�)�L<�3@�B��Ր!?-1Ma��@�m��o�ٿ�����@��ī��3@�4F��!?V?:����@�O"��ٿ�Z����@����?�3@���!?����9��@�O"��ٿ�Z����@����?�3@���!?����9��@�O"��ٿ�Z����@����?�3@���!?����9��@�O"��ٿ�Z����@����?�3@���!?����9��@ebF�ٿ!�H�>v�@=˃<��3@��uǐ!?+Ji���@�<���ٿ��V�"��@�Ȋ|W�3@�jn�ː!?��65�;�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@T��SF�ٿS�}9���@s��/�3@�h��!?�g9�@�]<�L�ٿ^#�C@��@���V�3@���ڐ!?�cFpI��@���	�ٿ�&�����@y�V���3@�-&B��!?tc��G��@WL� Ȥٿ�$�Z�@�<�x�3@e#�'��!?���p�@�B!�O�ٿ:m9 ^�@�Y `'�3@Uy���!?�o5����@�B!�O�ٿ:m9 ^�@�Y `'�3@Uy���!?�o5����@�B!�O�ٿ:m9 ^�@�Y `'�3@Uy���!?�o5����@�B!�O�ٿ:m9 ^�@�Y `'�3@Uy���!?�o5����@�B!�O�ٿ:m9 ^�@�Y `'�3@Uy���!?�o5����@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@N0�B��ٿL��j�@�Y~�x�3@y�`�!?�O)Ԁ��@~�T�5�ٿ�X�)�@P؇�r�3@��X��!?��z�@~�T�5�ٿ�X�)�@P؇�r�3@��X��!?��z�@l����ٿ��Vw$F�@x��"��3@4��A��!?F�W��@l����ٿ��Vw$F�@x��"��3@4��A��!?F�W��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@�����ٿqp�[ ��@�4]��3@���s
�!?���	��@vp�8�ٿ3$��ʺ�@�;�\�3@��H���!?0� kT�@vp�8�ٿ3$��ʺ�@�;�\�3@��H���!?0� kT�@vp�8�ٿ3$��ʺ�@�;�\�3@��H���!?0� kT�@vp�8�ٿ3$��ʺ�@�;�\�3@��H���!?0� kT�@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@���H�ٿV�w��&�@s�2l�3@���ݯ�!?�J�h���@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@%�e<�ٿp�b���@a�
���3@��w���!?��2v5��@��:���ٿ%~H	���@���+�3@���Ɛ!?6�.`<��@��:���ٿ%~H	���@���+�3@���Ɛ!?6�.`<��@��:���ٿ%~H	���@���+�3@���Ɛ!?6�.`<��@��:���ٿ%~H	���@���+�3@���Ɛ!?6�.`<��@��:���ٿ%~H	���@���+�3@���Ɛ!?6�.`<��@�����ٿQk:bf�@�>�tg�3@=��ѐ!?��6��C�@�����ٿQk:bf�@�>�tg�3@=��ѐ!?��6��C�@�����ٿQk:bf�@�>�tg�3@=��ѐ!?��6��C�@�����ٿQk:bf�@�>�tg�3@=��ѐ!?��6��C�@���'��ٿk����`�@�{���3@��H�!?�L*�Q1�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@�%P���ٿ�s��W�@����@�3@�˳^��!?�RKyr�@����ٿ�^{��O�@��Z&�3@��L��!?U�N%|��@����ٿ�^{��O�@��Z&�3@��L��!?U�N%|��@ܨy靖ٿۆ{Cϧ�@���v�3@h6܂Đ!?S�fc���@r� ��ٿ�-�~Ҵ�@y�  �3@��'�!?�S�{)A�@�R�@w�ٿƸb�w�@�HP��3@�#��!?������@�R�@w�ٿƸb�w�@�HP��3@�#��!?������@jW���ٿ׉")�@M�qws�3@�+����!?�X�����@jW���ٿ׉")�@M�qws�3@�+����!?�X�����@�{��t�ٿC�|'O��@�(����3@NOb\�!?d��$��@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@�>�ٿN�b�T��@Xkޒ_�3@[��!?~��1�@E�T ޝٿ^1�����@f+���3@�q.w��!?�* ��S�@E�T ޝٿ^1�����@f+���3@�q.w��!?�* ��S�@E�T ޝٿ^1�����@f+���3@�q.w��!?�* ��S�@E�T ޝٿ^1�����@f+���3@�q.w��!?�* ��S�@2)w��ٿ�=G��@zP{4@�a�-�!?��:�z��@�F�<n�ٿؗ��@�';��3@�"%�<�!?&���d�@�F�<n�ٿؗ��@�';��3@�"%�<�!?&���d�@�F�<n�ٿؗ��@�';��3@�"%�<�!?&���d�@�F�<n�ٿؗ��@�';��3@�"%�<�!?&���d�@�e��ٿ�s_�Hc�@������3@=`_���!?��H���@�e��ٿ�s_�Hc�@������3@=`_���!?��H���@�e��ٿ�s_�Hc�@������3@=`_���!?��H���@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@A'��ٿ����@�mB<��3@(%@;��!?~��z� �@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@WG�0��ٿ7��f�@f��%��3@��*�!?�p���@z�nx��ٿ���rW��@�5�Q��3@�G��Ɛ!?!z�s�@�C{!x�ٿtV�X���@�C���3@o�%�!?�>$g���@�C{!x�ٿtV�X���@�C���3@o�%�!?�>$g���@�C{!x�ٿtV�X���@�C���3@o�%�!?�>$g���@�C{!x�ٿtV�X���@�C���3@o�%�!?�>$g���@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@�^�Ѻ�ٿ�;���>�@"9�%�3@�9 �!?Ra��$�@��"���ٿ�/Ro"�@>eI���3@|!bZ�!?�I���@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@�`)ֻ�ٿ�0���.�@,���p�3@,P(��!?�\����@&�S�ٿ3�GJ�@)�x_��3@���̐!?VM��@&�S�ٿ3�GJ�@)�x_��3@���̐!?VM��@&�S�ٿ3�GJ�@)�x_��3@���̐!?VM��@�U3F=�ٿd
����@(����3@��S���!?�V�@�U3F=�ٿd
����@(����3@��S���!?�V�@�U3F=�ٿd
����@(����3@��S���!?�V�@�U3F=�ٿd
����@(����3@��S���!?�V�@�U3F=�ٿd
����@(����3@��S���!?�V�@�U3F=�ٿd
����@(����3@��S���!?�V�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@1n�Țٿ��\���@����>�3@�T����!?��wzF;�@���GԘٿ:����@��?f��3@�A�!?k	R�/	�@���GԘٿ:����@��?f��3@�A�!?k	R�/	�@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@w�MA�ٿd;#����@��ß��3@�ىА!?E�tn��@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@��F�١ٿ�����@bI���3@���5�!?�vv|�@���?�ٿA��%'!�@��5���3@����!?���Dq��@��H���ٿ�=$��@���	�3@؀�b��!?2������@�6�q�ٿ]�.��@��_��3@���܀�!?ہn�[��@��u:ˤٿN!�0i.�@�����3@�"�r��!?NjL~��@��u:ˤٿN!�0i.�@�����3@�"�r��!?NjL~��@<�$$�ٿ�6�Xc#�@�"��3@���.��!?�l+���@<�$$�ٿ�6�Xc#�@�"��3@���.��!?�l+���@<�$$�ٿ�6�Xc#�@�"��3@���.��!?�l+���@�s�[�ٿdkk�P�@k1���3@��K�Ӑ!?V��.���@�s�[�ٿdkk�P�@k1���3@��K�Ӑ!?V��.���@F�3��ٿ1��`b�@����3@�e��ɐ!?�g5�6t�@F�3��ٿ1��`b�@����3@�e��ɐ!?�g5�6t�@F�3��ٿ1��`b�@����3@�e��ɐ!?�g5�6t�@F�3��ٿ1��`b�@����3@�e��ɐ!?�g5�6t�@F�3��ٿ1��`b�@����3@�e��ɐ!?�g5�6t�@jw�B��ٿV(ǩ0+�@�5�I�3@6#��ސ!?�ҥ�=��@jw�B��ٿV(ǩ0+�@�5�I�3@6#��ސ!?�ҥ�=��@jw�B��ٿV(ǩ0+�@�5�I�3@6#��ސ!?�ҥ�=��@jw�B��ٿV(ǩ0+�@�5�I�3@6#��ސ!?�ҥ�=��@jw�B��ٿV(ǩ0+�@�5�I�3@6#��ސ!?�ҥ�=��@����ٿFӒ�b�@I�*�|�3@U<n̐!?�Z��k�@����ٿFӒ�b�@I�*�|�3@U<n̐!?�Z��k�@����ٿFӒ�b�@I�*�|�3@U<n̐!?�Z��k�@����ٿFӒ�b�@I�*�|�3@U<n̐!?�Z��k�@����ٿFӒ�b�@I�*�|�3@U<n̐!?�Z��k�@T�vb��ٿ߅k)��@û@�~�3@��Hc֐!?�� �a�@T�vb��ٿ߅k)��@û@�~�3@��Hc֐!?�� �a�@T�vb��ٿ߅k)��@û@�~�3@��Hc֐!?�� �a�@T�vb��ٿ߅k)��@û@�~�3@��Hc֐!?�� �a�@�.�H�ٿ(�UBd�@�`&�C�3@�_�А!?�<�1�K�@�.�H�ٿ(�UBd�@�`&�C�3@�_�А!?�<�1�K�@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�7�q�ٿ- A��@������3@�#���!?���F���@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�O�(,�ٿ�����@^�\���3@�X�j��!?�������@�����ٿ������@����3@��ڐ!?�˶�"�@�����ٿ������@����3@��ڐ!?�˶�"�@�����ٿ������@����3@��ڐ!?�˶�"�@�����ٿ������@����3@��ڐ!?�˶�"�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@��4��ٿ���@�u ��3@�J�W��!?��*LF�@`��şٿ/hwOQ��@	�����3@w'�e��!?�ݨ b�@`��şٿ/hwOQ��@	�����3@w'�e��!?�ݨ b�@`��şٿ/hwOQ��@	�����3@w'�e��!?�ݨ b�@3�bu�ٿ�����@������3@j�
��!?u�U����@3�bu�ٿ�����@������3@j�
��!?u�U����@���p�ٿx��7���@}H�u�3@г���!?No���7�@���p�ٿx��7���@}H�u�3@г���!?No���7�@���p�ٿx��7���@}H�u�3@г���!?No���7�@���p�ٿx��7���@}H�u�3@г���!?No���7�@���
�ٿ&&%��@{Q�:e�3@R3�?�!?	�O$4��@��	0�ٿ�]�-���@�K���3@����!?җ����@�� ���ٿ���A�F�@o碸�3@)2��ܐ!?�H^l�@*�@�G�ٿ�����@�����3@��M,��!?ߖ�o���@��Yk�ٿZ�+�"�@�C](��3@��ϔ�!?��a��@��Yk�ٿZ�+�"�@�C](��3@��ϔ�!?��a��@��Yk�ٿZ�+�"�@�C](��3@��ϔ�!?��a��@��Yk�ٿZ�+�"�@�C](��3@��ϔ�!?��a��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@&8�x9�ٿF����X�@���3@ܰ���!?�X�z��@1,_�)�ٿ�� �)�@W^C�3@>����!?�D����@b�^Ùٿ�\��V#�@��Q��3@�ˡ��!?/�"�T�@�6C�ٿ���<Ol�@�!ڱ��3@
T�Ր!?7\�(.��@�6C�ٿ���<Ol�@�!ڱ��3@
T�Ր!?7\�(.��@�6C�ٿ���<Ol�@�!ڱ��3@
T�Ր!?7\�(.��@���?�ٿ���Da�@�K��g�3@&\ɐ!?� �i]~�@'�Y�͜ٿrt�6��@��nlb�3@
��(��!?.���g4�@'�Y�͜ٿrt�6��@��nlb�3@
��(��!?.���g4�@'�Y�͜ٿrt�6��@��nlb�3@
��(��!?.���g4�@�)ZT5�ٿ�����@�'����3@;)��!?�^���L�@�)ZT5�ٿ�����@�'����3@;)��!?�^���L�@�n�s�ٿh�p��@Y;#p��3@JS��!?H�F~��@�n�s�ٿh�p��@Y;#p��3@JS��!?H�F~��@�n�s�ٿh�p��@Y;#p��3@JS��!?H�F~��@�n�s�ٿh�p��@Y;#p��3@JS��!?H�F~��@�n�s�ٿh�p��@Y;#p��3@JS��!?H�F~��@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@5Ҵu�ٿt��\�W�@�̦���3@���^�!?�u]�M�@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@��jE~�ٿ�P��Nu�@�r��3@�hS�!?�?�Y��@����ٿ�Tl.b�@b��2�3@J4��!?*�Ot���@����ٿ�Tl.b�@b��2�3@J4��!?*�Ot���@����ٿ�Tl.b�@b��2�3@J4��!?*�Ot���@bXn�ٿ>�¤���@�f�`z�3@_!;=�!?��§���@bXn�ٿ>�¤���@�f�`z�3@_!;=�!?��§���@bXn�ٿ>�¤���@�f�`z�3@_!;=�!?��§���@���;�ٿ:��q���@��C�3@G<J/�!?����\��@���;�ٿ:��q���@��C�3@G<J/�!?����\��@���;�ٿ:��q���@��C�3@G<J/�!?����\��@'���)�ٿ�'qGĮ�@Ah(�T�3@�8���!?|�&�|B�@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�8�6��ٿ4Ɓm��@���&��3@}A�:�!?�����@�w��F�ٿ�NU�Ι�@����`�3@�_���!?��'8��@8aUNџٿ��]%���@#cd��3@��֐!?V�Ӆ?�@��ɉ�ٿ�$��Z�@ʩ%G1�3@�τ���!?�9���@��ɉ�ٿ�$��Z�@ʩ%G1�3@�τ���!?�9���@��ɉ�ٿ�$��Z�@ʩ%G1�3@�τ���!?�9���@f!��ٿ_�k{V�@���P�3@W2���!?�4�k�N�@f!��ٿ_�k{V�@���P�3@W2���!?�4�k�N�@���&�ٿ�!�a��@�r�D��3@Orn�Ɛ!?rr�����@���&�ٿ�!�a��@�r�D��3@Orn�Ɛ!?rr�����@���&�ٿ�!�a��@�r�D��3@Orn�Ɛ!?rr�����@���&�ٿ�!�a��@�r�D��3@Orn�Ɛ!?rr�����@�F��ݥٿmz�@&$�@�݌V(�3@�殐!?�;���@�F��ݥٿmz�@&$�@�݌V(�3@�殐!?�;���@�F��ݥٿmz�@&$�@�݌V(�3@�殐!?�;���@��2�ٿª��@�i���3@x�z���!?�9j�K��@��2�ٿª��@�i���3@x�z���!?�9j�K��@��2�ٿª��@�i���3@x�z���!?�9j�K��@��2�ٿª��@�i���3@x�z���!?�9j�K��@��2�ٿª��@�i���3@x�z���!?�9j�K��@��2�ٿª��@�i���3@x�z���!?�9j�K��@B%�n��ٿ�ߖ4���@�xAE�3@ee�=��!?��:���@B%�n��ٿ�ߖ4���@�xAE�3@ee�=��!?��:���@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@.K:Jǝٿ}i�gLN�@Y�z��3@����!?�	�B#�@Qw�.u�ٿ\�u��8�@�l��U�3@�>ݐ!?Kf��2�@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@�0~�ٿ����H��@�74���3@��D1Ɛ!?�&�n��@���?�ٿj����>�@�6�H��3@bnw�Ð!?��<D�M�@���?�ٿj����>�@�6�H��3@bnw�Ð!?��<D�M�@���?�ٿj����>�@�6�H��3@bnw�Ð!?��<D�M�@�JM�ٿ�,�[��@�?�^��3@�t���!?���An"�@�JM�ٿ�,�[��@�?�^��3@�t���!?���An"�@�JM�ٿ�,�[��@�?�^��3@�t���!?���An"�@�JM�ٿ�,�[��@�?�^��3@�t���!?���An"�@g6B��ٿ�K^>���@4Ze^�3@,�D���!?뿉�3�@��:;�ٿx�w���@�ug�(�3@$a��!?�)�e&�@��L���ٿq�S���@` I���3@+U�F��!?���.޶�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@a����ٿI�.L�D�@���Y��3@.�̐!?XA]�2�@e�C'֞ٿ�K����@t�e��3@-e_���!?	�-���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Ӧz�)�ٿ~y�Y���@��37r�3@Ť�%��!?
���@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@Z�}�R�ٿ�'��2�@���<��3@�����!?��A�y��@i�zQ�ٿ�^���@%�'&��3@��ʧ�!?4|a���@i�zQ�ٿ�^���@%�'&��3@��ʧ�!?4|a���@i�zQ�ٿ�^���@%�'&��3@��ʧ�!?4|a���@i�zQ�ٿ�^���@%�'&��3@��ʧ�!?4|a���@i�zQ�ٿ�^���@%�'&��3@��ʧ�!?4|a���@_��b��ٿ�ԅ*��@����	�3@���h��!?�Y�*��@�~5m�ٿ��*�k�@�@�D3�3@�[�ϐ!?`q�z���@�~5m�ٿ��*�k�@�@�D3�3@�[�ϐ!?`q�z���@�~5m�ٿ��*�k�@�@�D3�3@�[�ϐ!?`q�z���@�~5m�ٿ��*�k�@�@�D3�3@�[�ϐ!?`q�z���@����ٿ��"N�@��)��3@�i�Ӑ!?�HIDM{�@����ٿ��"N�@��)��3@�i�Ӑ!?�HIDM{�@g̲L/�ٿPݾfX��@�n�>�3@��h�Ԑ!?�
}�LE�@g̲L/�ٿPݾfX��@�n�>�3@��h�Ԑ!?�
}�LE�@g̲L/�ٿPݾfX��@�n�>�3@��h�Ԑ!?�
}�LE�@g̲L/�ٿPݾfX��@�n�>�3@��h�Ԑ!?�
}�LE�@�is2�ٿC�4�@���E��3@���I��!?,��p,m�@�is2�ٿC�4�@���E��3@���I��!?,��p,m�@�is2�ٿC�4�@���E��3@���I��!?,��p,m�@�is2�ٿC�4�@���E��3@���I��!?,��p,m�@�M�nڝٿ�*��y�@o�O�3@,nz}��!?i�M�W�@�M�nڝٿ�*��y�@o�O�3@,nz}��!?i�M�W�@�M�nڝٿ�*��y�@o�O�3@,nz}��!?i�M�W�@�M�nڝٿ�*��y�@o�O�3@,nz}��!?i�M�W�@sn	���ٿ3��;	��@��);�3@c��kː!?��+���@sn	���ٿ3��;	��@��);�3@c��kː!?��+���@�;�@�ٿcی�ʁ�@�'U��3@���S�!?d�uF��@�;�@�ٿcی�ʁ�@�'U��3@���S�!?d�uF��@��ԣ��ٿ���7`�@�u�3@tOs ��!?�_�S�o�@��q���ٿ�YkOjB�@�U�'Z�3@�N�ő�!?�@����@��q���ٿ�YkOjB�@�U�'Z�3@�N�ő�!?�@����@;���i�ٿ��n��O�@�<9��3@�yA��!?��]փ�@;���i�ٿ��n��O�@�<9��3@�yA��!?��]փ�@;���i�ٿ��n��O�@�<9��3@�yA��!?��]փ�@;���i�ٿ��n��O�@�<9��3@�yA��!?��]փ�@;���i�ٿ��n��O�@�<9��3@�yA��!?��]փ�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@��0ģٿ'My��@2�\H�3@B�XJ�!?��<�@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@i����ٿR�l�b��@<��F��3@���P�!?e�j���@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@B�����ٿaxG50�@R���3@�y�<��!?5�z?��@�3���ٿ��IsS��@ ��(�3@���ꤐ!??*_��%�@�3���ٿ��IsS��@ ��(�3@���ꤐ!??*_��%�@�3���ٿ��IsS��@ ��(�3@���ꤐ!??*_��%�@�3���ٿ��IsS��@ ��(�3@���ꤐ!??*_��%�@�����ٿS=�:]��@fsqY��3@�䮴�!?�Bؠ���@�����ٿS=�:]��@fsqY��3@�䮴�!?�Bؠ���@�����ٿS=�:]��@fsqY��3@�䮴�!?�Bؠ���@�����ٿS=�:]��@fsqY��3@�䮴�!?�Bؠ���@C���ٿ#M7�]��@˒W���3@� 8���!?PQ��U��@C���ٿ#M7�]��@˒W���3@� 8���!?PQ��U��@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@a�d?Ţٿ�]J��l�@/�4P��3@�Ń��!?�=�$� �@C0�m��ٿ��B���@��^K��3@�DO0��!?䛄;��@C0�m��ٿ��B���@��^K��3@�DO0��!?䛄;��@C0�m��ٿ��B���@��^K��3@�DO0��!?䛄;��@C0�m��ٿ��B���@��^K��3@�DO0��!?䛄;��@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@If����ٿ4�H�@�/��3@#9���!?"�ئ�@�T���ٿ�1H�(�@ؖ��	�3@�R�u��!?o$�÷�@�T���ٿ�1H�(�@ؖ��	�3@�R�u��!?o$�÷�@����ٿ?��o���@J_�F�3@�:�k�!?��wR$$�@����ٿ?��o���@J_�F�3@�:�k�!?��wR$$�@�벙ٿ��)�ֺ�@�y����3@�CÐ!?�F&W�4�@�벙ٿ��)�ֺ�@�y����3@�CÐ!?�F&W�4�@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@C�r}�ٿ$>V�g��@m`(<�3@�̹�!?�i�_/��@\6P���ٿ���$.�@��jH�3@phH��!?��L���@�SA�ٿ���%$<�@�2y��3@~�9��!?�}c@��@�@�UW�ٿ�u�6��@�m���3@/[T�!?� �q���@�/"�<�ٿ������@����3@�2��!?��d�.��@�/"�<�ٿ������@����3@�2��!?��d�.��@���HI�ٿ�YD!1��@xлM��3@}Z��ݐ!?D���*�@���HI�ٿ�YD!1��@xлM��3@}Z��ݐ!?D���*�@�M�2�ٿm J|���@�[V'��3@������!?\���<�@"���v�ٿU���'�@#�)���3@��!?1~�{�@"���v�ٿU���'�@#�)���3@��!?1~�{�@"���v�ٿU���'�@#�)���3@��!?1~�{�@"���v�ٿU���'�@#�)���3@��!?1~�{�@ݗݬ��ٿ�ܚM��@Z�j�3@;�xՓ�!?����@(yR���ٿ�������@��o�w�3@=㙖�!?�C���Z�@(yR���ٿ�������@��o�w�3@=㙖�!?�C���Z�@(yR���ٿ�������@��o�w�3@=㙖�!?�C���Z�@��n��ٿ���V�R�@�7����3@-���!?=�;�f?�@��n��ٿ���V�R�@�7����3@-���!?=�;�f?�@��n��ٿ���V�R�@�7����3@-���!?=�;�f?�@��('��ٿ������@ݺ�J�3@u"�j��!?����M+�@��('��ٿ������@ݺ�J�3@u"�j��!?����M+�@��('��ٿ������@ݺ�J�3@u"�j��!?����M+�@��('��ٿ������@ݺ�J�3@u"�j��!?����M+�@c���ٿ���b�;�@�(H���3@�ؾ��!?�	0Re�@c���ٿ���b�;�@�(H���3@�ؾ��!?�	0Re�@c���ٿ���b�;�@�(H���3@�ؾ��!?�	0Re�@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@�jŘ~�ٿ~�%<��@|0��3@([�v��!?��ʀ,��@/�i���ٿ�$⪭��@3zgO��3@#4����!?t*h6�@/�i���ٿ�$⪭��@3zgO��3@#4����!?t*h6�@/�i���ٿ�$⪭��@3zgO��3@#4����!?t*h6�@/�i���ٿ�$⪭��@3zgO��3@#4����!?t*h6�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@�>����ٿ8�R=�@�!�@��3@�p4X��!?/ۋ�P�@;�� n�ٿtF��w��@�d���3@��'R��!?	Ӳ���@�M�W�ٿ\U�Df�@���G�3@ɣqb�!?��� ʫ�@n�C�5�ٿ����W�@W� ��3@%ik��!?��G�v�@n�C�5�ٿ����W�@W� ��3@%ik��!?��G�v�@n�C�5�ٿ����W�@W� ��3@%ik��!?��G�v�@�>y�Šٿ�웭�@:��ݲ�3@����Ð!?c�����@�~j�ٿ8e�_��@��V�m�3@g%@�!?UD� �E�@���̦�ٿt�}(EW�@_�e��3@[0	Һ�!?��+�n�@���̦�ٿt�}(EW�@_�e��3@[0	Һ�!?��+�n�@���̦�ٿt�}(EW�@_�e��3@[0	Һ�!?��+�n�@������ٿ,�l5���@�j.�%�3@�`��!?�9���@������ٿ,�l5���@�j.�%�3@�`��!?�9���@�eJ�9�ٿ�|;�M�@��@��3@S�'�!?��^����@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@ޮ��ٝٿQz����@4����3@�H���!?���G��@{ �٣�ٿ��4w��@��eV�3@}�a͐!?��6��@��,��ٿ�OL���@����3@�p���!?�ɠ)��@��,��ٿ�OL���@����3@�p���!?�ɠ)��@��,��ٿ�OL���@����3@�p���!?�ɠ)��@vp�Nߡٿ�r���j�@���o��3@>,DKː!?:fw��@vp�Nߡٿ�r���j�@���o��3@>,DKː!?:fw��@vp�Nߡٿ�r���j�@���o��3@>,DKː!?:fw��@vp�Nߡٿ�r���j�@���o��3@>,DKː!?:fw��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@�q4qОٿ����3�@p����3@W)�̐!?�q]@��@}�I,�ٿ/�N0���@6��R��3@N��3Ӑ!?�(�E��@}�I,�ٿ/�N0���@6��R��3@N��3Ӑ!?�(�E��@c�|z��ٿ�@�Zj��@�/js�3@�Y��!?�9�dT��@L]����ٿ��g�+��@�.:���3@A|�ѐ!?w( :���@L]����ٿ��g�+��@�.:���3@A|�ѐ!?w( :���@L]����ٿ��g�+��@�.:���3@A|�ѐ!?w( :���@��ճΤٿ�m�F���@�Ş���3@�.N�!?�,6�l��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@GفP��ٿ���k�W�@�?;_�3@�6�!?k8*��@ �_�P�ٿ����F�@��@���3@t�e�!?L�V��@ �_�P�ٿ����F�@��@���3@t�e�!?L�V��@ �_�P�ٿ����F�@��@���3@t�e�!?L�V��@87�բٿ���s���@�q&0��3@�%���!?����|�@87�բٿ���s���@�q&0��3@�%���!?����|�@87�բٿ���s���@�q&0��3@�%���!?����|�@�? ��ٿ�������@��?*��3@��ϐ!?N��=\��@�? ��ٿ�������@��?*��3@��ϐ!?N��=\��@�:ZF1�ٿ�&�ݲ~�@��Y��3@;!6˵�!?p�]��@�:ZF1�ٿ�&�ݲ~�@��Y��3@;!6˵�!?p�]��@�:ZF1�ٿ�&�ݲ~�@��Y��3@;!6˵�!?p�]��@�:ZF1�ٿ�&�ݲ~�@��Y��3@;!6˵�!?p�]��@�:ZF1�ٿ�&�ݲ~�@��Y��3@;!6˵�!?p�]��@D���'�ٿ<+�ͧ=�@�`j���3@���Ր!?گח���@D���'�ٿ<+�ͧ=�@�`j���3@���Ր!?گח���@D���'�ٿ<+�ͧ=�@�`j���3@���Ր!?گח���@sxIb#�ٿ�_r�%A�@�$!&b�3@�����!?���c��@ݾX��ٿ�<s�;E�@A_#ݬ�3@g���!?���j�@�5�
�ٿV7�%s��@�ױ��3@�)ܐ!?i�:����@�5�
�ٿV7�%s��@�ױ��3@�)ܐ!?i�:����@�5�
�ٿV7�%s��@�ױ��3@�)ܐ!?i�:����@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@�����ٿ7�o3#�@T�)��3@���ɐ!?���j܋�@��C�ٿ����0(�@�2�`�3@&�f��!?c�PY���@��C�ٿ����0(�@�2�`�3@&�f��!?c�PY���@� �ěٿ��6F���@�����3@�K�
��!?�O��51�@yꂁ�ٿ)�ۓ	�@�)�i#�3@�D[/�!?7���ȉ�@yꂁ�ٿ)�ۓ	�@�)�i#�3@�D[/�!?7���ȉ�@yꂁ�ٿ)�ۓ	�@�)�i#�3@�D[/�!?7���ȉ�@yꂁ�ٿ)�ۓ	�@�)�i#�3@�D[/�!?7���ȉ�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@����ٿ��8m�@;�Ha��3@Q]�6��!?~��b�@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@/��`��ٿ�8�7��@E�]�j�3@�˚I�!?� �̖��@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@��e���ٿW�
O �@������3@�\�ؐ!?B�\dY�@�Ȫ��ٿe����@�D�3@-wd��!?cu}I��@d.V�ٿ�o��0�@ϲ�I��3@�7*Y�!?XVYҝ��@d.V�ٿ�o��0�@ϲ�I��3@�7*Y�!?XVYҝ��@d����ٿg��)>��@�1����3@���_��!?��W��@��_no�ٿ�����i�@�T���3@&>�/��!?���	��@��3כٿ�����@� E@��3@�����!?������@��3כٿ�����@� E@��3@�����!?������@��3כٿ�����@� E@��3@�����!?������@ 9Ʈ��ٿ-��Uc�@!����3@v�wϐ!?׿��Q"�@���;�ٿ�=S*���@xe�@�4@
���|�!?%��%��@���;�ٿ�=S*���@xe�@�4@
���|�!?%��%��@�&J�ٿe~�#��@�[��& 4@����Y�!?CH4�3�@S��4]�ٿ�l����@2.��3@A��J��!?X���
�@S��4]�ٿ�l����@2.��3@A��J��!?X���
�@S��4]�ٿ�l����@2.��3@A��J��!?X���
�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@0�{K�ٿ�1\����@|nB�2�3@�1��!?��Lw�A�@�{xЦٿ@�m���@��Vk�3@Q%�2�!?���T
�@��>��ٿ��M �@L]g[��3@ ��~�!?��~� �@��>��ٿ��M �@L]g[��3@ ��~�!?��~� �@��>��ٿ��M �@L]g[��3@ ��~�!?��~� �@�N�N�ٿ �ȩ���@4v�t�3@;e�v�!?#���?�@]�� �ٿ����U�@���x�3@
�e���!?$��Z'<�@sެ��ٿ���R�@�)C��3@�s���!?ǡ	�cm�@sެ��ٿ���R�@�)C��3@�s���!?ǡ	�cm�@sެ��ٿ���R�@�)C��3@�s���!?ǡ	�cm�@sެ��ٿ���R�@�)C��3@�s���!?ǡ	�cm�@�%1��ٿ^J�Қ��@�]"}��3@ѲK0�!?۱� V�@�%1��ٿ^J�Қ��@�]"}��3@ѲK0�!?۱� V�@�%1��ٿ^J�Қ��@�]"}��3@ѲK0�!?۱� V�@��1��ٿ�h�~�u�@���`(�3@��NG�!?޻�"���@��1��ٿ�h�~�u�@���`(�3@��NG�!?޻�"���@��1��ٿ�h�~�u�@���`(�3@��NG�!?޻�"���@�X��y�ٿ		����@�����3@$͋���!?���� ��@�X��y�ٿ		����@�����3@$͋���!?���� ��@�X��y�ٿ		����@�����3@$͋���!?���� ��@�A=1�ٿa{�}��@�a�"��3@��m��!?�S����@�H���ٿ��'��@[��,�3@3RK�!?������@�H���ٿ��'��@[��,�3@3RK�!?������@�H���ٿ��'��@[��,�3@3RK�!?������@�H���ٿ��'��@[��,�3@3RK�!?������@�H���ٿ��'��@[��,�3@3RK�!?������@N����ٿ�u��[V�@)����3@��=d0�!? ߌ0�}�@N����ٿ�u��[V�@)����3@��=d0�!? ߌ0�}�@N����ٿ�u��[V�@)����3@��=d0�!? ߌ0�}�@N����ٿ�u��[V�@)����3@��=d0�!? ߌ0�}�@����ٿvْ���@������3@A%e�!?��/�Y�@����ٿvْ���@������3@A%e�!?��/�Y�@�[�f�ٿ!K:�~�@�>s!x�3@$]
�!?G�ܞR�@��Q���ٿ�]5lLS�@�� `��3@��"c
�!?$�l����@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@2���ٿ���T�@�K�z�3@��x�!?Ơ���#�@�mdn��ٿ���?���@�ژ��3@�OS�!?����C�@�mdn��ٿ���?���@�ژ��3@�OS�!?����C�@�mdn��ٿ���?���@�ژ��3@�OS�!?����C�@�mdn��ٿ���?���@�ژ��3@�OS�!?����C�@'�Fbȣٿ��^t
��@����3@B��e�!?�tC��]�@'�Fbȣٿ��^t
��@����3@B��e�!?�tC��]�@'�Fbȣٿ��^t
��@����3@B��e�!?�tC��]�@'�Fbȣٿ��^t
��@����3@B��e�!?�tC��]�@'�Fbȣٿ��^t
��@����3@B��e�!?�tC��]�@�)�`D�ٿs�w�@˱<���3@b��F��!?/&}h��@�)�`D�ٿs�w�@˱<���3@b��F��!?/&}h��@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�@�S�ٿ`�2�F��@��G���3@`��^��!?v��Jd�@�q�@�ٿ�T�&���@������3@F8�J��!?Dc*���@�q�@�ٿ�T�&���@������3@F8�J��!?Dc*���@����ٿZ��xY�@�"�3@{F�А!?a;�d�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@l�@R��ٿ�����@J7b7a�3@{'��ѐ!?*K�fk�@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@׈$<��ٿ1jgn��@2+�� 4@�[臐!?㸮i���@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@C!�V/�ٿ��&:"D�@��s���3@d���B�!?��׶A�@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@w���֠ٿ8M�`��@b��uw�3@�agϐ!?�/��@���l�ٿ������@�N����3@m�Y���!?fM)Y���@���l�ٿ������@�N����3@m�Y���!?fM)Y���@���l�ٿ������@�N����3@m�Y���!?fM)Y���@v�4��ٿ�G��@v#R~�3@Ӹ����!?ɒj@�K�@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@S�8?�ٿMYt�h�@�?1��3@c��^��!?z<�J��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@D�4T��ٿq`@U��@�3p1�3@�U���!?���|��@�h�Τٿ�pGkN�@������3@	{uPؐ!?�$���@�h�Τٿ�pGkN�@������3@	{uPؐ!?�$���@s?�(Z�ٿ��?�&�@������3@Ѐ��!?J�\L�@s?�(Z�ٿ��?�&�@������3@Ѐ��!?J�\L�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@�*�pޣٿ X=��"�@�М#�3@��fԐ!?�J�HN�@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@GC'tW�ٿ�(`�W��@�~�6�3@��J��!?'QXn��@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@И���ٿq���@l:�`�3@m�����!?M_B�ۥ�@9Ҩ(�ٿ[��@�1ͼ�3@�.TԨ�!?��V�5��@9Ҩ(�ٿ[��@�1ͼ�3@�.TԨ�!?��V�5��@�w>э�ٿU�M����@�+Hb�3@#��y�!?��>u�2�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@��C��ٿ%�b�@�/-9�3@�k*!!?s���"�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@����ٿ`}G��<�@�dV��3@P�����!?��7=�@\{�UE�ٿ�|v���@5 E��3@�B��Đ!?�;y�4�@�����ٿd��a�@�� ]��3@`�C��!?�N0ŽP�@�H�M��ٿX�!_���@vȤ�i�3@$П�А!?.`CB�@F�Z���ٿk���B��@ƌ`D�3@��u,�!?Oy��xT�@|�עٿ���R���@v�o�i�3@!$��̐!?ס0�5�@|�עٿ���R���@v�o�i�3@!$��̐!?ס0�5�@|�עٿ���R���@v�o�i�3@!$��̐!?ס0�5�@|�עٿ���R���@v�o�i�3@!$��̐!?ס0�5�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@�;(���ٿBUKK	��@swwe��3@��ѐ!?d��`aW�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@ҧ���ٿ=�3�b�@Uٴ{�3@�T���!?�ܤC*W�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�%t��ٿ������@��M?3�3@�Qs��!?$�94vM�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�:�Zx�ٿ��S����@k��.�3@�PV��!?�n�9/G�@�l�\�ٿ����Ύ�@�f���3@~<u�Ր!?�c�6Y�@�l�\�ٿ����Ύ�@�f���3@~<u�Ր!?�c�6Y�@�l�\�ٿ����Ύ�@�f���3@~<u�Ր!?�c�6Y�@�2|�ٿ~�Ф��@�3�I��3@]dk�А!?��6%��@�2|�ٿ~�Ф��@�3�I��3@]dk�А!?��6%��@�ns~~�ٿ�fK��@�n�$��3@�z
B��!?<�?�lp�@�ns~~�ٿ�fK��@�n�$��3@�z
B��!?<�?�lp�@�ns~~�ٿ�fK��@�n�$��3@�z
B��!?<�?�lp�@�ns~~�ٿ�fK��@�n�$��3@�z
B��!?<�?�lp�@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@@E\g��ٿ������@�s�M�3@0��ΐ!?-�:���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@���H�ٿ$�#��@Z����3@�*���!?+�E���@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@ԐZ)�ٿE����7�@��>�x�3@��FZ��!?0���u��@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@.�h�0�ٿ����K$�@�J�,�3@qO@�!?�Cw��u�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@_���ٿ�q8E���@]'�'��3@�/D�!?�n�s%�@˒�D�ٿ��r�J��@��}��3@D��ؐ!?�TKFi�@˒�D�ٿ��r�J��@��}��3@D��ؐ!?�TKFi�@˒�D�ٿ��r�J��@��}��3@D��ؐ!?�TKFi�@˒�D�ٿ��r�J��@��}��3@D��ؐ!?�TKFi�@˒�D�ٿ��r�J��@��}��3@D��ؐ!?�TKFi�@XČ8�ٿ�����@������3@�6�敖!?Ձ�֘�@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@����ٿʷ%��@�8�%7�3@���!?�Y(9��@�>����ٿ$���@vYV�3@+���!? �Q���@�>����ٿ$���@vYV�3@+���!? �Q���@�>����ٿ$���@vYV�3@+���!? �Q���@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�^����ٿ�����^�@����	�3@��~���!?����v-�@�Pi��ٿ(�V����@�V�KL�3@Z�3^�!?����m�@�Pi��ٿ(�V����@�V�KL�3@Z�3^�!?����m�@���.q�ٿDp،X.�@A�� J�3@���!?,����@�(%��ٿe�-!D��@�SN)2�3@�i��ǐ!?�+����@�(%��ٿe�-!D��@�SN)2�3@�i��ǐ!?�+����@��:}�ٿ:p~v0��@�v�tb�3@�ݫ㹐!?�J۬�l�@��:}�ٿ:p~v0��@�v�tb�3@�ݫ㹐!?�J۬�l�@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@t�Ao�ٿG����4�@�)FX4�3@��ა!?:'=����@�z/�¢ٿ��Ͻ�@�U5[L�3@/�ؐ!?�GR2
u�@�z/�¢ٿ��Ͻ�@�U5[L�3@/�ؐ!?�GR2
u�@�z/�¢ٿ��Ͻ�@�U5[L�3@/�ؐ!?�GR2
u�@��o"�ٿ�����@ ��L��3@Vbbz��!?h��*��@��o"�ٿ�����@ ��L��3@Vbbz��!?h��*��@��o"�ٿ�����@ ��L��3@Vbbz��!?h��*��@��o"�ٿ�����@ ��L��3@Vbbz��!?h��*��@��o"�ٿ�����@ ��L��3@Vbbz��!?h��*��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@Ѝ��f�ٿ��0j͜�@�T����3@�����!?��b��@ܓ�=��ٿ�U�͕��@�"��3@��[��!?O}�T��@ܓ�=��ٿ�U�͕��@�"��3@��[��!?O}�T��@ܓ�=��ٿ�U�͕��@�"��3@��[��!?O}�T��@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@�h��ٿI�gh
�@�A�MB�3@��z�ː!?���a�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@SYd�ٿ��-�?�@㻔���3@�d/Ȑ!?7�6F�R�@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�X�P@�ٿ@5_�'��@\`�e�3@�����!?���2/��@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�qt0\�ٿ,zRt�G�@����3@��3'��!?�˃0���@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�Q5g�ٿ�������@�ё�j�3@i4�T�!?��܉!�@�I(em�ٿ"F=����@]㕣 �3@{h���!?J?��n�@�I(em�ٿ"F=����@]㕣 �3@{h���!?J?��n�@�I(em�ٿ"F=����@]㕣 �3@{h���!?J?��n�@�I(em�ٿ"F=����@]㕣 �3@{h���!?J?��n�@��.�(�ٿc�ߋ��@��>k��3@)m%�!?�M,���@��.�(�ٿc�ߋ��@��>k��3@)m%�!?�M,���@/�4��ٿ�w�n��@q֗5�3@�bž�!?/��YT��@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@�����ٿ�gc3C��@b]�}�3@��Cɽ�!?��2���@����ٿʘ����@���3@9�̐!?�u�.S��@n.�I��ٿM�����@y�U���3@xD=IȐ!?s���v�@AT��ٿ#ȡ�(�@��]R�3@��A٪�!?a_�ؽ�@��*@��ٿx�E��@q
��	�3@�f�,d�!?Քۓ8�@��*@��ٿx�E��@q
��	�3@�f�,d�!?Քۓ8�@��*@��ٿx�E��@q
��	�3@�f�,d�!?Քۓ8�@��*@��ٿx�E��@q
��	�3@�f�,d�!?Քۓ8�@D�0�ٿ���ؗ�@?�,Y �3@��HAc�!?m����@D�0�ٿ���ؗ�@?�,Y �3@��HAc�!?m����@D�0�ٿ���ؗ�@?�,Y �3@��HAc�!?m����@D�0�ٿ���ؗ�@?�,Y �3@��HAc�!?m����@�:��>�ٿ'_�*�^�@��A�W�3@,n�3Ɛ!?�;�S��@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@s�1�G�ٿ_�;m'K�@&T�Kw�3@����ߐ!?K	Y Qs�@�& ���ٿ�-���@��
�3@v����!?��{�R��@�& ���ٿ�-���@��
�3@v����!?��{�R��@�& ���ٿ�-���@��
�3@v����!?��{�R��@�& ���ٿ�-���@��
�3@v����!?��{�R��@�& ���ٿ�-���@��
�3@v����!?��{�R��@�(�t�ٿ=
���A�@˴,�>�3@3����!?���^���@�3қٿZ�ZEݵ�@ ��`��3@X�Ð!?.��'B�@�rQ㧡ٿ��v��@�d[�E�3@B�t��!?�����;�@�rQ㧡ٿ��v��@�d[�E�3@B�t��!?�����;�@�rQ㧡ٿ��v��@�d[�E�3@B�t��!?�����;�@��$Y��ٿr<A����@ C��3@��cJ��!?�]J���@��$Y��ٿr<A����@ C��3@��cJ��!?�]J���@��$Y��ٿr<A����@ C��3@��cJ��!?�]J���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��,�.�ٿܶ�;�@�h��3@�j3��!?zW�t���@��p�դٿ��'�,�@+�y�&�3@{!���!?��uAP�@��p�դٿ��'�,�@+�y�&�3@{!���!?��uAP�@��p�դٿ��'�,�@+�y�&�3@{!���!?��uAP�@��p�դٿ��'�,�@+�y�&�3@{!���!?��uAP�@��ٙ�ٿ�ʶv��@R|�9u�3@�yC؛�!?�n�U��@��ٙ�ٿ�ʶv��@R|�9u�3@�yC؛�!?�n�U��@~�I��ٿ�'�,�U�@3 �4^�3@	3<_��!?�T�O>��@~�I��ٿ�'�,�U�@3 �4^�3@	3<_��!?�T�O>��@f��P�ٿG������@q����3@�"���!?�H�>���@f��P�ٿG������@q����3@�"���!?�H�>���@f��P�ٿG������@q����3@�"���!?�H�>���@f��P�ٿG������@q����3@�"���!?�H�>���@VovHn�ٿP�"~3�@����3@�й�!?�m�(F�@VovHn�ٿP�"~3�@����3@�й�!?�m�(F�@VovHn�ٿP�"~3�@����3@�й�!?�m�(F�@VovHn�ٿP�"~3�@����3@�й�!?�m�(F�@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@E4I��ٿXapAe�@�[�w�3@᭯���!?��`x���@��zW�ٿ��:0�@)�5���3@�A3���!?�����@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@��S�ٿ�������@o��?�3@�an�q�!?���T�@UEЀ�ٿ`�>S�A�@���3@��q�!?��.�,��@UEЀ�ٿ`�>S�A�@���3@��q�!?��.�,��@UEЀ�ٿ`�>S�A�@���3@��q�!?��.�,��@UEЀ�ٿ`�>S�A�@���3@��q�!?��.�,��@���=�ٿ�������@BhΌ<�3@̽��}�!?Q8ට��@���=�ٿ�������@BhΌ<�3@̽��}�!?Q8ට��@���=�ٿ�������@BhΌ<�3@̽��}�!?Q8ට��@���=�ٿ�������@BhΌ<�3@̽��}�!?Q8ට��@W��E�ٿ'�+�3��@��̻3�3@���!?��bW��@W��E�ٿ'�+�3��@��̻3�3@���!?��bW��@W��E�ٿ'�+�3��@��̻3�3@���!?��bW��@W��E�ٿ'�+�3��@��̻3�3@���!?��bW��@{z�8��ٿ��:�8�@B�2N?�3@���>�!?��>�D�@{z�8��ٿ��:�8�@B�2N?�3@���>�!?��>�D�@����ٿ����f�@%��6�3@��t�!?����^�@����ٿ����f�@%��6�3@��t�!?����^�@����ٿ����f�@%��6�3@��t�!?����^�@����ٿ����f�@%��6�3@��t�!?����^�@/�)�ԝٿ��n�r�@p����3@}�"&�!?���`�@/�)�ԝٿ��n�r�@p����3@}�"&�!?���`�@/�)�ԝٿ��n�r�@p����3@}�"&�!?���`�@/�)�ԝٿ��n�r�@p����3@}�"&�!?���`�@/�)�ԝٿ��n�r�@p����3@}�"&�!?���`�@�KJc�ٿ�&�9�@n�ˏ��3@����Ɛ!?����mU�@�KJc�ٿ�&�9�@n�ˏ��3@����Ɛ!?����mU�@�KJc�ٿ�&�9�@n�ˏ��3@����Ɛ!?����mU�@tzK퐨ٿ�F�����@��љ7�3@�_ps�!?ZX���l�@�U�:�ٿ�!����@�C�2��3@_�zMX�!?�H?TҨ�@"N<��ٿ�Vo�d��@"h�Y�3@�e��G�!?�of���@"N<��ٿ�Vo�d��@"h�Y�3@�e��G�!?�of���@"N<��ٿ�Vo�d��@"h�Y�3@�e��G�!?�of���@"N<��ٿ�Vo�d��@"h�Y�3@�e��G�!?�of���@"N<��ٿ�Vo�d��@"h�Y�3@�e��G�!?�of���@��_L�ٿ�m�72�@��	4�3@y�!?S��MK��@|�����ٿ�kS��[�@��G�3@QĽn�!?�Zj�l�@|�����ٿ�kS��[�@��G�3@QĽn�!?�Zj�l�@|�����ٿ�kS��[�@��G�3@QĽn�!?�Zj�l�@|�����ٿ�kS��[�@��G�3@QĽn�!?�Zj�l�@�(�F�ٿ���'�@2�p�j�3@.���!?��`1Ah�@�(�F�ٿ���'�@2�p�j�3@.���!?��`1Ah�@�(�F�ٿ���'�@2�p�j�3@.���!?��`1Ah�@�(�F�ٿ���'�@2�p�j�3@.���!?��`1Ah�@�(�F�ٿ���'�@2�p�j�3@.���!?��`1Ah�@]��ףٿa�h�Y�@<?���3@Wn��n�!?��Z���@]��ףٿa�h�Y�@<?���3@Wn��n�!?��Z���@]��ףٿa�h�Y�@<?���3@Wn��n�!?��Z���@�����ٿe^�$X�@5l#Av�3@��
Nv�!?|#{k��@�����ٿe^�$X�@5l#Av�3@��
Nv�!?|#{k��@�����ٿe^�$X�@5l#Av�3@��
Nv�!?|#{k��@�����ٿe^�$X�@5l#Av�3@��
Nv�!?|#{k��@�����ٿe^�$X�@5l#Av�3@��
Nv�!?|#{k��@7!;M�ٿBPu~S��@,v�ۑ�3@@��!?���)��@7!;M�ٿBPu~S��@,v�ۑ�3@@��!?���)��@7!;M�ٿBPu~S��@,v�ۑ�3@@��!?���)��@7!;M�ٿBPu~S��@,v�ۑ�3@@��!?���)��@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@�2�a�ٿ����z��@I~�bI�3@�]�X��!?U��~P�@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@D��	�ٿ�������@a"e��3@o[H׻�!?8�-���@=�_���ٿ��J����@�����3@�� E��!?��1���@=�_���ٿ��J����@�����3@�� E��!?��1���@=�_���ٿ��J����@�����3@�� E��!?��1���@5-�T��ٿ�E5���@������3@��S�!?Z��+��@5-�T��ٿ�E5���@������3@��S�!?Z��+��@5-�T��ٿ�E5���@������3@��S�!?Z��+��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@JĻ���ٿ2���m��@�L-Y��3@EK�w�!?�,G��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�y��&�ٿ�ƒ�@���`��3@aX���!?)�P��@�c�=�ٿ��~���@��Cd�3@�T!��!?�)'�e�@�c�=�ٿ��~���@��Cd�3@�T!��!?�)'�e�@�c�=�ٿ��~���@��Cd�3@�T!��!?�)'�e�@..�~3�ٿ@)�Y X�@v�^G=�3@��)���!?�p6�ߌ�@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@#d�t$�ٿ@���B��@���{�3@�(��!?Qq,����@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@�� ⪛ٿi}�O��@]3�ʺ�3@=r5��!?�ͺ$��@ms��ٿ��O~���@�t����3@c� GŐ!?�P0=��@ms��ٿ��O~���@�t����3@c� GŐ!?�P0=��@ms��ٿ��O~���@�t����3@c� GŐ!?�P0=��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@���ٿ���B��@��=]�3@.ɧ��!?xI��|��@O�+7.�ٿ,ۈE��@���f]�3@l�G�!?���,��@6c��ٿ�R�R�@CCl��3@�
����!?�D�G���@6c��ٿ�R�R�@CCl��3@�
����!?�D�G���@6c��ٿ�R�R�@CCl��3@�
����!?�D�G���@6c��ٿ�R�R�@CCl��3@�
����!?�D�G���@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@{ɡ�Ҟٿk��/�@�f����3@�*����!?�lU��@g����ٿL\e�;�@%-
��3@ᗐߐ!?�jK��@g����ٿL\e�;�@%-
��3@ᗐߐ!?�jK��@g����ٿL\e�;�@%-
��3@ᗐߐ!?�jK��@g����ٿL\e�;�@%-
��3@ᗐߐ!?�jK��@g����ٿL\e�;�@%-
��3@ᗐߐ!?�jK��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@ƀ��j�ٿ�:O��`�@	Pܧ�3@E 
4ܐ!?5��s��@�)�G��ٿ�+�\�;�@9�;�J�3@���Ǻ�!?��WP��@w
m�:�ٿ��V�Ff�@��Em�3@���h��!?�)
�r�@w
m�:�ٿ��V�Ff�@��Em�3@���h��!?�)
�r�@w
m�:�ٿ��V�Ff�@��Em�3@���h��!?�)
�r�@w
m�:�ٿ��V�Ff�@��Em�3@���h��!?�)
�r�@��$i8�ٿ�*c\��@�� \�3@/-ɐ�!?bA�j��@��$i8�ٿ�*c\��@�� \�3@/-ɐ�!?bA�j��@�\Vʣٿ�5�V���@���:�3@���!?�L��]�@,<�f��ٿg|&C�@�����3@�<)��!?i���@_%�^��ٿ(ch���@>o�;e�3@ёb�*�!?�,I�}��@_%�^��ٿ(ch���@>o�;e�3@ёb�*�!?�,I�}��@_%�^��ٿ(ch���@>o�;e�3@ёb�*�!?�,I�}��@.�byy�ٿ����D;�@�9	J!�3@J�F�o�!?d,�����@.�byy�ٿ����D;�@�9	J!�3@J�F�o�!?d,�����@.�byy�ٿ����D;�@�9	J!�3@J�F�o�!?d,�����@�RF�ٿ�3蹣�@�
U���3@�����!?�I��~�@�RF�ٿ�3蹣�@�
U���3@�����!?�I��~�@mˠ��ٿ=�����@f�k<c�3@�?�-�!? ����i�@mˠ��ٿ=�����@f�k<c�3@�?�-�!? ����i�@mˠ��ٿ=�����@f�k<c�3@�?�-�!? ����i�@mˠ��ٿ=�����@f�k<c�3@�?�-�!? ����i�@�s1�ٿ�c����@�o���3@�Y����!?�b��@�s1�ٿ�c����@�o���3@�Y����!?�b��@�s1�ٿ�c����@�o���3@�Y����!?�b��@�s1�ٿ�c����@�o���3@�Y����!?�b��@�s1�ٿ�c����@�o���3@�Y����!?�b��@�q���ٿ���<���@6��(�3@�5�.�!?���H�@ƞ$Y��ٿH��� ��@�W���3@����M�!?�T��$��@ƞ$Y��ٿH��� ��@�W���3@����M�!?�T��$��@ƞ$Y��ٿH��� ��@�W���3@����M�!?�T��$��@ƞ$Y��ٿH��� ��@�W���3@����M�!?�T��$��@ƞ$Y��ٿH��� ��@�W���3@����M�!?�T��$��@��Iԩٿ��b����@�[%��3@B����!?�Q��G�@'A�E�ٿ:	|����@/z�Cn�3@���HĐ!?G��y�@'A�E�ٿ:	|����@/z�Cn�3@���HĐ!?G��y�@'A�E�ٿ:	|����@/z�Cn�3@���HĐ!?G��y�@'A�E�ٿ:	|����@/z�Cn�3@���HĐ!?G��y�@'A�E�ٿ:	|����@/z�Cn�3@���HĐ!?G��y�@�&o*֪ٿe�ry"{�@�V�	�3@C��3��!?��|��@���
�ٿ�p���@יK��3@̲vs�!?et�e8�@���
�ٿ�p���@יK��3@̲vs�!?et�e8�@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@?�$�ٿ���z��@x�����3@Q�%��!?_ y���@�`~�3�ٿ��r%�@��:�H�3@?"�Ӑ!?��T^<�@�`~�3�ٿ��r%�@��:�H�3@?"�Ӑ!?��T^<�@�`~�3�ٿ��r%�@��:�H�3@?"�Ӑ!?��T^<�@�eP��ٿ���S���@/���u�3@�&��!?�3�t,�@�eP��ٿ���S���@/���u�3@�&��!?�3�t,�@���Z�ٿ�����@tqW�3@�>	��!?���5.r�@���Z�ٿ�����@tqW�3@�>	��!?���5.r�@���Z�ٿ�����@tqW�3@�>	��!?���5.r�@��-�ٿR̞\��@r9d��3@�l�cː!?���~@�@��-�ٿR̞\��@r9d��3@�l�cː!?���~@�@�KٿhI�+�R�@|���3@]ږN��!?AۚV[��@'ة�k�ٿh8g���@-,o��3@�����!?]M;����@'ة�k�ٿh8g���@-,o��3@�����!?]M;����@��C��ٿ���[�@v��l��3@@�5Y�!?^�r��	�@��C��ٿ���[�@v��l��3@@�5Y�!?^�r��	�@��C��ٿ���[�@v��l��3@@�5Y�!?^�r��	�@��C��ٿ���[�@v��l��3@@�5Y�!?^�r��	�@��C��ٿ���[�@v��l��3@@�5Y�!?^�r��	�@��7��ٿ�����@���|�3@0��z�!?��ߍ��@��7��ٿ�����@���|�3@0��z�!?��ߍ��@�Tj��ٿަ���@*���Q�3@|�j`�!?nw#�R"�@�Tj��ٿަ���@*���Q�3@|�j`�!?nw#�R"�@�Tj��ٿަ���@*���Q�3@|�j`�!?nw#�R"�@�Tj��ٿަ���@*���Q�3@|�j`�!?nw#�R"�@�Tj��ٿަ���@*���Q�3@|�j`�!?nw#�R"�@�K����ٿ�m�&��@\2. ��3@��*wu�!?&�٪L��@�K����ٿ�m�&��@\2. ��3@��*wu�!?&�٪L��@�K����ٿ�m�&��@\2. ��3@��*wu�!?&�٪L��@�<�թ�ٿ��g�~u�@�%_���3@���g��!?�� 6
W�@�<�թ�ٿ��g�~u�@�%_���3@���g��!?�� 6
W�@�<�թ�ٿ��g�~u�@�%_���3@���g��!?�� 6
W�@�<�թ�ٿ��g�~u�@�%_���3@���g��!?�� 6
W�@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@�(�p��ٿ%���k��@�~ s�3@iH��Đ!?Q�)��@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@]���ٿ��}xnK�@ϥ��3@��?��!?�M%z���@"#xݢٿ�0�̉d�@@gS#�3@)���!?��$m��@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@��t��ٿp���%�@�{�r�3@��Oߤ�!?ܣ� \�@������ٿ�H��%��@��+��3@3�u��!?�����L�@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@1��E�ٿN��Bt8�@�����3@��e��!?�M.���@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@lo�%ܡٿ�����l�@-��+�3@="	���!?���K`��@��� �ٿ��>�Q��@���S�3@��g���!?"�O/G��@��� �ٿ��>�Q��@���S�3@��g���!?"�O/G��@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@�z_�G�ٿ��2�@|%_g�3@�f˝�!?���@����f�ٿЋ�NP�@�V�\L�3@m���!?w/�C�[�@����f�ٿЋ�NP�@�V�\L�3@m���!?w/�C�[�@����f�ٿЋ�NP�@�V�\L�3@m���!?w/�C�[�@����f�ٿЋ�NP�@�V�\L�3@m���!?w/�C�[�@�.O��ٿ����Q�@�Q�M�3@H��#��!?J�w�@�.O��ٿ����Q�@�Q�M�3@H��#��!?J�w�@�.O��ٿ����Q�@�Q�M�3@H��#��!?J�w�@�.O��ٿ����Q�@�Q�M�3@H��#��!?J�w�@ۿ[g��ٿlscQ��@uQ{��3@�dn��!?�@Q����@ۿ[g��ٿlscQ��@uQ{��3@�dn��!?�@Q����@����ٿ=?�w{�@�Oʞ��3@u+���!?<0*�O�@����ٿ=?�w{�@�Oʞ��3@u+���!?<0*�O�@a�z/�ٿ}n�(�@.p��3@���d�!?fO*�L�@�)�.��ٿw��^	�@��Ŗ�3@S�(t�!?-��c�@���S��ٿ;Uf����@X���3@��m1��!?��lC+��@��*�ٿ�{�_���@�?G+!�3@�F&��!?}̭7�@RO���ٿa�q���@�L^b��3@Yf����!?Ԃ'��Y�@RO���ٿa�q���@�L^b��3@Yf����!?Ԃ'��Y�@RO���ٿa�q���@�L^b��3@Yf����!?Ԃ'��Y�@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@�#����ٿA޺��8�@(�]�3@pkQ�Ȑ!?_����@��ck��ٿC�1���@�x��3@%����!?���4��@��ck��ٿC�1���@�x��3@%����!?���4��@��f_<�ٿAy1g`��@k5�s�3@�OW&Ő!? �%��@��f_<�ٿAy1g`��@k5�s�3@�OW&Ő!? �%��@��f_<�ٿAy1g`��@k5�s�3@�OW&Ő!? �%��@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@_��zg�ٿ�A�|��@+ ��J�3@�f0�ې!?y������@6ԏ��ٿ)������@:T����3@/0�[H�!?��~� �@rz�\�ٿ)?�F\�@�0E�3@d�Z�!?��0���@rz�\�ٿ)?�F\�@�0E�3@d�Z�!?��0���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�'K>��ٿΕ�F���@��%��3@�<y�!?[n���@�ٶ�r�ٿ���R�@�QӠ�3@��Q��!?K� ���@�ٶ�r�ٿ���R�@�QӠ�3@��Q��!?K� ���@�ٶ�r�ٿ���R�@�QӠ�3@��Q��!?K� ���@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�7A�ٿW}H҈��@G�[�3@ɟ~"�!?d��9b�@�/׵ݠٿ�nM���@�ܻ���3@��\� �!?�����@�/׵ݠٿ�nM���@�ܻ���3@��\� �!?�����@���绦ٿ��a�8��@6n���3@�7.��!?��2{��@���绦ٿ��a�8��@6n���3@�7.��!?��2{��@��š��ٿd�tZ���@��˹"�3@�lײ�!?e>~z��@��o�~�ٿ~�S6\�@@y�ɏ�3@&M̵�!?���z�@��o�~�ٿ~�S6\�@@y�ɏ�3@&M̵�!?���z�@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@�ӏ�!�ٿ'�o�"�@���A]�3@G1sEА!?���y���@^�Q��ٿ��>�t	�@�Y���3@��M[ɐ!?]�0{�r�@^�Q��ٿ��>�t	�@�Y���3@��M[ɐ!?]�0{�r�@^�Q��ٿ��>�t	�@�Y���3@��M[ɐ!?]�0{�r�@^�Q��ٿ��>�t	�@�Y���3@��M[ɐ!?]�0{�r�@����+�ٿ�� �n��@I1p�7�3@ �W��!?��0�v0�@����+�ٿ�� �n��@I1p�7�3@ �W��!?��0�v0�@B!��|�ٿ��W��@�G�;��3@����!?,2���c�@B!��|�ٿ��W��@�G�;��3@����!?,2���c�@B!��|�ٿ��W��@�G�;��3@����!?,2���c�@B!��|�ٿ��W��@�G�;��3@����!?,2���c�@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@��麞ٿ4�K�3�@N˚a�3@E��ߐ!?y���4��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@t���S�ٿ�mH�#�@q�s���3@%�Ǚ�!?b��J��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@N�B�]�ٿT.��Wg�@U�k�3@�%����!?���,��@��m�ٿt���a��@��/�/�3@m�[��!?
.0O�Q�@��m�ٿt���a��@��/�/�3@m�[��!?
.0O�Q�@��m�ٿt���a��@��/�/�3@m�[��!?
.0O�Q�@��m�ٿt���a��@��/�/�3@m�[��!?
.0O�Q�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@����P�ٿ¦�G�G�@:��|^�3@j��ǐ!?���=�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�<���ٿ��j(+��@z��3@c�*E��!?Ҡ<XS�@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�3��*�ٿ<oG�_R�@yM��3�3@w�nUk�!?M|�v��@�\���ٿ٥����@2�|Av�3@� d͐!?�^y�@�\���ٿ٥����@2�|Av�3@� d͐!?�^y�@�\���ٿ٥����@2�|Av�3@� d͐!?�^y�@�\���ٿ٥����@2�|Av�3@� d͐!?�^y�@�\���ٿ٥����@2�|Av�3@� d͐!?�^y�@��3��ٿM&�d�i�@W�|h-�3@��Zr��!?Ǥ�K��@��3��ٿM&�d�i�@W�|h-�3@��Zr��!?Ǥ�K��@�O�Ѣٿ~-��%��@�]�Q6�3@�ϞdՐ!?�b~�%�@�O�Ѣٿ~-��%��@�]�Q6�3@�ϞdՐ!?�b~�%�@�O�Ѣٿ~-��%��@�]�Q6�3@�ϞdՐ!?�b~�%�@%���ٿ*.�����@|�6���3@u�~Ґ!?e�����@%���ٿ*.�����@|�6���3@u�~Ґ!?e�����@%���ٿ*.�����@|�6���3@u�~Ґ!?e�����@��'=��ٿG#�%#�@^ �3@fs�q֐!?��)�@��'=��ٿG#�%#�@^ �3@fs�q֐!?��)�@��'=��ٿG#�%#�@^ �3@fs�q֐!?��)�@��'=��ٿG#�%#�@^ �3@fs�q֐!?��)�@[G�r��ٿ�RGq��@l�,?��3@m����!?.�z�Q-�@[G�r��ٿ�RGq��@l�,?��3@m����!?.�z�Q-�@[G�r��ٿ�RGq��@l�,?��3@m����!?.�z�Q-�@�u�ky�ٿ��s�e��@wq��3@]w���!?�ma��@�u�ky�ٿ��s�e��@wq��3@]w���!?�ma��@K��"��ٿ9�/���@y�(�3@d�&���!?#c�D��@K��"��ٿ9�/���@y�(�3@d�&���!?#c�D��@K��"��ٿ9�/���@y�(�3@d�&���!?#c�D��@K��"��ٿ9�/���@y�(�3@d�&���!?#c�D��@K��"��ٿ9�/���@y�(�3@d�&���!?#c�D��@u!!2�ٿlvU�f��@��ٲ��3@'����!?�d%3#��@���Ɯٿ-�d�l��@����6�3@��o��!??̉�y��@���Ɯٿ-�d�l��@����6�3@��o��!??̉�y��@���Ɯٿ-�d�l��@����6�3@��o��!??̉�y��@a����ٿ�6�ܨ�@C{�T��3@�Y_��!?/ª���@�J�M��ٿ��q}��@n��x�3@mӕr�!?%�@brq�@�J�M��ٿ��q}��@n��x�3@mӕr�!?%�@brq�@�J�M��ٿ��q}��@n��x�3@mӕr�!?%�@brq�@~�쮥ٿ�6i]��@1*h���3@��N�!?���,�D�@~�쮥ٿ�6i]��@1*h���3@��N�!?���,�D�@���c�ٿ�������@u�ߞ�3@wqb�ߐ!??��$��@���c�ٿ�������@u�ߞ�3@wqb�ߐ!??��$��@:3ߠ�ٿ�
�c�]�@��d ��3@k
Ce��!?��:;_�@tw/4��ٿ�v�����@���ϣ�3@�ڂ\��!?Xw��j�@tw/4��ٿ�v�����@���ϣ�3@�ڂ\��!?Xw��j�@tw/4��ٿ�v�����@���ϣ�3@�ڂ\��!?Xw��j�@tw/4��ٿ�v�����@���ϣ�3@�ڂ\��!?Xw��j�@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@��ZE��ٿ4~9�7��@�>�[�3@�5��!?�;���@}Zg��ٿs����@�}�,�3@��v��!?������@}Zg��ٿs����@�}�,�3@��v��!?������@}Zg��ٿs����@�}�,�3@��v��!?������@"!��2�ٿ�FT���@��jP��3@��ֿ��!?��G6��@���c�ٿ#�%$��@Ce�k�3@���|�!?������@���c�ٿ#�%$��@Ce�k�3@���|�!?������@�ؗ.��ٿ�|F$��@�����3@��G�m�!?����vu�@�ؗ.��ٿ�|F$��@�����3@��G�m�!?����vu�@��0�	�ٿ�t�c �@�j���3@�\���!?�r���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@E�����ٿ�A��@p82[!�3@��=��!?��f
���@#�DX��ٿ#y�i��@PcV�(�3@��T�Ð!?I�Fl�I�@#�DX��ٿ#y�i��@PcV�(�3@��T�Ð!?I�Fl�I�@#�DX��ٿ#y�i��@PcV�(�3@��T�Ð!?I�Fl�I�@#�DX��ٿ#y�i��@PcV�(�3@��T�Ð!?I�Fl�I�@#�DX��ٿ#y�i��@PcV�(�3@��T�Ð!?I�Fl�I�@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@�����ٿ�k�k��@4>S��3@!�!Ő!?ـ�C��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@:�9��ٿ*����@B�t���3@.�����!?��0((��@�c�<Ԟٿ�d����@t��- 4@��u���!?�6�o�f�@�c�<Ԟٿ�d����@t��- 4@��u���!?�6�o�f�@�ܙ���ٿE�]}��@��/4@���!?h�K@$��@�ܙ���ٿE�]}��@��/4@���!?h�K@$��@�ܙ���ٿE�]}��@��/4@���!?h�K@$��@�ܙ���ٿE�]}��@��/4@���!?h�K@$��@5��Q�ٿ�9M�@R�ӝ4@z�,t&�!?H���-�@_�4l�ٿ�50��@k}E�4@z��!�!?&A���$�@_�4l�ٿ�50��@k}E�4@z��!�!?&A���$�@�FRF�ٿ� �/��@XH�R�3@����!?�x?8���@�FRF�ٿ� �/��@XH�R�3@����!?�x?8���@��OT[�ٿ�<�#�@������3@i�b��!?��a�!��@��OT[�ٿ�<�#�@������3@i�b��!?��a�!��@��OT[�ٿ�<�#�@������3@i�b��!?��a�!��@� �ࠥٿ��Y~�_�@�.NN��3@+���4�!?�V;@�l�@� �ࠥٿ��Y~�_�@�.NN��3@+���4�!?�V;@�l�@� �ࠥٿ��Y~�_�@�.NN��3@+���4�!?�V;@�l�@� �ࠥٿ��Y~�_�@�.NN��3@+���4�!?�V;@�l�@� �ࠥٿ��Y~�_�@�.NN��3@+���4�!?�V;@�l�@{��
�ٿ�@-2���@۠5��3@��g䜐!?َ�Y�@�����ٿ�}
4Z�@�ͺ��3@^�ѻ�!?�2#���@�����ٿ�}
4Z�@�ͺ��3@^�ѻ�!?�2#���@���̣ٿ��1��@\n��3@�	�΂�!?����a�@���̣ٿ��1��@\n��3@�	�΂�!?����a�@���̣ٿ��1��@\n��3@�	�΂�!?����a�@L&4G��ٿ}�'o1n�@O9� �3@���̐!?վ4�i��@���1٤ٿ]�SMa�@8����3@"J�Ȑ!?Kj�GA�@���1٤ٿ]�SMa�@8����3@"J�Ȑ!?Kj�GA�@���1٤ٿ]�SMa�@8����3@"J�Ȑ!?Kj�GA�@���1٤ٿ]�SMa�@8����3@"J�Ȑ!?Kj�GA�@�[��_�ٿ��L���@����3@ˮCf�!?�'�$	�@�[��_�ٿ��L���@����3@ˮCf�!?�'�$	�@�[��_�ٿ��L���@����3@ˮCf�!?�'�$	�@�[��_�ٿ��L���@����3@ˮCf�!?�'�$	�@�[��_�ٿ��L���@����3@ˮCf�!?�'�$	�@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@%�M5�ٿ3%��e��@���� �3@�퓐!?V�;���@O�(m��ٿQ� -��@4j�\3�3@������!?�!�'V�@O�(m��ٿQ� -��@4j�\3�3@������!?�!�'V�@O�(m��ٿQ� -��@4j�\3�3@������!?�!�'V�@O�(m��ٿQ� -��@4j�\3�3@������!?�!�'V�@����/�ٿ��j��@�6]v�3@e�nΐ!??G�0
t�@����/�ٿ��j��@�6]v�3@e�nΐ!??G�0
t�@����/�ٿ��j��@�6]v�3@e�nΐ!??G�0
t�@si�H�ٿ�?m�K�@lԌ��3@[�ӧ��!?�+��+&�@si�H�ٿ�?m�K�@lԌ��3@[�ӧ��!?�+��+&�@si�H�ٿ�?m�K�@lԌ��3@[�ӧ��!?�+��+&�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@�wG�Τٿ��j&�.�@ݺ&���3@�����!?�'rCY�@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@}�XHM�ٿ�R|���@���C��3@-���!?�Nv��@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@�q��ٿ�m�Ӊ��@�����3@��
�!??7���@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@��l��ٿ�a5�-�@�|V�'�3@<�w�!?���Q��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@�ax\�ٿ��9ɣ��@�UiN��3@�ۈ��!?M�T�y��@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��<���ٿ�/�`���@����3@6�r`ΐ!?�\Ih���@��iĬ�ٿ������@�!�g��3@#����!?#�W�$��@��iĬ�ٿ������@�!�g��3@#����!?#�W�$��@!.GX`�ٿ-p���@�����3@��E�!?.����@!.GX`�ٿ-p���@�����3@��E�!?.����@!.GX`�ٿ-p���@�����3@��E�!?.����@!.GX`�ٿ-p���@�����3@��E�!?.����@!.GX`�ٿ-p���@�����3@��E�!?.����@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@i��7Ȝٿ3X�/��@���a��3@s;��!?�@3h�/�@�_u(�ٿ�6����@^���3@V.2"��!?�%��<?�@�_u(�ٿ�6����@^���3@V.2"��!?�%��<?�@�_u(�ٿ�6����@^���3@V.2"��!?�%��<?�@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��B�ٿB@�T\��@U/#�E�3@�=�fÐ!?(�mؚ��@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@��Ajǡٿ����yH�@<玃r�3@E��%�!?�R���@�s旚ٿUՙ�
�@���	8�3@�>P�!?��1���@�@x�E�ٿ}%Ϛ�}�@��%@�3@q�e|�!?�NX���@��Ѻ��ٿ����@����3@�zs���!?��
t^��@��Ѻ��ٿ����@����3@�zs���!?��
t^��@�{ȸ�ٿ�E�ci�@���f�3@��MJi�!??zj�n�@S}�;�ٿ���'��@=θD�3@u�Fu�!?#6^��=�@S}�;�ٿ���'��@=θD�3@u�Fu�!?#6^��=�@S}�;�ٿ���'��@=θD�3@u�Fu�!?#6^��=�@S}�;�ٿ���'��@=θD�3@u�Fu�!?#6^��=�@S}�;�ٿ���'��@=θD�3@u�Fu�!?#6^��=�@X#L͟ٿ������@V�1�X�3@�<7w�!?��8��@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@`�q5�ٿ:�9�@�h�Z�3@G�E���!?�=8�
y�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@\�L�ϛٿ��i.�+�@�>� ��3@��η�!?��/�f>�@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@��@璝ٿ5%{G ��@�G����3@DFbp��!?�(,=��@vY���ٿ�l�����@�[��3@��^�Ð!?t&��t��@���n��ٿ���r���@�-d���3@>C�Đ!?{B4|��@���n��ٿ���r���@�-d���3@>C�Đ!?{B4|��@���n��ٿ���r���@�-d���3@>C�Đ!?{B4|��@���n��ٿ���r���@�-d���3@>C�Đ!?{B4|��@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�ɴZ�ٿ�i��H�@˕����3@�zYm�!?q\>�a�@�[/�N�ٿ/>�j��@Y�i�3@[��̐!?Й �j�@�[/�N�ٿ/>�j��@Y�i�3@[��̐!?Й �j�@�[/�N�ٿ/>�j��@Y�i�3@[��̐!?Й �j�@�[/�N�ٿ/>�j��@Y�i�3@[��̐!?Й �j�@�C����ٿ2ve��@%�:~�3@kRܤ��!?Z���N�@�C����ٿ2ve��@%�:~�3@kRܤ��!?Z���N�@�C����ٿ2ve��@%�:~�3@kRܤ��!?Z���N�@�C����ٿ2ve��@%�:~�3@kRܤ��!?Z���N�@�C����ٿ2ve��@%�:~�3@kRܤ��!?Z���N�@��vm�ٿ����@�hQC��3@��al��!?K&�i�@��vm�ٿ����@�hQC��3@��al��!?K&�i�@��vm�ٿ����@�hQC��3@��al��!?K&�i�@��vm�ٿ����@�hQC��3@��al��!?K&�i�@��vm�ٿ����@�hQC��3@��al��!?K&�i�@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@r��f��ٿoC�e+��@F�Cb�3@�����!?�Q����@�_x�)�ٿ�B��8'�@�ك1�3@��r�Ɛ!?��o�?��@�v�L3�ٿ��^�H��@�=�o�3@��&�ِ!?�<����@&�0���ٿd)���;�@���!�3@���U��!?Tq��W�@&�0���ٿd)���;�@���!�3@���U��!?Tq��W�@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@����ٿ;�d[���@m��O�3@�V�`��!?�(F#��@�Q���ٿ�g��>�@M��c��3@��-ڐ!?�-}�A�@�Q���ٿ�g��>�@M��c��3@��-ڐ!?�-}�A�@���6��ٿ�Z���D�@��r��3@�ד�ؐ!?}��i�@���6��ٿ�Z���D�@��r��3@�ד�ؐ!?}��i�@���6��ٿ�Z���D�@��r��3@�ד�ؐ!?}��i�@`����ٿ�]�����@gj����3@�2o��!?t�o��}�@`����ٿ�]�����@gj����3@�2o��!?t�o��}�@`����ٿ�]�����@gj����3@�2o��!?t�o��}�@`����ٿ�]�����@gj����3@�2o��!?t�o��}�@-�F	��ٿ�F=!��@�ɹ�3@10�8�!?6��^Z��@��H�;�ٿ��[�g�@��c�3@z?s��!?(�a!���@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�h��L�ٿA55���@�	[�3@��Į��!?j�
����@�-���ٿΘ:lk�@��(%��3@����!?ց��c��@�-���ٿΘ:lk�@��(%��3@����!?ց��c��@`ݨ���ٿ�m�	�@Wb��3@�
�ݵ�!?Ά0��@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@{���ٿY�Mܲ5�@��H�(�3@ϯh���!?S���@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@vj6/ �ٿ� ��Y�@��|�V�3@�!+��!?�|�G��@e��{�ٿf���9��@NږK��3@�lS2�!?X�ޛ���@e��{�ٿf���9��@NږK��3@�lS2�!?X�ޛ���@e��{�ٿf���9��@NږK��3@�lS2�!?X�ޛ���@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@U���ٿz�h���@�fy �3@�Jf��!?)~��A�@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@��m{c�ٿVYc/��@�JƟ��3@����!?v��"��@~�T�ٿ�dô��@����o�3@�����!?l
�%���@~�T�ٿ�dô��@����o�3@�����!?l
�%���@�|դٿ����4�@�G�V��3@��$2ؐ!?T�,��@�����ٿCe�Qn�@F�S�Q�3@�-�ː!?���<��@�����ٿCe�Qn�@F�S�Q�3@�-�ː!?���<��@�����ٿCe�Qn�@F�S�Q�3@�-�ː!?���<��@�����ٿCe�Qn�@F�S�Q�3@�-�ː!?���<��@�����ٿCe�Qn�@F�S�Q�3@�-�ː!?���<��@E�O|�ٿ�n�j�u�@�&�z(�3@a����!?����@E�O|�ٿ�n�j�u�@�&�z(�3@a����!?����@E�O|�ٿ�n�j�u�@�&�z(�3@a����!?����@$f䆦ٿG�,xuN�@���C��3@X8�!?��Sr��@`�YH��ٿ6�+#���@������3@#�|�!?��][R�@��*,��ٿӷ&0W��@bTLo�3@������!?_4�w�@;�Ic�ٿ��OMi��@��~(��3@eYޥ�!?�O���[�@;�Ic�ٿ��OMi��@��~(��3@eYޥ�!?�O���[�@;�Ic�ٿ��OMi��@��~(��3@eYޥ�!?�O���[�@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@c�?�	�ٿ"l�![�@�c����3@��`ɰ�!?�B�%���@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�i0�=�ٿ(�]�X�@�
����3@6��f��!?T�%0�@�a�4_�ٿ���!���@�[�u��3@7O�Ő!?vb���@�a�4_�ٿ���!���@�[�u��3@7O�Ő!?vb���@�a�4_�ٿ���!���@�[�u��3@7O�Ő!?vb���@�a�4_�ٿ���!���@�[�u��3@7O�Ő!?vb���@�a�4_�ٿ���!���@�[�u��3@7O�Ő!?vb���@gv�>�ٿ(q��U�@O;K��3@q몆��!?�,.��@gv�>�ٿ(q��U�@O;K��3@q몆��!?�,.��@gv�>�ٿ(q��U�@O;K��3@q몆��!?�,.��@gv�>�ٿ(q��U�@O;K��3@q몆��!?�,.��@gv�>�ٿ(q��U�@O;K��3@q몆��!?�,.��@#̼y�ٿ1�eI�@�Ę��3@#�Uא!?�l/��@#̼y�ٿ1�eI�@�Ę��3@#�Uא!?�l/��@#̼y�ٿ1�eI�@�Ę��3@#�Uא!?�l/��@#̼y�ٿ1�eI�@�Ę��3@#�Uא!?�l/��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@�5$>�ٿ�mo�p��@窢���3@U�>��!?���=Y��@ӠǠ͝ٿ#W~���@M�Nd��3@__&Hڐ!?�X$x���@#�<�S�ٿ�UQZ|.�@A�,^��3@+�ː!?7p�W�@��)�ٿM�1�S�@����g�3@���h�!?�^�x��@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@�~b�ߝٿ�ٝ��F�@�oH�3@2����!?M̸���@L��^�ٿ�E�pAI�@[����3@�\!<��!?��:��@L��^�ٿ�E�pAI�@[����3@�\!<��!?��:��@o��i��ٿ]bZ_��@��ӫ��3@πW��!?CKE�I��@���ڦٿ2M���@R�6�!�3@?�|\��!?��/L��@�-B촡ٿ�UO���@V>�W��3@���!?/:�`��@�-B촡ٿ�UO���@V>�W��3@���!?/:�`��@�-B촡ٿ�UO���@V>�W��3@���!?/:�`��@�-B촡ٿ�UO���@V>�W��3@���!?/:�`��@�-B촡ٿ�UO���@V>�W��3@���!?/:�`��@�m�&ȥٿ2ܓ�6�@�&o���3@�H���!?O�W���@�m�&ȥٿ2ܓ�6�@�&o���3@�H���!?O�W���@�UПٿ| M�_��@�3(4�3@� �H�!?��['�u�@�UПٿ| M�_��@�3(4�3@� �H�!?��['�u�@n	h3śٿ�����%�@ !����3@T�E�!?F|�K|i�@n	h3śٿ�����%�@ !����3@T�E�!?F|�K|i�@n	h3śٿ�����%�@ !����3@T�E�!?F|�K|i�@n	h3śٿ�����%�@ !����3@T�E�!?F|�K|i�@HѳWx�ٿ!_�f�@hȸ��3@v>@���!?{B_X�T�@HѳWx�ٿ!_�f�@hȸ��3@v>@���!?{B_X�T�@HѳWx�ٿ!_�f�@hȸ��3@v>@���!?{B_X�T�@S-�6��ٿ<JS���@��4h��3@A.n�ǐ!?%���@S-�6��ٿ<JS���@��4h��3@A.n�ǐ!?%���@S-�6��ٿ<JS���@��4h��3@A.n�ǐ!?%���@S-�6��ٿ<JS���@��4h��3@A.n�ǐ!?%���@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@�W�̙ٿ���p��@�����3@6� Đ!?�t���1�@zo&��ٿA�8���@��?ap�3@��I��!?��pv��@zo&��ٿA�8���@��?ap�3@��I��!?��pv��@zo&��ٿA�8���@��?ap�3@��I��!?��pv��@zo&��ٿA�8���@��?ap�3@��I��!?��pv��@�
��ٿC��1���@W3�}E�3@Ն31�!?PݹX�@�
��ٿC��1���@W3�}E�3@Ն31�!?PݹX�@�
��ٿC��1���@W3�}E�3@Ն31�!?PݹX�@�
��ٿC��1���@W3�}E�3@Ն31�!?PݹX�@�
��ٿC��1���@W3�}E�3@Ն31�!?PݹX�@\���k�ٿ�|�c��@X"&a��3@�o-���!?Ņ%��@\���k�ٿ�|�c��@X"&a��3@�o-���!?Ņ%��@\���k�ٿ�|�c��@X"&a��3@�o-���!?Ņ%��@\���k�ٿ�|�c��@X"&a��3@�o-���!?Ņ%��@s~����ٿ2e�����@ˀA=��3@��.��!?/��� �@s~����ٿ2e�����@ˀA=��3@��.��!?/��� �@�cY`	�ٿS/D0X0�@\YCz�3@%B/i��!?E�F�3��@�cY`	�ٿS/D0X0�@\YCz�3@%B/i��!?E�F�3��@�cY`	�ٿS/D0X0�@\YCz�3@%B/i��!?E�F�3��@�cY`	�ٿS/D0X0�@\YCz�3@%B/i��!?E�F�3��@�g��c�ٿ·���v�@˵��3@��Í��!?�jD��@�w1�)�ٿ"��m�@aG7��3@�0���!?�»9'�@�w1�)�ٿ"��m�@aG7��3@�0���!?�»9'�@�w1�)�ٿ"��m�@aG7��3@�0���!?�»9'�@�w1�)�ٿ"��m�@aG7��3@�0���!?�»9'�@�w1�)�ٿ"��m�@aG7��3@�0���!?�»9'�@��U�ٿ��i"��@�v���3@7��;ː!?V�2yq�@��U�ٿ��i"��@�v���3@7��;ː!?V�2yq�@��U�ٿ��i"��@�v���3@7��;ː!?V�2yq�@6h�g4�ٿ[w�Vw�@>�1cx�3@`�X�̐!?�[0�p�@f+����ٿ������@t?�:|�3@���O�!?�8�-C�@o��r�ٿ ��6���@�m�3�3@��u�!?8l�orA�@o��r�ٿ ��6���@�m�3�3@��u�!?8l�orA�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@B ᓴ�ٿ̣kz�?�@P���v�3@Y���!?6*�F9X�@���	*�ٿ%��k���@ߴT�H�3@Sqڷ�!?l�Q���@���	*�ٿ%��k���@ߴT�H�3@Sqڷ�!?l�Q���@��k"�ٿa��*`��@���w4�3@�tx��!?O�����@蘅��ٿ�o=9�-�@�+�}�3@��p���!?BM���@蘅��ٿ�o=9�-�@�+�}�3@��p���!?BM���@蘅��ٿ�o=9�-�@�+�}�3@��p���!?BM���@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@(~JT�ٿTV�����@:ݣ��3@�K\c��!?�Vϳf�@8O� Τٿ1�Bc9��@A�^K�3@�[�M|�!?�K�2�@�����ٿ���f�@�4��3@^���!?}�0�ė�@�����ٿ���f�@�4��3@^���!?}�0�ė�@�����ٿ���f�@�4��3@^���!?}�0�ė�@�����ٿ���f�@�4��3@^���!?}�0�ė�@�����ٿ���f�@�4��3@^���!?}�0�ė�@�����ٿ���f�@�4��3@^���!?}�0�ė�@f����ٿ�'��x�@��)�3@S%ePؐ!?mH�d���@f����ٿ�'��x�@��)�3@S%ePؐ!?mH�d���@,J�㐤ٿe"Qړ'�@?�Q?]�3@B;�!?�s>c$�@,J�㐤ٿe"Qړ'�@?�Q?]�3@B;�!?�s>c$�@�A��<�ٿ���/]$�@p{����3@�~��!?�p����@�A��<�ٿ���/]$�@p{����3@�~��!?�p����@��Ԕ�ٿ\�ʥ��@�Y�#7�3@��*А!?�rڶ�	�@��Ԕ�ٿ\�ʥ��@�Y�#7�3@��*А!?�rڶ�	�@��|=�ٿ����g��@�P+�J�3@`�P���!?�fc_eK�@��|=�ٿ����g��@�P+�J�3@`�P���!?�fc_eK�@V5�ٝٿ�O|� ��@�=��3@_0_���!?�}��@V5�ٝٿ�O|� ��@�=��3@_0_���!?�}��@S`n�ٿRe��BC�@�I���3@/� ��!?���x��@S`n�ٿRe��BC�@�I���3@/� ��!?���x��@S`n�ٿRe��BC�@�I���3@/� ��!?���x��@S`n�ٿRe��BC�@�I���3@/� ��!?���x��@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@���Ϝٿ�\Wn"R�@�8x�K�3@�-��!?7�h
�)�@�s��
�ٿ��ɐ�@�W|���3@�����!?������@�s��
�ٿ��ɐ�@�W|���3@�����!?������@�s��
�ٿ��ɐ�@�W|���3@�����!?������@��=엟ٿ�	g�	��@M����3@5L��!?�a��n��@��=엟ٿ�	g�	��@M����3@5L��!?�a��n��@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@����N�ٿ�m2Q� �@�&����3@����!?�a?�[J�@�#��̞ٿ��$�Q\�@�l���3@P�#ސ!?.X���@�#��̞ٿ��$�Q\�@�l���3@P�#ސ!?.X���@�#��̞ٿ��$�Q\�@�l���3@P�#ސ!?.X���@�#��̞ٿ��$�Q\�@�l���3@P�#ސ!?.X���@D�4�ٟٿנ�.m�@
K���3@���ݐ!?���|�@D�4�ٟٿנ�.m�@
K���3@���ݐ!?���|�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@f��D�ٿ��	�}�@#yX��3@]�P{�!?^rL!�@'����ٿ^N��@/��[�3@n�G:Ȑ!?�!2ڭ�@w���ٿ�׷�Ww�@#����3@꿗䜐!?����n�@w���ٿ�׷�Ww�@#����3@꿗䜐!?����n�@;����ٿ��y�t�@/#�{�3@#���!?d�W��@;����ٿ��y�t�@/#�{�3@#���!?d�W��@;����ٿ��y�t�@/#�{�3@#���!?d�W��@;����ٿ��y�t�@/#�{�3@#���!?d�W��@�$�E@�ٿUr�6���@�8�2�3@Hf��!?&!>x|S�@�$�E@�ٿUr�6���@�8�2�3@Hf��!?&!>x|S�@ZaޑA�ٿ#�zD�6�@�ʽ˕�3@i5�*��!?���#���@ZaޑA�ٿ#�zD�6�@�ʽ˕�3@i5�*��!?���#���@ZaޑA�ٿ#�zD�6�@�ʽ˕�3@i5�*��!?���#���@ZaޑA�ٿ#�zD�6�@�ʽ˕�3@i5�*��!?���#���@ZaޑA�ٿ#�zD�6�@�ʽ˕�3@i5�*��!?���#���@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@MON�,�ٿ>��S`��@8�3D��3@��h��!?Yr� 9�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@Irdަ�ٿ2*���B�@y�%���3@g�%D��!?L�j,�@�fl�ٿ�CIb��@������3@:��7Ȑ!?�9p�Y�@�fl�ٿ�CIb��@������3@:��7Ȑ!?�9p�Y�@}6��ٿ�u�'��@����}�3@^$���!?�C��'�@w�rM�ٿTRl�x�@�f��k�3@�p�+�!?p�����@ۓ�/��ٿ��5���@����P�3@�4ٖː!?#���n��@ۓ�/��ٿ��5���@����P�3@�4ٖː!?#���n��@�n[��ٿ�;���M�@>2�%��3@%�N�!?�����@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@��f���ٿ��
+x�@��x,�3@���z��!?�R�{\_�@�d���ٿ:l,V)�@�)g�3@<)ߥ��!?��_8z�@�d���ٿ:l,V)�@�)g�3@<)ߥ��!?��_8z�@�d���ٿ:l,V)�@�)g�3@<)ߥ��!?��_8z�@��V\g�ٿ�AcN��@VGW��3@z�MU��!?��	�ek�@��V\g�ٿ�AcN��@VGW��3@z�MU��!?��	�ek�@��V\g�ٿ�AcN��@VGW��3@z�MU��!?��	�ek�@��K�ٿ�E�'�I�@���(�3@�9�p�!?�0� ܩ�@��K�ٿ�E�'�I�@���(�3@�9�p�!?�0� ܩ�@��K�ٿ�E�'�I�@���(�3@�9�p�!?�0� ܩ�@B ��ٿ�j��,��@�!R`�3@��׬��!?�u�i1�@h;i�ٿU�6%׃�@��.	�3@��Z�ǐ!?��RO���@h;i�ٿU�6%׃�@��.	�3@��Z�ǐ!?��RO���@h;i�ٿU�6%׃�@��.	�3@��Z�ǐ!?��RO���@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@g���ٿm7fύ��@�+��3@4,�ڐ!?R�9ۃ��@�~�_�ٿ��=	��@�u6��3@!]�0��!?���wB�@�~�_�ٿ��=	��@�u6��3@!]�0��!?���wB�@����ٿ�Ɠ�#]�@u�1��3@[xi�!?����Aj�@����ٿ�Ɠ�#]�@u�1��3@[xi�!?����Aj�@�+����ٿ+j=�SG�@�����3@�*q���!?���h�l�@�+����ٿ+j=�SG�@�����3@�*q���!?���h�l�@����j�ٿɾc���@��/.��3@=�~T��!?=Q�yls�@����j�ٿɾc���@��/.��3@=�~T��!?=Q�yls�@����j�ٿɾc���@��/.��3@=�~T��!?=Q�yls�@����j�ٿɾc���@��/.��3@=�~T��!?=Q�yls�@����ٿu��&/�@�;�3@F\���!?W�q: R�@o"!"d�ٿ؇�q�a�@zd�~��3@��զ�!?�|�L4��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@�#q�ٿg  8|�@.Үgt�3@a�'pܐ!?M�[ ��@T}�{��ٿ�����G�@��G���3@��++�!?+/�_�I�@T}�{��ٿ�����G�@��G���3@��++�!?+/�_�I�@T}�{��ٿ�����G�@��G���3@��++�!?+/�_�I�@T}�{��ٿ�����G�@��G���3@��++�!?+/�_�I�@<T�U֜ٿ\�kB�@����3@z����!?�	���@<T�U֜ٿ\�kB�@����3@z����!?�	���@�%��'�ٿ/�8����@�b�]�3@T�KO�!?)�|����@�%��'�ٿ/�8����@�b�]�3@T�KO�!?)�|����@�%��'�ٿ/�8����@�b�]�3@T�KO�!?)�|����@�%��'�ٿ/�8����@�b�]�3@T�KO�!?)�|����@�%��'�ٿ/�8����@�b�]�3@T�KO�!?)�|����@�Z�x�ٿ:t��-+�@�$Fu��3@ݨ�
ِ!?�������@�Z�x�ٿ:t��-+�@�$Fu��3@ݨ�
ِ!?�������@�Z�x�ٿ:t��-+�@�$Fu��3@ݨ�
ِ!?�������@�Ai1�ٿKbP�}��@/~j�y�3@5b�9�!?�Қ�c:�@�Ai1�ٿKbP�}��@/~j�y�3@5b�9�!?�Қ�c:�@A��튠ٿ��d"Q��@s#�;�3@�)�!?��eb/�@Kt�6�ٿ�cv>�@��� ��3@�	��ِ!?a�Ȱ�r�@��XX��ٿ*Г�[�@E���F�3@e2���!?L��i��@��XX��ٿ*Г�[�@E���F�3@e2���!?L��i��@i��8�ٿ���?2��@���
��3@�0(z�!?dXg�T�@i��8�ٿ���?2��@���
��3@�0(z�!?dXg�T�@i��8�ٿ���?2��@���
��3@�0(z�!?dXg�T�@i��8�ٿ���?2��@���
��3@�0(z�!?dXg�T�@i��8�ٿ���?2��@���
��3@�0(z�!?dXg�T�@x�ӜٿG�nŦ��@n�,�!�3@od�
�!?N?��1n�@x�ӜٿG�nŦ��@n�,�!�3@od�
�!?N?��1n�@������ٿ� �����@��i��3@�s�!?E:��c��@������ٿ� �����@��i��3@�s�!?E:��c��@������ٿ� �����@��i��3@�s�!?E:��c��@E�u���ٿ��z�@7@�T�3@3Pw9�!?��	�#�@E�u���ٿ��z�@7@�T�3@3Pw9�!?��	�#�@E�u���ٿ��z�@7@�T�3@3Pw9�!?��	�#�@���.�ٿ��W�@�K�3@J�S��!?Z~3�(��@���.�ٿ��W�@�K�3@J�S��!?Z~3�(��@���.�ٿ��W�@�K�3@J�S��!?Z~3�(��@���.�ٿ��W�@�K�3@J�S��!?Z~3�(��@���.�ٿ��W�@�K�3@J�S��!?Z~3�(��@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@[��D��ٿ[�,�JD�@�^q�j�3@ۘ��!?���1�@X���p�ٿ�'�V?��@�	���3@ޔ�=ʐ!?$���TF�@X���p�ٿ�'�V?��@�	���3@ޔ�=ʐ!?$���TF�@X���p�ٿ�'�V?��@�	���3@ޔ�=ʐ!?$���TF�@%��A��ٿ���U%1�@�z��3@�����!?ꂻE
��@2 �6�ٿ:~N���@�9�{��3@��3��!?%���n��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�)�E�ٿ� 5	�@>n
���3@g�����!?{D��Q��@�/��ٿ�`U3���@O�<�{�3@�:-�!?i��A��@�/��ٿ�`U3���@O�<�{�3@�:-�!?i��A��@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@�i��ٿu[�x��@.2��$�3@���q�!?�A�����@��(�Ǡٿ�7\"U��@z��T��3@��A8!�!?���cf�@+\�^�ٿ�����@S�����3@߸� �!?�1�'�(�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@�F��;�ٿr��9��@�e��3@��u�א!?�l�|J5�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@��T�ٿ���P�@�_����3@��Ґ!?x�'Kb�@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@*���ܝٿ��켹q�@�m��3@�b��!?�P5 �@�傩e�ٿJ�_x$�@���s�3@�z� �!?�
��7�@%�PC�ٿ���zfO�@}���3@7�����!?�����R�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@CW�}�ٿ�Iu�Z�@_،H�3@_��E��!?GF-ƍ*�@/�B��ٿ-����U�@�Bڷ��3@��Z���!?�֛��m�@/�B��ٿ-����U�@�Bڷ��3@��Z���!?�֛��m�@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@�DE��ٿ'������@�8=�"�3@�q͹k�!?)�?&���@��E�ʛٿ����;�@}44@�3@1�M*�!?p��-��@��E�ʛٿ����;�@}44@�3@1�M*�!?p��-��@��E�ʛٿ����;�@}44@�3@1�M*�!?p��-��@��E�ʛٿ����;�@}44@�3@1�M*�!?p��-��@1CINڞٿ)mV@��@�Xb�j�3@�Zy\'�!?NA�݁�@1CINڞٿ)mV@��@�Xb�j�3@�Zy\'�!?NA�݁�@1CINڞٿ)mV@��@�Xb�j�3@�Zy\'�!?NA�݁�@1CINڞٿ)mV@��@�Xb�j�3@�Zy\'�!?NA�݁�@7֡���ٿ"]�¾��@�~R�Y�3@f����!?���9	g�@7֡���ٿ"]�¾��@�~R�Y�3@f����!?���9	g�@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@>{��ٿ������@�-#��3@�⧏�!?���S��@�GVI͢ٿ{�S�� �@��Z��3@V"ʁ��!?�+���@�GVI͢ٿ{�S�� �@��Z��3@V"ʁ��!?�+���@�GVI͢ٿ{�S�� �@��Z��3@V"ʁ��!?�+���@�GVI͢ٿ{�S�� �@��Z��3@V"ʁ��!?�+���@�Ĵ&�ٿ�#��@p���3@�\�!?� T���@N�_�P�ٿ���!�@��7m��3@h�vΐ!?А���D�@N�_�P�ٿ���!�@��7m��3@h�vΐ!?А���D�@N�_�P�ٿ���!�@��7m��3@h�vΐ!?А���D�@�mF�r�ٿ�gB���@p����3@3��!?�/�,ic�@�mF�r�ٿ�gB���@p����3@3��!?�/�,ic�@����ٿ�!�#��@�G<#5�3@7�e��!?�%�T>j�@����ٿ�!�#��@�G<#5�3@7�e��!?�%�T>j�@%`4|��ٿ*��D^��@�� VM�3@"!��<�!?��$Pr�@��Pۛٿ{̗Y@��@�
��\�3@��@C�!?�֒��@��Pۛٿ{̗Y@��@�
��\�3@��@C�!?�֒��@��Pۛٿ{̗Y@��@�
��\�3@��@C�!?�֒��@��Pۛٿ{̗Y@��@�
��\�3@��@C�!?�֒��@
� �ٿ��Y�m�@�,pMQ�3@��w�!?O�K7���@
� �ٿ��Y�m�@�,pMQ�3@��w�!?O�K7���@�r),�ٿ�����@!�cg* 4@n��J�!?a��9o��@T͊�A�ٿ��-��@�û�C�3@����!?t�1@�@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@�p�ğ�ٿ.I����@S��˹�3@rdM�!?�� ��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@m��w�ٿ����uc�@���3��3@d�n֐!?_~֛X��@�ɏ8z�ٿ׉����@F8<}�3@��(�c�!?��:H�@�ɏ8z�ٿ׉����@F8<}�3@��(�c�!?��:H�@�ɏ8z�ٿ׉����@F8<}�3@��(�c�!?��:H�@�ɏ8z�ٿ׉����@F8<}�3@��(�c�!?��:H�@�1�P�ٿ,����@k��7��3@�+%�w�!?>�⨈v�@�1�P�ٿ,����@k��7��3@�+%�w�!?>�⨈v�@�1�P�ٿ,����@k��7��3@�+%�w�!?>�⨈v�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@>5���ٿ�]��[�@�����3@2�����!?���<2%�@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@?��ٿ)&��z�@���t�3@���q��!?,i��N��@w�)��ٿa~r�'�@�=����3@��fHK�!?>DF}m��@w�)��ٿa~r�'�@�=����3@��fHK�!?>DF}m��@w�)��ٿa~r�'�@�=����3@��fHK�!?>DF}m��@w�)��ٿa~r�'�@�=����3@��fHK�!?>DF}m��@~6��͞ٿen�m;�@���T�3@E�;��!?1��~�@~6��͞ٿen�m;�@���T�3@E�;��!?1��~�@~6��͞ٿen�m;�@���T�3@E�;��!?1��~�@}׍$ٿ�OM@i�@�R,�}�3@Ja~�!?IT����@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@¸Ez�ٿt`��@�kP��3@�!���!?�4"ob��@U��j��ٿ��s��@᯲"��3@�%��!?C�&��@U��j��ٿ��s��@᯲"��3@�%��!?C�&��@U��j��ٿ��s��@᯲"��3@�%��!?C�&��@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@�cd��ٿ�.P�"��@P�K��3@eEQ4��!?C9eR�@57��ݝٿ�Ֆ>�@���\��3@	˭�!?
78-��@Q�Y���ٿ� }�?�@A�q�3@��!�!?�qgv;2�@�h����ٿ�~XwF�@�>���3@���8�!??mU�!��@�h����ٿ�~XwF�@�>���3@���8�!??mU�!��@�h����ٿ�~XwF�@�>���3@���8�!??mU�!��@�h����ٿ�~XwF�@�>���3@���8�!??mU�!��@�����ٿ����t�@[xl�	�3@�3�C��!?o�`�j��@�����ٿ����t�@[xl�	�3@�3�C��!?o�`�j��@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�	��'�ٿ�@���@"�P�3@�jr�͐!?�I�	�h�@�Y�<h�ٿ�9+:��@V����3@$	c1o�!?�:�ޛ�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@4� 6�ٿ�e]j��@�O��3@"ja�!?m�|�w�@	����ٿW�����@`QG+�3@E.`iy�!?���A���@�h]�ٿ��H	�@:\�d�3@W����!?/x��@�h]�ٿ��H	�@:\�d�3@W����!?/x��@�h]�ٿ��H	�@:\�d�3@W����!?/x��@�h]�ٿ��H	�@:\�d�3@W����!?/x��@�h]�ٿ��H	�@:\�d�3@W����!?/x��@�h]�ٿ��H	�@:\�d�3@W����!?/x��@5���ٿ�p�{���@k�',�3@� \(�!?5�A{���@5���ٿ�p�{���@k�',�3@� \(�!?5�A{���@5���ٿ�p�{���@k�',�3@� \(�!?5�A{���@5���ٿ�p�{���@k�',�3@� \(�!?5�A{���@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@�8	��ٿ�g�3�9�@���.��3@τǌW�!?�!L��'�@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@\*\s�ٿd0?̸��@5�Ղ7�3@N��|�!?�Z����@A�6��ٿS�?�FC�@�x\��3@^6���!?�q/G��@�Q����ٿ�O�Y�{�@uF)�3@��F��!?�X�&��@�Q����ٿ�O�Y�{�@uF)�3@��F��!?�X�&��@�Q����ٿ�O�Y�{�@uF)�3@��F��!?�X�&��@�Q����ٿ�O�Y�{�@uF)�3@��F��!?�X�&��@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@��ܛٿ(���@��FXV�3@��8���!?{�g&ц�@#۴��ٿ�^��-�@�ܖ��3@�,r���!?:�J!�@#۴��ٿ�^��-�@�ܖ��3@�,r���!?:�J!�@#۴��ٿ�^��-�@�ܖ��3@�,r���!?:�J!�@#۴��ٿ�^��-�@�ܖ��3@�,r���!?:�J!�@#۴��ٿ�^��-�@�ܖ��3@�,r���!?:�J!�@�lʱ�ٿ_4�u�@ҧH�3@Hb����!?5�Zn$��@�lʱ�ٿ_4�u�@ҧH�3@Hb����!?5�Zn$��@�lʱ�ٿ_4�u�@ҧH�3@Hb����!?5�Zn$��@�lʱ�ٿ_4�u�@ҧH�3@Hb����!?5�Zn$��@�lʱ�ٿ_4�u�@ҧH�3@Hb����!?5�Zn$��@�� �<�ٿ��H����@� %y�3@�Ύɽ�!?���0��@�� �<�ٿ��H����@� %y�3@�Ύɽ�!?���0��@�%|ꁛٿ��K�M��@C:�ZY�3@}WBBؐ!?�k�Ο�@�%|ꁛٿ��K�M��@C:�ZY�3@}WBBؐ!?�k�Ο�@�%|ꁛٿ��K�M��@C:�ZY�3@}WBBؐ!?�k�Ο�@�%|ꁛٿ��K�M��@C:�ZY�3@}WBBؐ!?�k�Ο�@ᕌ�"�ٿ�~ ��$�@�Q瑋�3@��!?��qJ�@g����ٿ:C� 1H�@F�L�3@_^|x�!?�2aʽU�@�l��U�ٿ/�A�e�@2~��3@Mx���!?Bh�B�@�l��U�ٿ/�A�e�@2~��3@Mx���!?Bh�B�@�M��+�ٿ4C��K�@�L��X�3@�m�[ݐ!?E�`sLf�@�Q���ٿ"������@Z����3@j1�!?�{���@�Q���ٿ"������@Z����3@j1�!?�{���@�Q���ٿ"������@Z����3@j1�!?�{���@�Q���ٿ"������@Z����3@j1�!?�{���@�Q���ٿ"������@Z����3@j1�!?�{���@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@�qB@~�ٿ�<�b�@vӟv%�3@���~Ő!?�z��m�@#^��j�ٿ��zY��@����3@����!?DL���I�@#^��j�ٿ��zY��@����3@����!?DL���I�@#^��j�ٿ��zY��@����3@����!?DL���I�@��\>�ٿ�q�x��@�D���3@P̐!?�6^/�H�@�;�ٿ�ַ�x��@�����3@�>�Đ!?`kdm�@�;�ٿ�ַ�x��@�����3@�>�Đ!?`kdm�@�;�ٿ�ַ�x��@�����3@�>�Đ!?`kdm�@�"�RQ�ٿ�.�9�3�@.����3@��=��!?X�磧�@�"�RQ�ٿ�.�9�3�@.����3@��=��!?X�磧�@�"�RQ�ٿ�.�9�3�@.����3@��=��!?X�磧�@.����ٿ�.CA���@�4tq�3@�V��!?�����@.����ٿ�.CA���@�4tq�3@�V��!?�����@.����ٿ�.CA���@�4tq�3@�V��!?�����@.����ٿ�.CA���@�4tq�3@�V��!?�����@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@G�X�X�ٿ�& �q�@2����3@	����!?-�v���@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@�[���ٿ=�eZ��@W@HGF�3@&}-��!?�f��@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@� Ή�ٿ�w�k��@�]>@��3@�;���!?�Uа�@դDC٢ٿwp>��l�@��q��3@�]����!?��?F��@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��d���ٿO���/�@'��*E�3@��}�z�!?9ίf:�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@��j:�ٿ���֌�@i�^�d�3@�Y�]{�!?p�U�r3�@J�1m�ٿ<)�u1�@&�j4�3@��b�Y�!?�T��@J�1m�ٿ<)�u1�@&�j4�3@��b�Y�!?�T��@r���3�ٿ�8 ���@� �9D�3@���K}�!?���f���@�Тٿ@Rs(�@�w�|�3@F��1��!?�?Ö��@�Тٿ@Rs(�@�w�|�3@F��1��!?�?Ö��@Q><��ٿ��M����@���I{�3@%@�µ�!?���e�@Q><��ٿ��M����@���I{�3@%@�µ�!?���e�@Q><��ٿ��M����@���I{�3@%@�µ�!?���e�@(��%��ٿ\]ITM��@�C*�3@]
����!?9%�5v�@(��%��ٿ\]ITM��@�C*�3@]
����!?9%�5v�@(��%��ٿ\]ITM��@�C*�3@]
����!?9%�5v�@(��%��ٿ\]ITM��@�C*�3@]
����!?9%�5v�@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@+O�#ިٿ��د�@��d��3@�C4�z�!?���B��@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@��D�ٿX�J�@6��|��3@�jI��!?�,D߼+�@�9����ٿ��@����@�2� 4@nTo<��!?�B>�l:�@�9����ٿ��@����@�2� 4@nTo<��!?�B>�l:�@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@l�K��ٿ��r��@��q��3@H?1M�!?�A^WV��@:�F��ٿbᥲF�@���9X�3@�;ʐ!?A�q�BM�@:�F��ٿbᥲF�@���9X�3@�;ʐ!?A�q�BM�@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@�+�/�ٿƂ�%���@�c����3@jh�b��!?R�����@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@@�ߣ��ٿϱ,�%��@V!��~�3@�1�h��!?��� u��@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@���;�ٿ��0¨��@H��f��3@��;���!?Fb�dV�@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@W�ԛC�ٿw"Ni���@�O���3@�)���!?�6�w��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@����ٿ�/�/��@=v�,��3@̘A�$�!?4O��+��@t�-���ٿ`�����@kb�f�3@��B'�!?'����@�:���ٿ���ܮ��@3�;M��3@Iܵ���!?�����@��HKv�ٿ�s�\�@�Z1b��3@�&h�А!?*M*L��@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@l��Mj�ٿ_N_���@Q3�"��3@O��mb�!?g� _�@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@��WWêٿ�8\��@Z�	��3@f��y�!?�A���@�dv T�ٿ'5���@$^����3@U/����!?�1�Y1�@�6|��ٿ3kU�@:D���3@�ub���!?�
j�P�@�o�[�ٿef#�@�a��3@�dѓ��!?�������@�o�[�ٿef#�@�a��3@�dѓ��!?�������@gv�OT�ٿ�B]U*�@f��N��3@^�
EĐ!?pm�>���@gv�OT�ٿ�B]U*�@f��N��3@^�
EĐ!?pm�>���@gv�OT�ٿ�B]U*�@f��N��3@^�
EĐ!?pm�>���@gv�OT�ٿ�B]U*�@f��N��3@^�
EĐ!?pm�>���@��:��ٿz�`kR�@�"2�V�3@c��ѐ!?�D}�n2�@ک��ٿ��,0���@3�0���3@l ?��!?$�	<�@ک��ٿ��,0���@3�0���3@l ?��!?$�	<�@ک��ٿ��,0���@3�0���3@l ?��!?$�	<�@ک��ٿ��,0���@3�0���3@l ?��!?$�	<�@�Ѣ��ٿr��1�@���3@����\�!?�hxPYR�@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@*?�ٿt������@�f��3@:�w��!?�,&l��@�+Ƥٿ�dKO4-�@y�����3@2�ʐ!?vCG�|>�@�+Ƥٿ�dKO4-�@y�����3@2�ʐ!?vCG�|>�@�+Ƥٿ�dKO4-�@y�����3@2�ʐ!?vCG�|>�@�+Ƥٿ�dKO4-�@y�����3@2�ʐ!?vCG�|>�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�J��͝ٿ����9�@�G��3@z�|�!?&LE�J�@�C�8~�ٿh\ި���@���o��3@���Đ!?42���e�@�C�8~�ٿh\ި���@���o��3@���Đ!?42���e�@f��	�ٿ7o�?�@�����3@����!?n�7�3z�@f��	�ٿ7o�?�@�����3@����!?n�7�3z�@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@�M�ٿ�8��68�@5e��x�3@�-���!?A�j7��@��)�ٿ� k
R�@�����3@�#v���!?xʛB)�@{�f5�ٿ����~�@�B�2��3@uߨ���!?n�K�ZB�@{�f5�ٿ����~�@�B�2��3@uߨ���!?n�K�ZB�@{�f5�ٿ����~�@�B�2��3@uߨ���!?n�K�ZB�@��Z
Пٿa�E:��@WW����3@��wSȐ!?��A���@��Z
Пٿa�E:��@WW����3@��wSȐ!?��A���@��Z
Пٿa�E:��@WW����3@��wSȐ!?��A���@��Z
Пٿa�E:��@WW����3@��wSȐ!?��A���@%�h���ٿ���}�@�(�F>�3@��{��!?d�e����@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@Lp�ۘ�ٿp�_���@rⵍ�3@e'�.t�!?����F�@�@�'�ٿ�f���$�@,���3@x#d�y�!?�Z[��@t;y}��ٿ�+�]�@��4��3@W/�!?���R��@t;y}��ٿ�+�]�@��4��3@W/�!?���R��@t;y}��ٿ�+�]�@��4��3@W/�!?���R��@抖��ٿ��? ���@j�&���3@sv�oz�!?�:@.a;�@抖��ٿ��? ���@j�&���3@sv�oz�!?�:@.a;�@抖��ٿ��? ���@j�&���3@sv�oz�!?�:@.a;�@抖��ٿ��? ���@j�&���3@sv�oz�!?�:@.a;�@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@䡸���ٿE"f��@ �����3@#�4a�!?]ފy��@�ו)�ٿP�N���@�(��h�3@r幚��!?�C)��G�@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@�	NE��ٿ�}^����@n�ȁ��3@���s��!?�aq����@b�H���ٿ���{N��@��B���3@�]�a��!?^���V��@b�H���ٿ���{N��@��B���3@�]�a��!?^���V��@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@����&�ٿp�Qt��@��c0��3@�
���!?~k��+�@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@8S���ٿշN5��@D�2��3@�mօ�!?��PA��@PE�!J�ٿ���:��@�J�� �3@��&���!?�c�۰a�@PE�!J�ٿ���:��@�J�� �3@��&���!?�c�۰a�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@|@�N�ٿ	�����@Qn����3@q��ʝ�!?�U�z�G�@�1	�ʝٿЄgDB�@�ir�3@��qd�!?�����@�1	�ʝٿЄgDB�@�ir�3@��qd�!?�����@��.��ٿ����/�@z� ���3@p�8I��!?yq)�E��@��.��ٿ����/�@z� ���3@p�8I��!?yq)�E��@��.��ٿ����/�@z� ���3@p�8I��!?yq)�E��@��R��ٿЅ�J�@!@���3@�s��f�!?4�4(���@��R��ٿЅ�J�@!@���3@�s��f�!?4�4(���@	�L�ٿӒ�u �@�v�?�3@Ғ=u��!?��ɑ��@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@����T�ٿ0�U��@��d4@�3@ټ;�s�!?�L�/�Q�@Y� ؤٿ��jy��@��j`�3@�%��!?�l�����@Y� ؤٿ��jy��@��j`�3@�%��!?�l�����@Y� ؤٿ��jy��@��j`�3@�%��!?�l�����@Y� ؤٿ��jy��@��j`�3@�%��!?�l�����@eХ��ٿ��x[&�@Ry����3@�iм�!?�����@eХ��ٿ��x[&�@Ry����3@�iм�!?�����@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@�Mh�ٿwF栤�@���e�3@�vbdِ!?<�?b ��@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@֝o�Ρٿ�!����@�EG@+�3@���ː!?�z���@R�4p$�ٿ�]m�F��@�����3@��
+��!?�V�,��@R�4p$�ٿ�]m�F��@�����3@��
+��!?�V�,��@R�4p$�ٿ�]m�F��@�����3@��
+��!?�V�,��@R�4p$�ٿ�]m�F��@�����3@��
+��!?�V�,��@m��{�ٿj򢆀�@ͫ��n�3@E��lx�!?��'��@m��{�ٿj򢆀�@ͫ��n�3@E��lx�!?��'��@m��{�ٿj򢆀�@ͫ��n�3@E��lx�!?��'��@m��{�ٿj򢆀�@ͫ��n�3@E��lx�!?��'��@m��{�ٿj򢆀�@ͫ��n�3@E��lx�!?��'��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@���8��ٿ�%���@��!���3@%]�z�!?��U@��@� ;LΛٿ��~Q�@D����3@i�g���!?�a1rc��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@^��ٿP�A��Y�@D�[>R�3@c�/�s�!?��q�:��@��ߩ��ٿ'/*=6��@,�"��3@vc�n�!?�μ�Ҿ�@��ߩ��ٿ'/*=6��@,�"��3@vc�n�!?�μ�Ҿ�@��ߩ��ٿ'/*=6��@,�"��3@vc�n�!?�μ�Ҿ�@��ߩ��ٿ'/*=6��@,�"��3@vc�n�!?�μ�Ҿ�@��ߩ��ٿ'/*=6��@,�"��3@vc�n�!?�μ�Ҿ�@}��s��ٿ���t��@��j�t�3@��,蛐!?X]�{��@}��s��ٿ���t��@��j�t�3@��,蛐!?X]�{��@}��s��ٿ���t��@��j�t�3@��,蛐!?X]�{��@�����ٿU�O�/�@[�'u��3@6�����!?a�XX���@	��� �ٿf�;�X�@]p�3@J�MȐ!?�'M����@	��� �ٿf�;�X�@]p�3@J�MȐ!?�'M����@	��� �ٿf�;�X�@]p�3@J�MȐ!?�'M����@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@���-�ٿ4��%^;�@(S�S�3@'{O���!?��oQ�,�@�?.�ٿ�V�@���l��3@����ǐ!?3̳cS�@�?.�ٿ�V�@���l��3@����ǐ!?3̳cS�@����ٿG����'�@F2E]��3@h5�֒�!?��l��@����ٿG����'�@F2E]��3@h5�֒�!?��l��@����ٿG����'�@F2E]��3@h5�֒�!?��l��@����ٿG����'�@F2E]��3@h5�֒�!?��l��@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@����ٿG~[��@5����3@��@{�!?C��S���@�C�d�ٿ �η�@�"����3@"\	6А!?Z�0�@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�C?g]�ٿ0�����@'Z/��3@�)}�ʐ!?�~e��@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@�}��ٿ�OYI�@��8�^�3@�0T�ѐ!?��z݋�@g��k�ٿ�9_���@ڜ�Á�3@����!?��ay�@g��k�ٿ�9_���@ڜ�Á�3@����!?��ay�@g��k�ٿ�9_���@ڜ�Á�3@����!?��ay�@�g˥��ٿ��Wi�@M�d�3@���k��!?o�z\���@�g˥��ٿ��Wi�@M�d�3@���k��!?o�z\���@�g˥��ٿ��Wi�@M�d�3@���k��!?o�z\���@۠���ٿ͟P6O��@Sgiv�3@��lW��!?�EA����@۠���ٿ͟P6O��@Sgiv�3@��lW��!?�EA����@۠���ٿ͟P6O��@Sgiv�3@��lW��!?�EA����@۠���ٿ͟P6O��@Sgiv�3@��lW��!?�EA����@�D�=��ٿц�����@S���3@�UO�q�!?E���	��@�D�=��ٿц�����@S���3@�UO�q�!?E���	��@������ٿc�"c]�@ܮ�4�3@ ��ɐ!?�y�O�@������ٿc�"c]�@ܮ�4�3@ ��ɐ!?�y�O�@������ٿc�"c]�@ܮ�4�3@ ��ɐ!?�y�O�@������ٿc�"c]�@ܮ�4�3@ ��ɐ!?�y�O�@�K?�ٿ���:��@q�Z*s�3@�g��o�!?ǀ��E�@�K?�ٿ���:��@q�Z*s�3@�g��o�!?ǀ��E�@�K?�ٿ���:��@q�Z*s�3@�g��o�!?ǀ��E�@pb�U�ٿ��/�k��@�ը��3@�>��f�!?Y;.B�-�@C��ٿ6�>
Z�@#�]���3@d$���!? $h�@m���R�ٿ���>�@x��U�3@�0��b�!?�� F���@m���R�ٿ���>�@x��U�3@�0��b�!?�� F���@m���R�ٿ���>�@x��U�3@�0��b�!?�� F���@m���R�ٿ���>�@x��U�3@�0��b�!?�� F���@m���R�ٿ���>�@x��U�3@�0��b�!?�� F���@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@om��ٿ�Ch��@� �ػ�3@��+��!?�2T��@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@~^�eנٿ�
���@x#���3@MWX�ʐ!?r_=����@ؼp\�ٿ$�nOrT�@uD__\�3@$k�!?=C�G��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@����ٿ:�����@/�Mw�3@����{�!?�՞D��@�?���ٿR�p�RP�@.^A���3@����!?�؅����@l"Q���ٿ3i�Nh�@�ns?�3@�����!?~���4�@/����ٿ���fJ��@:͹��3@Av��ǐ!?�L0�L�@/����ٿ���fJ��@:͹��3@Av��ǐ!?�L0�L�@/����ٿ���fJ��@:͹��3@Av��ǐ!?�L0�L�@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@
U�=��ٿ�7�W��@{�e���3@�pض�!?�����@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@���s��ٿ;(uM|�@��6�3@T�Ɛ!?Ad-��@#�;hK�ٿH�KD�@z����3@�\$��!?-4"C��@#�;hK�ٿH�KD�@z����3@�\$��!?-4"C��@#�;hK�ٿH�KD�@z����3@�\$��!?-4"C��@���]�ٿI�p��@�%����3@���J~�!?CQ��8�@���p�ٿ���]��@�'o4 �3@���蟐!?���ٗ��@���p�ٿ���]��@�'o4 �3@���蟐!?���ٗ��@E<��i�ٿ�6�� ��@^���2�3@�ďܐ!?�2U��@E<��i�ٿ�6�� ��@^���2�3@�ďܐ!?�2U��@��j�Þٿ�\�h��@λ���3@��@�!?����W�@��j�Þٿ�\�h��@λ���3@��@�!?����W�@��j�Þٿ�\�h��@λ���3@��@�!?����W�@��j�Þٿ�\�h��@λ���3@��@�!?����W�@J���M�ٿ9�C���@M0	���3@�oص8�!?C�H���@J���M�ٿ9�C���@M0	���3@�oص8�!?C�H���@�C4�ٿH�4�>�@��a-��3@R�%=�!?�����@�C4�ٿH�4�>�@��a-��3@R�%=�!?�����@�C4�ٿH�4�>�@��a-��3@R�%=�!?�����@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@�e��՛ٿ�Z��$�@D��F�3@�v�O��!?�K,5h��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@yV.۸�ٿ��"W��@F��_��3@�}縐!?<��
��@q�a���ٿ)�0P��@���!�3@��p멐!?:g��X��@��	��ٿ	3����@my�|9�3@b�m���!?�ۀ�b,�@��	��ٿ	3����@my�|9�3@b�m���!?�ۀ�b,�@��	��ٿ	3����@my�|9�3@b�m���!?�ۀ�b,�@��	��ٿ	3����@my�|9�3@b�m���!?�ۀ�b,�@��	��ٿ	3����@my�|9�3@b�m���!?�ۀ�b,�@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@<ai��ٿ7�"����@���x�3@��/'��!?O�'.��@+�ɟ�ٿ�
�^���@>z?n�3@@M��!?�	�-�@+�ɟ�ٿ�
�^���@>z?n�3@@M��!?�	�-�@+�ɟ�ٿ�
�^���@>z?n�3@@M��!?�	�-�@+�ɟ�ٿ�
�^���@>z?n�3@@M��!?�	�-�@+�ɟ�ٿ�
�^���@>z?n�3@@M��!?�	�-�@�+��ٿ9�>LHp�@
�q�3@���܏�!?��8?�k�@�+��ٿ9�>LHp�@
�q�3@���܏�!?��8?�k�@�+��ٿ9�>LHp�@
�q�3@���܏�!?��8?�k�@�(�`�ٿ|]u��@�PC���3@v�-�!?��gN	��@�(�`�ٿ|]u��@�PC���3@v�-�!?��gN	��@�(�`�ٿ|]u��@�PC���3@v�-�!?��gN	��@�(�`�ٿ|]u��@�PC���3@v�-�!?��gN	��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@E�˝ٿ��S΄�@xS-a�3@p��ː!?9�~7d��@��-h�ٿ�t/a�}�@XFaX��3@�:ߐ��!?9aN�@��-h�ٿ�t/a�}�@XFaX��3@�:ߐ��!?9aN�@��-h�ٿ�t/a�}�@XFaX��3@�:ߐ��!?9aN�@b�����ٿ����@;�����3@���]ΐ!?k���ۿ�@b�����ٿ����@;�����3@���]ΐ!?k���ۿ�@b�����ٿ����@;�����3@���]ΐ!?k���ۿ�@b�����ٿ����@;�����3@���]ΐ!?k���ۿ�@p��xǟٿD�筷�@e�"p�3@9��Y �!?��4�@p��xǟٿD�筷�@e�"p�3@9��Y �!?��4�@˟Ȯ��ٿ��kpƀ�@4�)�`�3@��N�+�!?"�f�!�@˟Ȯ��ٿ��kpƀ�@4�)�`�3@��N�+�!?"�f�!�@b;<7ۣٿ��D�1\�@��(��3@�6�!?}Ҍ�f�@b;<7ۣٿ��D�1\�@��(��3@�6�!?}Ҍ�f�@b;<7ۣٿ��D�1\�@��(��3@�6�!?}Ҍ�f�@��6s�ٿKR���@��F_/4@�f���!?��Qw�@'�f��ٿU�!��x�@�Pj�4@�8Z���!?J�ܛ�@'�f��ٿU�!��x�@�Pj�4@�8Z���!?J�ܛ�@Z~��ٿ�`��k�@%�� ��3@��(�ې!?��6����@Z~��ٿ�`��k�@%�� ��3@��(�ې!?��6����@Z~��ٿ�`��k�@%�� ��3@��(�ې!?��6����@Z~��ٿ�`��k�@%�� ��3@��(�ې!?��6����@Z~��ٿ�`��k�@%�� ��3@��(�ې!?��6����@|���ٿP���f��@����3@^�}�x�!?�	C,�@|���ٿP���f��@����3@^�}�x�!?�	C,�@|���ٿP���f��@����3@^�}�x�!?�	C,�@|���ٿP���f��@����3@^�}�x�!?�	C,�@��zٔ�ٿ��WI"�@�WI�,�3@Ġ���!?�]�
��@��zٔ�ٿ��WI"�@�WI�,�3@Ġ���!?�]�
��@�vZ�ݟٿ�� ��@=|���3@ji��!?��Ql�@bO/���ٿW`8�S;�@��`���3@=�4�Ȑ!?��8e�r�@bO/���ٿW`8�S;�@��`���3@=�4�Ȑ!?��8e�r�@ւ�c�ٿ,��e�@��&V�3@�N�Ym�!?K�7tou�@Z)j��ٿp���|��@�^X��3@f!�_�!?��k��@Z)j��ٿp���|��@�^X��3@f!�_�!?��k��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@6��K۟ٿҾH\?��@�oܸ�3@�M&��!?�۟\&��@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@tP��_�ٿ����0�@�n#�3@L�#�z�!?��c����@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@К�i�ٿr���7$�@�Ope��3@Ձ�X�!?�F�'-��@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@N�
D��ٿ2�DpZ�@���.�3@�Ar�!?C�m��4�@*�}���ٿ$�����@Үq��3@D�h�v�!?�x�&1�@*�}���ٿ$�����@Үq��3@D�h�v�!?�x�&1�@*�}���ٿ$�����@Үq��3@D�h�v�!?�x�&1�@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@73�ƣ�ٿ�+�)�w�@�M,��3@�����!?=Jsa>��@o{�Ϥٿ�|��7[�@!8 9��3@:��o��!?�k��vW�@o{�Ϥٿ�|��7[�@!8 9��3@:��o��!?�k��vW�@o{�Ϥٿ�|��7[�@!8 9��3@:��o��!?�k��vW�@�xwj�ٿ����|%�@�!�	��3@��:��!?�����@�xwj�ٿ����|%�@�!�	��3@��:��!?�����@�xwj�ٿ����|%�@�!�	��3@��:��!?�����@�xwj�ٿ����|%�@�!�	��3@��:��!?�����@�xwj�ٿ����|%�@�!�	��3@��:��!?�����@T���ٿ�d?(�@��uB��3@Rǘ�!?i�~����@T���ٿ�d?(�@��uB��3@Rǘ�!?i�~����@T���ٿ�d?(�@��uB��3@Rǘ�!?i�~����@ڿ�8מٿheݶ[��@}�Y��3@�\�'�!?UA#7f�@ڿ�8מٿheݶ[��@}�Y��3@�\�'�!?UA#7f�@}u'��ٿ�1���@,lÀ��3@�9�vԐ!?kt��O��@}u'��ٿ�1���@,lÀ��3@�9�vԐ!?kt��O��@}u'��ٿ�1���@,lÀ��3@�9�vԐ!?kt��O��@}u'��ٿ�1���@,lÀ��3@�9�vԐ!?kt��O��@%o�Ҡ�ٿ~����@�~#�e�3@��7]Đ!?ø<=�k�@%o�Ҡ�ٿ~����@�~#�e�3@��7]Đ!?ø<=�k�@%o�Ҡ�ٿ~����@�~#�e�3@��7]Đ!?ø<=�k�@%o�Ҡ�ٿ~����@�~#�e�3@��7]Đ!?ø<=�k�@%o�Ҡ�ٿ~����@�~#�e�3@��7]Đ!?ø<=�k�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@�.-#ٿȌ�fS��@a�B��3@jK�!?�K̪zk�@+v�|w�ٿ�#>_��@Q٫�W�3@��wĺ�!?��gw�@+v�|w�ٿ�#>_��@Q٫�W�3@��wĺ�!?��gw�@+v�|w�ٿ�#>_��@Q٫�W�3@��wĺ�!?��gw�@+v�|w�ٿ�#>_��@Q٫�W�3@��wĺ�!?��gw�@+v�|w�ٿ�#>_��@Q٫�W�3@��wĺ�!?��gw�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@�XqP�ٿT{����@e�ac�3@dĽPt�!?���u$�@_k���ٿv���@��C��3@{Y��ΐ!?^��4��@K ���ٿC�����@����3@�o����!?E�6+�@����8�ٿ˹�&o�@�h;���3@��+;��!?zo�ߤ��@����8�ٿ˹�&o�@�h;���3@��+;��!?zo�ߤ��@��I�ٿ�W<_]��@�����3@K]�k�!?V��g���@'�|y �ٿI�Rʫ��@GJ��3@pv�p�!?�1`�n�@'�|y �ٿI�Rʫ��@GJ��3@pv�p�!?�1`�n�@'�|y �ٿI�Rʫ��@GJ��3@pv�p�!?�1`�n�@�F�[�ٿ�69�@���y�3@7U+!��!?�'7
��@�F�[�ٿ�69�@���y�3@7U+!��!?�'7
��@�F�[�ٿ�69�@���y�3@7U+!��!?�'7
��@�F�[�ٿ�69�@���y�3@7U+!��!?�'7
��@���7�ٿ���g���@e�2.�3@�����!?z��Pd�@���7�ٿ���g���@e�2.�3@�����!?z��Pd�@���7�ٿ���g���@e�2.�3@�����!?z��Pd�@���7�ٿ���g���@e�2.�3@�����!?z��Pd�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@� K�ٿڑ�����@f�)���3@�\)ސ!?N�v؂�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@�ѓ_�ٿ7� U�@�f��D�3@o�j/��!?Su�iV�@��c`�ٿ^At ~��@4?���3@��^2��!?^��*%W�@��c`�ٿ^At ~��@4?���3@��^2��!?^��*%W�@��c`�ٿ^At ~��@4?���3@��^2��!?^��*%W�@��c`�ٿ^At ~��@4?���3@��^2��!?^��*%W�@�6h�y�ٿ���!{��@P,#W�3@�~�Ȑ!?����9�@'�ٿ^P�9&:�@l%9��3@YT`G�!?��K��t�@'�ٿ^P�9&:�@l%9��3@YT`G�!?��K��t�@��
˥ٿ�����@�t�~�3@�vp��!?u�<���@��
˥ٿ�����@�t�~�3@�vp��!?u�<���@��
˥ٿ�����@�t�~�3@�vp��!?u�<���@��
˥ٿ�����@�t�~�3@�vp��!?u�<���@<Ea�ٿʉ]�ZO�@S2c�5�3@����Ӑ!?�(�)�2�@)�bL@�ٿ�����@h%�p�3@��^+t�!?��h1���@)�bL@�ٿ�����@h%�p�3@��^+t�!?��h1���@)�bL@�ٿ�����@h%�p�3@��^+t�!?��h1���@)�bL@�ٿ�����@h%�p�3@��^+t�!?��h1���@)�bL@�ٿ�����@h%�p�3@��^+t�!?��h1���@G�uB�ٿޔ����@x��h�3@����Đ!?VkQ��"�@G�uB�ٿޔ����@x��h�3@����Đ!?VkQ��"�@G�uB�ٿޔ����@x��h�3@����Đ!?VkQ��"�@G�uB�ٿޔ����@x��h�3@����Đ!?VkQ��"�@G�uB�ٿޔ����@x��h�3@����Đ!?VkQ��"�@�6$u�ٿi5\q4,�@q��dU�3@�u$ϐ�!?P��R"K�@�6$u�ٿi5\q4,�@q��dU�3@�u$ϐ�!?P��R"K�@�6$u�ٿi5\q4,�@q��dU�3@�u$ϐ�!?P��R"K�@�6$u�ٿi5\q4,�@q��dU�3@�u$ϐ�!?P��R"K�@%����ٿ�PA��$�@ɴ�҈�3@j
;Đ!?|���@%����ٿ�PA��$�@ɴ�҈�3@j
;Đ!?|���@%����ٿ�PA��$�@ɴ�҈�3@j
;Đ!?|���@��-}�ٿ$JS��"�@0��}�3@�G6�ʐ!?����G��@��-}�ٿ$JS��"�@0��}�3@�G6�ʐ!?����G��@��-}�ٿ$JS��"�@0��}�3@�G6�ʐ!?����G��@��-}�ٿ$JS��"�@0��}�3@�G6�ʐ!?����G��@��-}�ٿ$JS��"�@0��}�3@�G6�ʐ!?����G��@|H~آٿ\*T�UD�@�q�3@��O	��!?��N6�@|H~آٿ\*T�UD�@�q�3@��O	��!?��N6�@|H~آٿ\*T�UD�@�q�3@��O	��!?��N6�@|H~آٿ\*T�UD�@�q�3@��O	��!?��N6�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@j8>u~�ٿ���?-��@/5o �3@)�9��!?a"�Jγ�@�A����ٿ����c�@�k��3@哖L��!?�[�E�@��'Тٿt�%�o��@����3@?�2Ð!?*��L��@멟Eߢٿ��%�[��@�k`�k�3@ �b�!?E��J���@멟Eߢٿ��%�[��@�k`�k�3@ �b�!?E��J���@멟Eߢٿ��%�[��@�k`�k�3@ �b�!?E��J���@g%J��ٿ���A���@�.���3@��`��!?��@��@g%J��ٿ���A���@�.���3@��`��!?��@��@g%J��ٿ���A���@�.���3@��`��!?��@��@g%J��ٿ���A���@�.���3@��`��!?��@��@I_L=�ٿ|z�1t�@�e���3@-��q�!?��M�<�@I_L=�ٿ|z�1t�@�e���3@-��q�!?��M�<�@I_L=�ٿ|z�1t�@�e���3@-��q�!?��M�<�@I_L=�ٿ|z�1t�@�e���3@-��q�!?��M�<�@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@Z,�!(�ٿ�瀬���@T���3@��ݲ�!?�C�q��@��T͠ٿ�H��}��@ռ��3@�.�3��!?��n���@��T͠ٿ�H��}��@ռ��3@�.�3��!?��n���@{\�Y9�ٿ���X��@n�C]_�3@l޴��!?�S�C�9�@{\�Y9�ٿ���X��@n�C]_�3@l޴��!?�S�C�9�@{\�Y9�ٿ���X��@n�C]_�3@l޴��!?�S�C�9�@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@V���{�ٿ�hɍ�j�@�!#��3@X�X�ǐ!?�&�fp��@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@���֞ٿ��rt��@U���3@�$\�ː!?�$�l�@�}�j��ٿf�SOo�@��
��3@Ú�ː!?�����@�}�j��ٿf�SOo�@��
��3@Ú�ː!?�����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@�Ձn�ٿN�f�,�@F֦���3@�v����!?meh����@V]W�>�ٿC1,���@/��;��3@p�rs7�!?�'7��@V]W�>�ٿC1,���@/��;��3@p�rs7�!?�'7��@V]W�>�ٿC1,���@/��;��3@p�rs7�!?�'7��@����͞ٿ�((W��@pf|	�3@�a�Of�!?o�YF*�@���ٿu��~t��@\�tg�3@�Bgt$�!?e�={=�@���ٿu��~t��@\�tg�3@�Bgt$�!?e�={=�@�Q���ٿdE��g�@�e�U�3@<-�%�!?���R`�@�Q���ٿdE��g�@�e�U�3@<-�%�!?���R`�@�Q���ٿdE��g�@�e�U�3@<-�%�!?���R`�@�Q���ٿdE��g�@�e�U�3@<-�%�!?���R`�@�Q���ٿdE��g�@�e�U�3@<-�%�!?���R`�@�k&k�ٿ�-#��@1��d�3@��V�@�!?h��CG��@�k&k�ٿ�-#��@1��d�3@��V�@�!?h��CG��@�k&k�ٿ�-#��@1��d�3@��V�@�!?h��CG��@�k&k�ٿ�-#��@1��d�3@��V�@�!?h��CG��@�k&k�ٿ�-#��@1��d�3@��V�@�!?h��CG��@��ҕH�ٿ?H��>h�@{}�-�3@�zw��!?���v�@��ҕH�ٿ?H��>h�@{}�-�3@�zw��!?���v�@��ҕH�ٿ?H��>h�@{}�-�3@�zw��!?���v�@�_O��ٿ>�>����@ ��Z�3@��7�!?g,}6��@�_O��ٿ>�>����@ ��Z�3@��7�!?g,}6��@����1�ٿ2��^<��@c��R�3@'2K��!?K��j�.�@�f��ߘٿ������@:LX���3@�J�qŐ!?�;^�G�@>"H��ٿ��}+N��@���]�3@�����!?FE�)�@>"H��ٿ��}+N��@���]�3@�����!?FE�)�@>"H��ٿ��}+N��@���]�3@�����!?FE�)�@��$�I�ٿ��"�lt�@��~��3@��+\�!?K
�8�)�@��$�I�ٿ��"�lt�@��~��3@��+\�!?K
�8�)�@��$�I�ٿ��"�lt�@��~��3@��+\�!?K
�8�)�@��$�I�ٿ��"�lt�@��~��3@��+\�!?K
�8�)�@��$�I�ٿ��"�lt�@��~��3@��+\�!?K
�8�)�@�z�7�ٿ��K����@zoZ2��3@yS֐!?�h����@�z�7�ٿ��K����@zoZ2��3@yS֐!?�h����@�z�7�ٿ��K����@zoZ2��3@yS֐!?�h����@�z�7�ٿ��K����@zoZ2��3@yS֐!?�h����@�z�7�ٿ��K����@zoZ2��3@yS֐!?�h����@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@#�PMx�ٿ�m�!���@������3@T=Jǐ!?
 Z,��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@�0p��ٿW��p�@�A5��3@0��L��!?�ￜ��@;~�&�ٿ�����@�����3@�� ��!?ܪ�����@;~�&�ٿ�����@�����3@�� ��!?ܪ�����@;~�&�ٿ�����@�����3@�� ��!?ܪ�����@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@����j�ٿ��dt��@�aq�y�3@�1����!?7�o���@��ؘ��ٿ.�L��V�@�)�ד�3@7#�ސ!?��L�	�@��ؘ��ٿ.�L��V�@�)�ד�3@7#�ސ!?��L�	�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@gd�9X�ٿ�������@Z:)�I�3@��e��!?�~��v�@����ٿ�ڹx%��@�@S�3@JQ����!?6�o|]�@����ٿ�ڹx%��@�@S�3@JQ����!?6�o|]�@����ٿ�ڹx%��@�@S�3@JQ����!?6�o|]�@����ٿ�ڹx%��@�@S�3@JQ����!?6�o|]�@����ٿ�ڹx%��@�@S�3@JQ����!?6�o|]�@�8�w�ٿJ�9�P�@%����3@L1��Ґ!?Agt�p��@kkb?��ٿd���@���3R�3@�9��z�!?���6���@kkb?��ٿd���@���3R�3@�9��z�!?���6���@kkb?��ٿd���@���3R�3@�9��z�!?���6���@޽^���ٿ���D�@��\�3@W��Ґ!?��#�h��@
*�/�ٿ8#e��@�����3@PỠ��!?�f7,���@
*�/�ٿ8#e��@�����3@PỠ��!?�f7,���@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@S"f@��ٿ�&e[Yq�@�녙��3@�>�ΐ!?�K��x�@����ٿ5}#d��@�چ.��3@ܰ��!?��#O�@����ٿ5}#d��@�چ.��3@ܰ��!?��#O�@����ٿ5}#d��@�چ.��3@ܰ��!?��#O�@/��Q��ٿ/i��@Q���3@�����!?>xN���@/��Q��ٿ/i��@Q���3@�����!?>xN���@/��Q��ٿ/i��@Q���3@�����!?>xN���@Qh1d�ٿ��r���@�<�t��3@�,�ϐ!?�I!�@Qh1d�ٿ��r���@�<�t��3@�,�ϐ!?�I!�@Qh1d�ٿ��r���@�<�t��3@�,�ϐ!?�I!�@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@f�𮣠ٿ�� �;��@�����3@��̽ߐ!?�}���@��͂יٿ������@�l�n�3@b	�~��!?W�n�փ�@��͂יٿ������@�l�n�3@b	�~��!?W�n�փ�@���v�ٿ^@���[�@�����3@)�1���!?l���(��@���v�ٿ^@���[�@�����3@)�1���!?l���(��@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@	�J_'�ٿ�,��T2�@�hN�q�3@~揩��!?�.DC�m�@�%�Ϛٿj*�7��@X�M��3@�tNlڐ!?�V�T}�@�%�Ϛٿj*�7��@X�M��3@�tNlڐ!?�V�T}�@z0	�ٿ'�x��}�@��7��3@��z��!?=ը��%�@z0	�ٿ'�x��}�@��7��3@��z��!?=ը��%�@ÿ�3��ٿyv���@�6Z C�3@+r^�ΐ!?1�U+]^�@ÿ�3��ٿyv���@�6Z C�3@+r^�ΐ!?1�U+]^�@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@3Hˍ��ٿ�'m�@@V�׌�3@�^
��!?�7�P��@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@�ȅ%֡ٿ;$�o_h�@�����3@��S�!?��[��^�@^	���ٿ� Ȕ���@����/�3@S��S��!?�T9X�@^	���ٿ� Ȕ���@����/�3@S��S��!?�T9X�@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@;X�ٿQ�v�[�@k ����3@�`�亐!?�d4$1��@c%���ٿum3
S�@�#���3@�4��}�!?�*�Z1��@c%���ٿum3
S�@�#���3@�4��}�!?�*�Z1��@c%���ٿum3
S�@�#���3@�4��}�!?�*�Z1��@�K�@�ٿ�M����@6����3@�L�ِ!?|�D��@�K�@�ٿ�M����@6����3@�L�ِ!?|�D��@�K�@�ٿ�M����@6����3@�L�ِ!?|�D��@�K�@�ٿ�M����@6����3@�L�ِ!?|�D��@N 8��ٿ��8Ǳ[�@$����3@`�f�!?���y�@|��f�ٿ2�|���@5��R�3@uӞr�!?��5�N��@�'����ٿ?��Y~��@F�֣��3@t��W�!?�B}/�@�)��v�ٿ!�"��@eV����3@���V�!?�g���@�)��v�ٿ!�"��@eV����3@���V�!?�g���@�)��v�ٿ!�"��@eV����3@���V�!?�g���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���\��ٿE�R��@�e@6�3@4=7m�!?��Ɩ���@���z1�ٿp�AX��@� �/2�3@�n�預!?�?���@���z1�ٿp�AX��@� �/2�3@�n�預!?�?���@ȫ�ᮡٿd�	���@���Q�3@v ��ؐ!?[ ���@.�c��ٿF��Z�@7S����3@�L�k��!?o*���@.�c��ٿF��Z�@7S����3@�L�k��!?o*���@.�c��ٿF��Z�@7S����3@�L�k��!?o*���@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�L��£ٿ���Ŵ��@x~سw�3@v��0�!?�&�!j�@�sP��ٿ��~����@����>�3@�t6Y��!?Z���և�@wn;y�ٿϤ]e_��@��7��3@�SK��!?:�l+��@wn;y�ٿϤ]e_��@��7��3@�SK��!?:�l+��@wn;y�ٿϤ]e_��@��7��3@�SK��!?:�l+��@wn;y�ٿϤ]e_��@��7��3@�SK��!?:�l+��@R!��ٿ��!_���@���N��3@��뒜�!?�ZP���@R!��ٿ��!_���@���N��3@��뒜�!?�ZP���@R!��ٿ��!_���@���N��3@��뒜�!?�ZP���@���ᮦٿ��"���@��3��3@#T����!?��b��.�@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@RU���ٿ�ѽ�O��@G�w t�3@J�Ő!?cP�8��@�F�&��ٿ�5�>	�@�HЙ�3@��|��!?{.�F��@�2Q�*�ٿߧ���E�@'�sͦ�3@���!?��#H�@�2Q�*�ٿߧ���E�@'�sͦ�3@���!?��#H�@�2Q�*�ٿߧ���E�@'�sͦ�3@���!?��#H�@�2Q�*�ٿߧ���E�@'�sͦ�3@���!?��#H�@��[p�ٿ<�v�9��@'�f��3@�EJ���!?�J�DC�@��[p�ٿ<�v�9��@'�f��3@�EJ���!?�J�DC�@��[p�ٿ<�v�9��@'�f��3@�EJ���!?�J�DC�@L�Ux��ٿ����@"��)�3@���Ј�!?)3���@���V�ٿ<]���P�@�q6Q�3@C�P��!?P���?<�@���V�ٿ<]���P�@�q6Q�3@C�P��!?P���?<�@���V�ٿ<]���P�@�q6Q�3@C�P��!?P���?<�@���V�ٿ<]���P�@�q6Q�3@C�P��!?P���?<�@���V�ٿ<]���P�@�q6Q�3@C�P��!?P���?<�@A9���ٿ���m�@��{��3@�pҐ!?�K	�@A9���ٿ���m�@��{��3@�pҐ!?�K	�@A9���ٿ���m�@��{��3@�pҐ!?�K	�@A9���ٿ���m�@��{��3@�pҐ!?�K	�@A9���ٿ���m�@��{��3@�pҐ!?�K	�@�xQ.�ٿF�.0�@� P��3@ߩ���!?��!�*~�@�xQ.�ٿF�.0�@� P��3@ߩ���!?��!�*~�@�xQ.�ٿF�.0�@� P��3@ߩ���!?��!�*~�@�xQ.�ٿF�.0�@� P��3@ߩ���!?��!�*~�@?�����ٿLB%�=�@5����3@��u0Ð!?V�.�7�@?�����ٿLB%�=�@5����3@��u0Ð!?V�.�7�@?�����ٿLB%�=�@5����3@��u0Ð!?V�.�7�@?�����ٿLB%�=�@5����3@��u0Ð!?V�.�7�@vg����ٿ|ٲ�w�@�e��3@���{��!?_�	�bq�@vg����ٿ|ٲ�w�@�e��3@���{��!?_�	�bq�@vg����ٿ|ٲ�w�@�e��3@���{��!?_�	�bq�@�;�l�ٿi��D�s�@Ʌp3�3@�s�9��!?�6̞��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@2����ٿ+Z)��M�@H^�R:�3@�-���!?Q#�"'��@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�R`�$�ٿ�4l\��@("��3@3�q��!?@��J�@�����ٿ�뚦Q�@1����3@���)�!?��Нw�@�����ٿ�뚦Q�@1����3@���)�!?��Нw�@�����ٿ�뚦Q�@1����3@���)�!?��Нw�@�����ٿ�뚦Q�@1����3@���)�!?��Нw�@	Xc��ٿL��43�@h	\��3@ ,ʐ!?af08��@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@�\]sR�ٿ�����5�@����~�3@�L
j��!?�a��_�@v
�,��ٿ1�FI�%�@�QS�3@�Q\]�!?�%�����@v
�,��ٿ1�FI�%�@�QS�3@�Q\]�!?�%�����@v
�,��ٿ1�FI�%�@�QS�3@�Q\]�!?�%�����@v
�,��ٿ1�FI�%�@�QS�3@�Q\]�!?�%�����@v
�,��ٿ1�FI�%�@�QS�3@�Q\]�!?�%�����@ڷ,��ٿ��J��b�@;Q��3@�!�P`�!?�����@*��O�ٿPm��4�@da�Pb�3@V����!?�3���V�@*��O�ٿPm��4�@da�Pb�3@V����!?�3���V�@*��O�ٿPm��4�@da�Pb�3@V����!?�3���V�@*��O�ٿPm��4�@da�Pb�3@V����!?�3���V�@���_�ٿ�Di���@\L�N��3@dtN��!?�W���@���_�ٿ�Di���@\L�N��3@dtN��!?�W���@���_�ٿ�Di���@\L�N��3@dtN��!?�W���@���_�ٿ�Di���@\L�N��3@dtN��!?�W���@���_�ٿ�Di���@\L�N��3@dtN��!?�W���@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@��
3?�ٿ�.��Z�@����5�3@�5w��!?��/��M�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@����ٿ�'�:�N�@u��v��3@��w<�!?R�x�G�@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@ q.=a�ٿ�j~�� �@���J��3@�*֪֐!?<Q[���@}	�y�ٿ�,�\�@�h��3@ ��[��!?[��l��@Ke�n��ٿ���2]��@�a��3@]��S��!?���6�@����k�ٿbbMSa�@D��	��3@	��[�!?غ��M��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@hwx��ٿ�0<\F�@F���3@-&��!?����
��@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@!D�R��ٿl����@,�fM~�3@W/�pՐ!?2F>U���@#<��@�ٿq��E�u�@��xo*�3@�8W��!?_����@#<��@�ٿq��E�u�@��xo*�3@�8W��!?_����@#<��@�ٿq��E�u�@��xo*�3@�8W��!?_����@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@�����ٿ��R�G5�@�W)S��3@|:zȯ�!?�^�'���@.ܥy�ٿ�i�8g��@o�����3@b�]z�!?������@f �Ɲٿ�oA�%��@�(��s�3@�C]d��!?�\W�~��@f �Ɲٿ�oA�%��@�(��s�3@�C]d��!?�\W�~��@Je��Ӣٿ��UE��@��Ě��3@3�h̊�!?r��+��@Je��Ӣٿ��UE��@��Ě��3@3�h̊�!?r��+��@�}�d�ٿr��U0d�@���o��3@���_�!?��Sxf��@�}�d�ٿr��U0d�@���o��3@���_�!?��Sxf��@�}�d�ٿr��U0d�@���o��3@���_�!?��Sxf��@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@��L���ٿ�9b8C�@)�1���3@�Soc�!?�����@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@!���>�ٿiQMd��@�k����3@L��ǻ�!?�ڍ���@��cB9�ٿ����@�����3@_�&���!?#�L����@��cB9�ٿ����@�����3@_�&���!?#�L����@��cB9�ٿ����@�����3@_�&���!?#�L����@��cB9�ٿ����@�����3@_�&���!?#�L����@��cB9�ٿ����@�����3@_�&���!?#�L����@��cB9�ٿ����@�����3@_�&���!?#�L����@f�U���ٿH����&�@�-/��3@{�,!?�*w�� �@f�U���ٿH����&�@�-/��3@{�,!?�*w�� �@f�U���ٿH����&�@�-/��3@{�,!?�*w�� �@����w�ٿ�N,1��@W�%v3�3@�͍2�!?J{��c��@����w�ٿ�N,1��@W�%v3�3@�͍2�!?J{��c��@��'�ٿȌ�X���@�$��3@�\�W%�!?-�-���@�r�S�ٿ6#~�w�@�x	�L�3@LfJn�!?n��Er�@�r�S�ٿ6#~�w�@�x	�L�3@LfJn�!?n��Er�@�r�S�ٿ6#~�w�@�x	�L�3@LfJn�!?n��Er�@�r�S�ٿ6#~�w�@�x	�L�3@LfJn�!?n��Er�@tM�,�ٿA�A�ME�@�f�3@)BĐ!?\)��I�@tM�,�ٿA�A�ME�@�f�3@)BĐ!?\)��I�@tM�,�ٿA�A�ME�@�f�3@)BĐ!?\)��I�@tM�,�ٿA�A�ME�@�f�3@)BĐ!?\)��I�@tM�,�ٿA�A�ME�@�f�3@)BĐ!?\)��I�@w��¡ٿŨ�|5��@���V�3@��\\��!?�N��Qq�@w��¡ٿŨ�|5��@���V�3@��\\��!?�N��Qq�@w��¡ٿŨ�|5��@���V�3@��\\��!?�N��Qq�@w��¡ٿŨ�|5��@���V�3@��\\��!?�N��Qq�@����%�ٿ���#q�@�iĬ��3@��h�!?�y�v���@����%�ٿ���#q�@�iĬ��3@��h�!?�y�v���@����%�ٿ���#q�@�iĬ��3@��h�!?�y�v���@����%�ٿ���#q�@�iĬ��3@��h�!?�y�v���@TP�K�ٿ��;L��@|���7�3@Y@Y�!?M̌���@Ol��ٿ������@gt}�o�3@#,¤�!?�h5�*`�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@��8��ٿ���o_�@�r����3@˼���!?;���	�@�ڛ|�ٿ�����@�#˷w�3@r��I�!?h��6`�@�ڛ|�ٿ�����@�#˷w�3@r��I�!?h��6`�@�ڛ|�ٿ�����@�#˷w�3@r��I�!?h��6`�@A����ٿrFQ�L�@`��w��3@�z ��!?�� x��@A����ٿrFQ�L�@`��w��3@�z ��!?�� x��@A����ٿrFQ�L�@`��w��3@�z ��!?�� x��@A����ٿrFQ�L�@`��w��3@�z ��!?�� x��@a�KEd�ٿyS���@�ѡ���3@ )7�ސ!?K�~��@a�KEd�ٿyS���@�ѡ���3@ )7�ސ!?K�~��@a�KEd�ٿyS���@�ѡ���3@ )7�ސ!?K�~��@a�KEd�ٿyS���@�ѡ���3@ )7�ސ!?K�~��@a�KEd�ٿyS���@�ѡ���3@ )7�ސ!?K�~��@ͬP��ٿ�{DQ�+�@���;��3@Ҩ3���!?�� �9�@ͬP��ٿ�{DQ�+�@���;��3@Ҩ3���!?�� �9�@Ӎ�n�ٿ�6�_�#�@a2rr��3@<�(k�!?�7[��@Ӎ�n�ٿ�6�_�#�@a2rr��3@<�(k�!?�7[��@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@AU.�ٿ1��k�t�@d�T�3@��M.�!?NWW�>'�@Oz����ٿ��U~���@*AQ3#�3@�s�2�!?��P�2�@Oz����ٿ��U~���@*AQ3#�3@�s�2�!?��P�2�@Oz����ٿ��U~���@*AQ3#�3@�s�2�!?��P�2�@Oz����ٿ��U~���@*AQ3#�3@�s�2�!?��P�2�@m"��Ǣٿ��i�,�@x���!�3@�9VB�!?���T���@��U�t�ٿP��`��@E���l�3@�1B#�!?t�����@��U�t�ٿP��`��@E���l�3@�1B#�!?t�����@��U�t�ٿP��`��@E���l�3@�1B#�!?t�����@<��I�ٿ�>�TG��@y#��3@��gِ!?�������@<:��ٿX���j��@��6���3@������!?p�7<hV�@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@������ٿ&�
3��@�����3@l�ɐ!?I�����@�oš�ٿ:X�s���@̘}A�3@~Qu��!?�f)���@�oš�ٿ:X�s���@̘}A�3@~Qu��!?�f)���@�oš�ٿ:X�s���@̘}A�3@~Qu��!?�f)���@�oš�ٿ:X�s���@̘}A�3@~Qu��!?�f)���@�oš�ٿ:X�s���@̘}A�3@~Qu��!?�f)���@M�vb��ٿ��)�6��@�s���3@��%ϐ!?o����m�@c\��2�ٿ��q{E��@A <ؠ�3@��/���!?��ݖ2j�@A��աٿ�og%���@����3@�n����!?�<=�^��@�6M�ٿm<J�@�d��3@��d��!?0: �/��@�6M�ٿm<J�@�d��3@��d��!?0: �/��@�6M�ٿm<J�@�d��3@��d��!?0: �/��@�6M�ٿm<J�@�d��3@��d��!?0: �/��@�6M�ٿm<J�@�d��3@��d��!?0: �/��@�&��W�ٿ���o�@�=��3@��OP�!?��}cF�@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@@8{X��ٿlC�V��@V'�љ�3@:Q�!?��?�� �@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@������ٿ%ׇ��q�@�N1�3@�+�Ɛ!?+, ��@�#�ݪ�ٿ!�DU���@S gH#�3@nzJ?Ґ!?ĘOC;�@�#�ݪ�ٿ!�DU���@S gH#�3@nzJ?Ґ!?ĘOC;�@�ؘ��ٿV�����@��xI�3@�0&Đ!?��$|^�@�ؘ��ٿV�����@��xI�3@�0&Đ!?��$|^�@�ؘ��ٿV�����@��xI�3@�0&Đ!?��$|^�@�ؘ��ٿV�����@��xI�3@�0&Đ!?��$|^�@@u1o�ٿ,cTƔ�@��U�'�3@���[��!?%X�/:�@@u1o�ٿ,cTƔ�@��U�'�3@���[��!?%X�/:�@@u1o�ٿ,cTƔ�@��U�'�3@���[��!?%X�/:�@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@� Ή�ٿK�a����@C=`OV�3@��U�}�!?�x�F���@��ӕٿ��7+��@2Z�Z_�3@�	U���!?X�R �@��ӕٿ��7+��@2Z�Z_�3@�	U���!?X�R �@��ӕٿ��7+��@2Z�Z_�3@�	U���!?X�R �@�-�Q�ٿsLOV��@?��@M�3@�7_�4�!?ʺ]���@�ь�F�ٿ���j�@Q��3@oї��!?Y=q����@�^�ٿrc�,�_�@`�8���3@zobN�!?�ǔW��@"j#uڟٿ��&�6�@����
�3@rd"f�!?������@"j#uڟٿ��&�6�@����
�3@rd"f�!?������@oi�0�ٿ���,���@���7�3@b��*��!?�ul72��@�����ٿN��7[��@2�Q,�3@���Z��!?٢Zj��@�����ٿN��7[��@2�Q,�3@���Z��!?٢Zj��@�����ٿN��7[��@2�Q,�3@���Z��!?٢Zj��@�����ٿN��7[��@2�Q,�3@���Z��!?٢Zj��@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@
R)ٿ�;�����@�����3@�jpΐ!?��́.�@��驡ٿ�7����@��D�(�3@#��!?T\}�$�@��驡ٿ�7����@��D�(�3@#��!?T\}�$�@�'�ٿYty`VB�@g��J��3@��u�Ґ!?�*�S�@�'�ٿYty`VB�@g��J��3@��u�Ґ!?�*�S�@�'�ٿYty`VB�@g��J��3@��u�Ґ!?�*�S�@�"N��ٿ�i��@6|�F��3@�9mj�!?��ҁ�@�"N��ٿ�i��@6|�F��3@�9mj�!?��ҁ�@�����ٿe��pQ�@@�C��3@��vﲐ!?��m[̚�@�����ٿe��pQ�@@�C��3@��vﲐ!?��m[̚�@�����ٿe��pQ�@@�C��3@��vﲐ!?��m[̚�@�����ٿe��pQ�@@�C��3@��vﲐ!?��m[̚�@�����ٿe��pQ�@@�C��3@��vﲐ!?��m[̚�@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@,��\�ٿS�]���@��^�e�3@do�e�!?,�HX���@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@�H��ٿ>K"SV�@�XJ_�3@���!?;ȳ0��@ж���ٿv��@;��@��\TR�3@MQ����!?���!S�@ж���ٿv��@;��@��\TR�3@MQ����!?���!S�@t�J�٠ٿp�8���@�O��3@������!?e
J���@���d�ٿ���##�@d\�ty�3@����!?��L��@���d�ٿ���##�@d\�ty�3@����!?��L��@��
ƽ�ٿ-���,�@�y��3@o����!?�>�ޥ	�@�F�[t�ٿ���X��@��Y=v�3@i����!?쫰�%��@�Wzo��ٿy�|\7�@��%vw�3@nu���!?l�e�?k�@�Wzo��ٿy�|\7�@��%vw�3@nu���!?l�e�?k�@�Wzo��ٿy�|\7�@��%vw�3@nu���!?l�e�?k�@�Wzo��ٿy�|\7�@��%vw�3@nu���!?l�e�?k�@<e����ٿ�9-�@d��d$�3@3��L��!?�ɽ�Nh�@m&����ٿ�B�����@ ��Z��3@��y�!?����@m&����ٿ�B�����@ ��Z��3@��y�!?����@m&����ٿ�B�����@ ��Z��3@��y�!?����@�}�{�ٿ�+��kM�@����3@֕��h�!?ڐ����@�}�{�ٿ�+��kM�@����3@֕��h�!?ڐ����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@۠�4�ٿ/��.���@)�Ԑ�3@u-x���!?:�����@�Ϳ�3�ٿ���>��@1�A�&�3@#A�c��!?j���-�@���{�ٿ�Ѝ���@,�j���3@�˂Ր!?ArJ8��@��f���ٿ�ek��/�@#�z�U�3@Y���!?��+�jS�@��f���ٿ�ek��/�@#�z�U�3@Y���!?��+�jS�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@��zj�ٿa��7���@�����3@O,%�!?�^e� J�@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@�S��8�ٿ��H�7�@T���3@8����!?���@���	��ٿdU]�tc�@?�G=�3@�1�#b�!?�S�;,�@���	��ٿdU]�tc�@?�G=�3@�1�#b�!?�S�;,�@���	��ٿdU]�tc�@?�G=�3@�1�#b�!?�S�;,�@���	��ٿdU]�tc�@?�G=�3@�1�#b�!?�S�;,�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���6�ٿ��ɑ#��@3m"�D�3@v�}ة�!?��6h�@���ٿ���}]�@�T(��3@��ؐ!?E9 �n�@���ٿ���}]�@�T(��3@��ؐ!?E9 �n�@���ٿ���}]�@�T(��3@��ؐ!?E9 �n�@���ٿ���}]�@�T(��3@��ؐ!?E9 �n�@���ٿ���}]�@�T(��3@��ؐ!?E9 �n�@��~��ٿWH����@�6氚�3@�Z��Ð!?���Y{��@��~��ٿWH����@�6氚�3@�Z��Ð!?���Y{��@��~��ٿWH����@�6氚�3@�Z��Ð!?���Y{��@��~��ٿWH����@�6氚�3@�Z��Ð!?���Y{��@�%�K��ٿ|�����@1j�GD�3@�C�c�!?!�����@d���ٿZO��l�@L�Т��3@�����!?#�B�;�@d���ٿZO��l�@L�Т��3@�����!?#�B�;�@d���ٿZO��l�@L�Т��3@�����!?#�B�;�@d���ٿZO��l�@L�Т��3@�����!?#�B�;�@e�7	�ٿ�����@>��M3�3@��2��!?��6�y��@e�7	�ٿ�����@>��M3�3@��2��!?��6�y��@����F�ٿ!Q{����@59�x~�3@���Ő!?.H����@����F�ٿ!Q{����@59�x~�3@���Ő!?.H����@^P r��ٿA�y
�@�"uy��3@'l�j�!?�f{����@^P r��ٿA�y
�@�"uy��3@'l�j�!?�f{����@^P r��ٿA�y
�@�"uy��3@'l�j�!?�f{����@^P r��ٿA�y
�@�"uy��3@'l�j�!?�f{����@��F�ٿvm{���@.��-�3@������!?��7����@��F�ٿvm{���@.��-�3@������!?��7����@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@h���ٿ78��u�@>w�|�3@�9?@��!?��!�\��@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@K���ٿTLwp��@���'�3@�B�Ǿ�!?�O��m�@�uꍹ�ٿ�Y�xDT�@4�$]��3@;KΩ��!?��A��@º91̤ٿ����\��@�x���3@W���!?P��[q��@º91̤ٿ����\��@�x���3@W���!?P��[q��@º91̤ٿ����\��@�x���3@W���!?P��[q��@dCj	ݣٿ�^�j�@쫰~�3@���Ӑ!??j~qi��@dCj	ݣٿ�^�j�@쫰~�3@���Ӑ!??j~qi��@dCj	ݣٿ�^�j�@쫰~�3@���Ӑ!??j~qi��@e���ٿ)�M���@�p!.��3@8p��!?����O��@e���ٿ)�M���@�p!.��3@8p��!?����O��@f�=2�ٿ�p�7Qf�@�dJ��3@�Ʉ|�!?�:����@f�=2�ٿ�p�7Qf�@�dJ��3@�Ʉ|�!?�:����@;>��~�ٿ�I0�OZ�@�s�S�3@��� ��!?&�K��@;>��~�ٿ�I0�OZ�@�s�S�3@��� ��!?&�K��@;>��~�ٿ�I0�OZ�@�s�S�3@��� ��!?&�K��@��ٿ�2l�]��@闑��3@7�,ʣ�!?��
���@��ٿ�2l�]��@闑��3@7�,ʣ�!?��
���@��ٿ�2l�]��@闑��3@7�,ʣ�!?��
���@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�3��d�ٿ���έ�@�wn�i�3@�V���!?XO��7��@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�m�>ژٿh�R�:�@m�L��3@R�#N��!?�F�C���@�+j^�ٿL~R"s"�@�.�q��3@i�Wː!?���D��@�+j^�ٿL~R"s"�@�.�q��3@i�Wː!?���D��@u�Q<��ٿ�?3kEI�@���Y�3@s�C���!?i�"I��@u�Q<��ٿ�?3kEI�@���Y�3@s�C���!?i�"I��@��Gn�ٿ�؃ۮ?�@�xq3��3@�Y�ø�!?�Q�*���@��Gn�ٿ�؃ۮ?�@�xq3��3@�Y�ø�!?�Q�*���@�r�8�ٿ�ܜn�{�@Օ�p�3@w�+�!?�T�L)��@�r�8�ٿ�ܜn�{�@Օ�p�3@w�+�!?�T�L)��@�r�8�ٿ�ܜn�{�@Օ�p�3@w�+�!?�T�L)��@�r�8�ٿ�ܜn�{�@Օ�p�3@w�+�!?�T�L)��@�۹�)�ٿ|UT9�@G��}O�3@�Ƿ���!?�Q⟺��@�۹�)�ٿ|UT9�@G��}O�3@�Ƿ���!?�Q⟺��@�۹�)�ٿ|UT9�@G��}O�3@�Ƿ���!?�Q⟺��@�۹�)�ٿ|UT9�@G��}O�3@�Ƿ���!?�Q⟺��@u�snԢٿ5���L��@R"���3@k	0 ��!?E'����@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�[�?��ٿL]��D��@�٭N�3@�	򀭐!?�E�+���@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�X">�ٿ�U�:T�@M�Wd�3@�S��!?L�'��@�<'[��ٿ��W���@�
[~��3@ݡ��!?�G;z҉�@�<'[��ٿ��W���@�
[~��3@ݡ��!?�G;z҉�@���䔡ٿC����@�<���3@Lb�{�!?���L�@���䔡ٿC����@�<���3@Lb�{�!?���L�@���䔡ٿC����@�<���3@Lb�{�!?���L�@���䔡ٿC����@�<���3@Lb�{�!?���L�@���䔡ٿC����@�<���3@Lb�{�!?���L�@[t��ٿ�wk�!z�@���>�3@ۖٱ��!?������@[t��ٿ�wk�!z�@���>�3@ۖٱ��!?������@[t��ٿ�wk�!z�@���>�3@ۖٱ��!?������@w-���ٿ<�W\��@y9�U<�3@-K8�̐!?|C�<�@w-���ٿ<�W\��@y9�U<�3@-K8�̐!?|C�<�@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@;a��ٿ~�"?Z?�@J®� �3@K�W��!?)Pȷ��@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@���ٿW������@n׸��3@����!?�V
���@ ���Νٿ]}����@f��3@��cV��!?��Y���@܊1���ٿɈ�&h�@�ah��3@�iJ~��!?P[D>��@܊1���ٿɈ�&h�@�ah��3@�iJ~��!?P[D>��@/���ٿ�q|]��@����3@|�쏐!?$H��{�@/���ٿ�q|]��@����3@|�쏐!?$H��{�@/���ٿ�q|]��@����3@|�쏐!?$H��{�@/���ٿ�q|]��@����3@|�쏐!?$H��{�@/���ٿ�q|]��@����3@|�쏐!?$H��{�@��8�ٿA͈"s��@���_�3@��򍌐!?D�#���@,-�8��ٿI�$�zC�@l%����3@�->�!?��3͙��@I��%Q�ٿݝ�M��@�"�Y��3@a�;ǐ!?��@I��%Q�ٿݝ�M��@�"�Y��3@a�;ǐ!?��@I��%Q�ٿݝ�M��@�"�Y��3@a�;ǐ!?��@I��%Q�ٿݝ�M��@�"�Y��3@a�;ǐ!?��@I��%Q�ٿݝ�M��@�"�Y��3@a�;ǐ!?��@�iKI�ٿ$���@���#T�3@O�C�!?vIG���@�iKI�ٿ$���@���#T�3@O�C�!?vIG���@�� �ٿ5ۖ���@;���3@���E��!?�Ea��@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@p�~
�ٿr ����@��ٿ��3@"4�ې!?ª�y���@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@y��\�ٿi�̐��@2ZD���3@P�l�!?Y	{�@�S����ٿ�4 %�@��ұ{�3@�frz�!?���g���@z�/�ٿLb�2�N�@�@|���3@͠���!?,�� @v�@z�/�ٿLb�2�N�@�@|���3@͠���!?,�� @v�@�X-�Ӝٿ$�*��@D��g��3@��[���!?/��S��@Gp���ٿ광F���@�p}��3@�'�<�!?����`Z�@Gp���ٿ광F���@�p}��3@�'�<�!?����`Z�@/���ٿ�����K�@��Lڿ�3@����ʐ!?/���y�@/���ٿ�����K�@��Lڿ�3@����ʐ!?/���y�@/���ٿ�����K�@��Lڿ�3@����ʐ!?/���y�@ƌJ��ٿ�GE�ơ�@��Z��3@_Ư�!?������@ƌJ��ٿ�GE�ơ�@��Z��3@_Ư�!?������@ƌJ��ٿ�GE�ơ�@��Z��3@_Ư�!?������@ᵾ9�ٿ�������@�AJ{�3@�"X|��!?�h"���@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@��ac�ٿ�"�����@�����3@0๓��!?Z�T'k(�@�L�9ԣٿUA�y�@�O�B��3@>��Ð!?3�3��@�L�9ԣٿUA�y�@�O�B��3@>��Ð!?3�3��@��׽��ٿ�H�|0��@��V�3@Kc��ΐ!?cʑ��C�@��׽��ٿ�H�|0��@��V�3@Kc��ΐ!?cʑ��C�@��׽��ٿ�H�|0��@��V�3@Kc��ΐ!?cʑ��C�@ER�d��ٿKlFI���@��"~ 4@̀�ݐ!?�<-|P�@4S�A��ٿ B/�0�@���R��3@C(���!?aLd���@4S�A��ٿ B/�0�@���R��3@C(���!?aLd���@S����ٿԻ�����@�KT�3@K�57�!?Ij�����@S����ٿԻ�����@�KT�3@K�57�!?Ij�����@1OnեٿDa<�@�m|d��3@�Z^ѐ!?��H��@�@1OnեٿDa<�@�m|d��3@�Z^ѐ!?��H��@�@1OnեٿDa<�@�m|d��3@�Z^ѐ!?��H��@�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@�=����ٿ�H_� �@�����3@xN��!?"]om�@��m���ٿ	�m�S�@��i��3@{I�¼�!?��o�@�zjѹ�ٿ����E�@�`�x��3@�}5�!?�� �Ϙ�@4T�0�ٿ��U�:h�@����w�3@��el!?��9���@K��1�ٿSuhZ���@�����3@v�#m��!?!�l�m��@K��1�ٿSuhZ���@�����3@v�#m��!?!�l�m��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@a�#!�ٿ�~�z+�@F��@�3@�h\�!?1%��@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@@`1�ٿb��.�@����g�3@������!?}-�5 E�@'{V�4�ٿ���L-�@����}�3@�AL8��!?�:"2��@D��ٿ=P�0*��@�0�.�3@�?!�!?������@D��ٿ=P�0*��@�0�.�3@�?!�!?������@D��ٿ=P�0*��@�0�.�3@�?!�!?������@D��ٿ=P�0*��@�0�.�3@�?!�!?������@D��ٿ=P�0*��@�0�.�3@�?!�!?������@D��ٿ=P�0*��@�0�.�3@�?!�!?������@�R/��ٿdF((��@�P�#��3@�Q�m�!?!���@�R/��ٿdF((��@�P�#��3@�Q�m�!?!���@�R/��ٿdF((��@�P�#��3@�Q�m�!?!���@�R/��ٿdF((��@�P�#��3@�Q�m�!?!���@�R/��ٿdF((��@�P�#��3@�Q�m�!?!���@�
�2�ٿ=��)���@��t���3@�N�K�!?�h �d��@�
�2�ٿ=��)���@��t���3@�N�K�!?�h �d��@RY�\V�ٿ<�����@�z����3@8'��Ԑ!?[�/�@����ٿW?.x��@9�i�3@j�p=ߐ!?��Ч�@�1�ٿk�hA�@����U�3@��lO�!?Yb�i�@�1�ٿk�hA�@����U�3@��lO�!?Yb�i�@�1�ٿk�hA�@����U�3@��lO�!?Yb�i�@�1�ٿk�hA�@����U�3@��lO�!?Yb�i�@�1�ٿk�hA�@����U�3@��lO�!?Yb�i�@�+��ٿ��q�c��@��h���3@�n�U��!?� S�O�@�+��ٿ��q�c��@��h���3@�n�U��!?� S�O�@�+��ٿ��q�c��@��h���3@�n�U��!?� S�O�@�+��ٿ��q�c��@��h���3@�n�U��!?� S�O�@�+��ٿ��q�c��@��h���3@�n�U��!?� S�O�@�J�K �ٿ?=E'�@�����3@��`.�!?M��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@VuB�ٿ�=�`l��@�:��4@�Ҿ���!?9�e��@s�m/r�ٿOI��@H�_�3@�M���!?k�����@s�m/r�ٿOI��@H�_�3@�M���!?k�����@X���ٿҽ%�Z�@�����3@��A��!?4B]�j�@X���ٿҽ%�Z�@�����3@��A��!?4B]�j�@:����ٿg��H\g�@P߾!��3@�e���!?��*A�@:����ٿg��H\g�@P߾!��3@�e���!?��*A�@���(�ٿ��؄���@~	6x��3@o[�S�!?|�UU���@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@P��ϟٿ��),���@��BFi�3@���a�!?�S�#!�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@�	&���ٿ��(%�@�-�j
�3@Ỳ��!?P���x�@*�.��ٿ�U�����@�T���3@����+�!?���ZB�@*�.��ٿ�U�����@�T���3@����+�!?���ZB�@vYJ�2�ٿ!��5�_�@����l�3@����!?��c�4��@vYJ�2�ٿ!��5�_�@����l�3@����!?��c�4��@�h(�O�ٿ���:J�@ų��3@���%��!?AdU�@�h(�O�ٿ���:J�@ų��3@���%��!?AdU�@�h(�O�ٿ���:J�@ų��3@���%��!?AdU�@�h(�O�ٿ���:J�@ų��3@���%��!?AdU�@�h(�O�ٿ���:J�@ų��3@���%��!?AdU�@V� ���ٿ�[��؆�@N���3@CU�~�!?8e��5S�@V� ���ٿ�[��؆�@N���3@CU�~�!?8e��5S�@V� ���ٿ�[��؆�@N���3@CU�~�!?8e��5S�@V� ���ٿ�[��؆�@N���3@CU�~�!?8e��5S�@V� ���ٿ�[��؆�@N���3@CU�~�!?8e��5S�@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�*;�ٿ�$����@��8�3@���_W�!?9˗�Q��@�%Dy��ٿ���(��@�ڤ�@�3@��~�!�!?WA���@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@'�GL��ٿz�^5��@�#z�3@q�cސ!?�e��\%�@��C���ٿ�&Y��@н��3@�#�ې!?���'�@��C���ٿ�&Y��@н��3@�#�ې!?���'�@��C���ٿ�&Y��@н��3@�#�ې!?���'�@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@X~�v"�ٿ��S�[�@g�	js�3@�?��!?�D�r"��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@d}QN��ٿ�ʳs���@�rQ���3@�|T��!?"hqm��@��r��ٿ�j:���@���<�3@g��"��!?ͱ���T�@��r��ٿ�j:���@���<�3@g��"��!?ͱ���T�@��r��ٿ�j:���@���<�3@g��"��!?ͱ���T�@���ٿ����q�@H �t�3@��е�!?"�� ��@���ٿ����q�@H �t�3@��е�!?"�� ��@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@���R)�ٿ#�hƉ��@�����3@X�xo��!?&]�6���@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@q��4�ٿ-S��_��@Go���3@W�ソ�!?����:�@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@�@����ٿ[�N+��@�}��3@�ͼ��!?+g[c��@q:�ٿn�Q�N�@}��dH�3@l�ې!?�[$�Z�@q:�ٿn�Q�N�@}��dH�3@l�ې!?�[$�Z�@q:�ٿn�Q�N�@}��dH�3@l�ې!?�[$�Z�@q:�ٿn�Q�N�@}��dH�3@l�ې!?�[$�Z�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@����{�ٿ�s�6�W�@��V+�3@��]��!?L�&�#=�@ܭR��ٿ����<��@��kS�3@{4�"|�!?n��}��@ܭR��ٿ����<��@��kS�3@{4�"|�!?n��}��@ܭR��ٿ����<��@��kS�3@{4�"|�!?n��}��@ܭR��ٿ����<��@��kS�3@{4�"|�!?n��}��@ܭR��ٿ����<��@��kS�3@{4�"|�!?n��}��@�ȍ�:�ٿyz��-��@��>�3@�b�t��!?E0=����@�ȍ�:�ٿyz��-��@��>�3@�b�t��!?E0=����@
8��ٿc[���@[.u��3@�U3}��!?��es��@$�j���ٿQZ����@��1K�3@�0|��!?d\���@$�j���ٿQZ����@��1K�3@�0|��!?d\���@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@p�V�q�ٿ���	�1�@��f�3@!�y��!?��fV��@Ϲ���ٿ�Z��@L��3@��Rν�!?]J'�'�@Ϲ���ٿ�Z��@L��3@��Rν�!?]J'�'�@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��^��ٿ�S�NQ6�@h\ ��3@��a^��!?�Eo��@��y�N�ٿ�:ȫ�@�1���3@��d���!?0Y���l�@��y�N�ٿ�:ȫ�@�1���3@��d���!?0Y���l�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@ƌ�W�ٿ�..���@�`%G=�3@��@Ð!?�h���/�@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@s�Fq�ٿb�#��@�Ot�
�3@H
�㮐!?�I��K��@J�L�ٿ�0N
���@7u�K[�3@�@����!?��ss�@J�L�ٿ�0N
���@7u�K[�3@�@����!?��ss�@J�L�ٿ�0N
���@7u�K[�3@�@����!?��ss�@J�L�ٿ�0N
���@7u�K[�3@�@����!?��ss�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@�ҍ�k�ٿpy;����@'\���3@�@4�!?���+ U�@M�; z�ٿF�/��@=��S��3@Zm-s�!?� Voʕ�@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@z��s�ٿ�5d��@�̵�� 4@$L�y�!?�4����@DQ]*ݡٿ�������@��cG�3@�u����!?&�g��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@h���Ԣٿ��p��@�����3@���x�!?mϴ_��@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@m�6@�ٿ�)��R�@%����3@�#Y ��!?Lp����@��ٿ�������@'F����3@��WK��!?%�5f�@��ٿ�������@'F����3@��WK��!?%�5f�@��ٿ�������@'F����3@��WK��!?%�5f�@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@O����ٿ4�����@��^�:�3@{u�ܐ!?Ue�R��@��k���ٿȫ����@��֤a�3@^�֥ɐ!?==jO���@��k���ٿȫ����@��֤a�3@^�֥ɐ!?==jO���@��k���ٿȫ����@��֤a�3@^�֥ɐ!?==jO���@��fh�ٿ&g绀t�@4�铺�3@q��!?9?��;�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@�9Y�u�ٿ\���L�@&!��+�3@m�ّ�!?+ߡ�l�@f���ٿ^��Q�7�@���9��3@��ʧ�!?℃�n�@f���ٿ^��Q�7�@���9��3@��ʧ�!?℃�n�@f���ٿ^��Q�7�@���9��3@��ʧ�!?℃�n�@f���ٿ^��Q�7�@���9��3@��ʧ�!?℃�n�@f���ٿ^��Q�7�@���9��3@��ʧ�!?℃�n�@�<�S��ٿ�� GO��@�3��y�3@N]N��!?������@�<�S��ٿ�� GO��@�3��y�3@N]N��!?������@�<�S��ٿ�� GO��@�3��y�3@N]N��!?������@]���ٿ�6�k�@�:����3@��S��!?�룢��@]���ٿ�6�k�@�:����3@��S��!?�룢��@]���ٿ�6�k�@�:����3@��S��!?�룢��@]���ٿ�6�k�@�:����3@��S��!?�룢��@]���ٿ�6�k�@�:����3@��S��!?�룢��@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@���ٿ��ۍ��@dw�,7�3@��@���!?�	���@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@��:F�ٿ��|��@m��2��3@3M?���!?^��kT��@nG�e��ٿ��[�:�@�����3@�$`��!?o�.�R(�@nG�e��ٿ��[�:�@�����3@�$`��!?o�.�R(�@U�~�m�ٿ�h�@��r�3@�5]tؐ!?������@G���8�ٿ2}Yb��@�k�y�3@z]�D�!?�#�n�@�'%V�ٿᝃk���@�e�r�3@���%�!?�x���e�@d�Q���ٿ��W��@H���m�3@AO�s�!?Y9R��@d�Q���ٿ��W��@H���m�3@AO�s�!?Y9R��@d�Q���ٿ��W��@H���m�3@AO�s�!?Y9R��@�Q�s�ٿ�U4��@�/On��3@d��uP�!?�J����@�Q�s�ٿ�U4��@�/On��3@d��uP�!?�J����@�Q�s�ٿ�U4��@�/On��3@d��uP�!?�J����@�3O�L�ٿ�uu����@�T��e�3@&#�cW�!?n@B���@}ޞ���ٿ�i�+�@*��.Q�3@�u[m�!?�hԚ���@}ޞ���ٿ�i�+�@*��.Q�3@�u[m�!?�hԚ���@}ޞ���ٿ�i�+�@*��.Q�3@�u[m�!?�hԚ���@}ޞ���ٿ�i�+�@*��.Q�3@�u[m�!?�hԚ���@x�(i��ٿ�M�A��@��C��3@�n�p�!?Fh�/i�@x�(i��ٿ�M�A��@��C��3@�n�p�!?Fh�/i�@x�(i��ٿ�M�A��@��C��3@�n�p�!?Fh�/i�@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@i��P�ٿ������@�s��3@IHam��!?��S5��@���ٿ�=�+w�@CH����3@�Ej�e�!?�u�C��@���ٿ�=�+w�@CH����3@�Ej�e�!?�u�C��@~���ٿ��}�~�@9#��Q�3@L���ݐ!?�ᐿ�+�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�T+�9�ٿ\6l�@�X�q2�3@��I���!?9���X/�@�.}
�ٿ�y��@ӹ��3@�CD�Ő!?���P��@�.}
�ٿ�y��@ӹ��3@�CD�Ő!?���P��@�.}
�ٿ�y��@ӹ��3@�CD�Ő!?���P��@�.}
�ٿ�y��@ӹ��3@�CD�Ő!?���P��@�.}
�ٿ�y��@ӹ��3@�CD�Ő!?���P��@���ۧ�ٿ�����@{�߿��3@	��甐!?�t;�4�@���ۧ�ٿ�����@{�߿��3@	��甐!?�t;�4�@���ۧ�ٿ�����@{�߿��3@	��甐!?�t;�4�@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@�QeN�ٿ�$��7��@�FU��3@`-��!?�3ix��@,E]뎞ٿB� 3��@2͝��3@Ѫ5�!?��:��@,E]뎞ٿB� 3��@2͝��3@Ѫ5�!?��:��@,E]뎞ٿB� 3��@2͝��3@Ѫ5�!?��:��@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@!�^Cc�ٿh5�+~��@?�O�7�3@=��s��!?���{�@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@��_�"�ٿ/.��b�@úL#��3@�X�G�!?�fe��@:1:��ٿx�6�Vf�@��n|E�3@��{���!?:�	0���@:1:��ٿx�6�Vf�@��n|E�3@��{���!?:�	0���@:1:��ٿx�6�Vf�@��n|E�3@��{���!?:�	0���@:1:��ٿx�6�Vf�@��n|E�3@��{���!?:�	0���@W|u�1�ٿ�j9�	�@�$J0,�3@���!?��Q�r��@W|u�1�ٿ�j9�	�@�$J0,�3@���!?��Q�r��@��i6��ٿO��ҁ�@�	a/��3@P>��z�!?g�l��@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@���^��ٿL��S�@C�P�3@�+|�y�!?�X���@����ٿ��4��@WBP"��3@�n�Ӑ!?���-AM�@����ٿ��4��@WBP"��3@�n�Ӑ!?���-AM�@����ٿ��4��@WBP"��3@�n�Ӑ!?���-AM�@����ٿ��4��@WBP"��3@�n�Ӑ!?���-AM�@����ٿ��4��@WBP"��3@�n�Ӑ!?���-AM�@��jl�ٿ�Zu
y��@�!P�3@�v/Ɛ!?�)h�\��@��jl�ٿ�Zu
y��@�!P�3@�v/Ɛ!?�)h�\��@��jl�ٿ�Zu
y��@�!P�3@�v/Ɛ!?�)h�\��@��jl�ٿ�Zu
y��@�!P�3@�v/Ɛ!?�)h�\��@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@�բ�ٿ�����@�i�3@Jv�!?�� JHp�@,5�
*�ٿX����r�@kԤk��3@��L�H�!?����Q�@G]���ٿ�B-0
1�@($�_F�3@L����!?
H�r��@G]���ٿ�B-0
1�@($�_F�3@L����!?
H�r��@G]���ٿ�B-0
1�@($�_F�3@L����!?
H�r��@����ٿL/܆`��@uo5��3@;Y����!?uu4J�@����ٿL/܆`��@uo5��3@;Y����!?uu4J�@����ٿL/܆`��@uo5��3@;Y����!?uu4J�@����ٿL/܆`��@uo5��3@;Y����!?uu4J�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@&�we�ٿ����X��@r���3@��M��!?��}�g�@BpVw�ٿ��(���@�K�3@�o��!?��P*���@������ٿf=X�=��@6uI�3@~�Zq��!?dHw灿�@������ٿf=X�=��@6uI�3@~�Zq��!?dHw灿�@������ٿf=X�=��@6uI�3@~�Zq��!?dHw灿�@������ٿf=X�=��@6uI�3@~�Zq��!?dHw灿�@������ٿf=X�=��@6uI�3@~�Zq��!?dHw灿�@����ٿ	��P��@��e�3@�^��!?�Ƈ���@����ٿ	��P��@��e�3@�^��!?�Ƈ���@$��b�ٿ?�O\��@�Nٗ��3@P=�c�!?��uP���@����%�ٿ}t�&���@N���3@��訐!?sw��ZY�@����%�ٿ}t�&���@N���3@��訐!?sw��ZY�@μL*h�ٿ�y���@���\�3@
�3���!?�!��L�@μL*h�ٿ�y���@���\�3@
�3���!?�!��L�@���ٿ]���@�F�$H�3@�d���!?�������@���ٿ]���@�F�$H�3@�d���!?�������@���ٿ]���@�F�$H�3@�d���!?�������@$�*P�ٿH���k�@ڝ�r>�3@̥2�͐!?�隲=��@$�*P�ٿH���k�@ڝ�r>�3@̥2�͐!?�隲=��@$�*P�ٿH���k�@ڝ�r>�3@̥2�͐!?�隲=��@$�*P�ٿH���k�@ڝ�r>�3@̥2�͐!?�隲=��@$�*P�ٿH���k�@ڝ�r>�3@̥2�͐!?�隲=��@iį|��ٿ|����%�@�bm�$�3@�i*�!?����`_�@iį|��ٿ|����%�@�bm�$�3@�i*�!?����`_�@iį|��ٿ|����%�@�bm�$�3@�i*�!?����`_�@iį|��ٿ|����%�@�bm�$�3@�i*�!?����`_�@����U�ٿܜ�pi�@�a�k��3@�}��Ő!?۔����@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@U���ٿ���l��@C�5� �3@�ԄI��!?�RQj���@2�ۋ�ٿ�YF��K�@�@D-�3@���+��!?���S���@2�ۋ�ٿ�YF��K�@�@D-�3@���+��!?���S���@V�3d�ٿ�W)x3��@D�pCR�3@��f`�!?�:�5�5�@V�3d�ٿ�W)x3��@D�pCR�3@��f`�!?�:�5�5�@V�3d�ٿ�W)x3��@D�pCR�3@��f`�!?�:�5�5�@V�3d�ٿ�W)x3��@D�pCR�3@��f`�!?�:�5�5�@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@��� �ٿ�cRB�5�@��h�3@BͣE��!?YzP���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@o��m �ٿPm����@�m؈b�3@EҞ�!?�W_���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@�+o�6�ٿ�z]�{��@��{b�3@�����!?�6�}���@{�n��ٿ��*���@q����3@��'�Ր!?w�����@{�n��ٿ��*���@q����3@��'�Ր!?w�����@{�n��ٿ��*���@q����3@��'�Ր!?w�����@{�n��ٿ��*���@q����3@��'�Ր!?w�����@{�n��ٿ��*���@q����3@��'�Ր!?w�����@�-lڠٿ��N�@��#U�3@크�ې!?_����@�-lڠٿ��N�@��#U�3@크�ې!?_����@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@o��[;�ٿIWdp<��@��3@Q,��!?v�c:��@��2B�ٿ�� ͇7�@Ϊ��k�3@���8�!?�����@��2B�ٿ�� ͇7�@Ϊ��k�3@���8�!?�����@��T_�ٿN ����@E����3@@!v˺�!?Ƶ����@��T_�ٿN ����@E����3@@!v˺�!?Ƶ����@��T_�ٿN ����@E����3@@!v˺�!?Ƶ����@i�+_[�ٿ���Nc�@8� �S�3@��Uݐ!?`���d�@i�+_[�ٿ���Nc�@8� �S�3@��Uݐ!?`���d�@�5N�g�ٿ�r.,���@�t�9\�3@��Eo��!?vQ.�L�@�5N�g�ٿ�r.,���@�t�9\�3@��Eo��!?vQ.�L�@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@��K?��ٿC���l�@kB���3@.P*��!?~'����@RNz*�ٿ ����@�`���3@����Ր!?�n�U�@RNz*�ٿ ����@�`���3@����Ր!?�n�U�@RNz*�ٿ ����@�`���3@����Ր!?�n�U�@T��o�ٿN8�)<�@/��p�3@�k~��!?�3U���@T��o�ٿN8�)<�@/��p�3@�k~��!?�3U���@��s�%�ٿ�0Jy��@
�|���3@蒂S�!?~�l �!�@l�T;�ٿ���ˌ��@)�r�3@[����!?[�oH�?�@l�T;�ٿ���ˌ��@)�r�3@[����!?[�oH�?�@l�T;�ٿ���ˌ��@)�r�3@[����!?[�oH�?�@�Fiޚٿ&d���@f%S���3@u�rWΐ!?FJ�ή��@b�f�ٿl�+�X�@����j�3@>5����!?���Tq�@b�f�ٿl�+�X�@����j�3@>5����!?���Tq�@b�f�ٿl�+�X�@����j�3@>5����!?���Tq�@b�f�ٿl�+�X�@����j�3@>5����!?���Tq�@��ȅt�ٿ:(KƱk�@����3@8���ϐ!?� ߁�~�@��ȅt�ٿ:(KƱk�@����3@8���ϐ!?� ߁�~�@��ȅt�ٿ:(KƱk�@����3@8���ϐ!?� ߁�~�@�x��ٿKgi���@�]����3@�:�`�!?@=�O���@eqh#�ٿ��yHҕ�@�� ��3@D��֐!?Y�Yd�>�@eqh#�ٿ��yHҕ�@�� ��3@D��֐!?Y�Yd�>�@eqh#�ٿ��yHҕ�@�� ��3@D��֐!?Y�Yd�>�@eqh#�ٿ��yHҕ�@�� ��3@D��֐!?Y�Yd�>�@�k���ٿ������@���J�3@��1!?9�QG�@�k���ٿ������@���J�3@��1!?9�QG�@�k���ٿ������@���J�3@��1!?9�QG�@�k���ٿ������@���J�3@��1!?9�QG�@���m�ٿX����Q�@�iE��3@��*ݐ�!?g�DD���@���m�ٿX����Q�@�iE��3@��*ݐ�!?g�DD���@�*E�ٿ���;��@�}�u�3@?_sﺐ!?��C�L�@ń�ٿ��R�i%�@A+-��3@13'��!?��S�2�@����ٿ���%D�@��g3%�3@�����!?�@m-�O�@����ٿ���%D�@��g3%�3@�����!?�@m-�O�@����ٿ���%D�@��g3%�3@�����!?�@m-�O�@����ٿ���%D�@��g3%�3@�����!?�@m-�O�@t�C���ٿ# ��D�@L���Y�3@4� i��!?���(�:�@t�C���ٿ# ��D�@L���Y�3@4� i��!?���(�:�@��k�ٿ���3��@�m�0�3@��q���!?�p�����@��k�ٿ���3��@�m�0�3@��q���!?�p�����@��k�ٿ���3��@�m�0�3@��q���!?�p�����@��k�ٿ���3��@�m�0�3@��q���!?�p�����@��k�ٿ���3��@�m�0�3@��q���!?�p�����@��k�ٿ���3��@�m�0�3@��q���!?�p�����@XY�
��ٿ/p�+�y�@�,���3@�ZM��!?.K,b���@XY�
��ٿ/p�+�y�@�,���3@�ZM��!?.K,b���@XY�
��ٿ/p�+�y�@�,���3@�ZM��!?.K,b���@XY�
��ٿ/p�+�y�@�,���3@�ZM��!?.K,b���@J�N�ٿ��O� �@kB�x�3@ݕo���!?A9�	��@J�N�ٿ��O� �@kB�x�3@ݕo���!?A9�	��@J�N�ٿ��O� �@kB�x�3@ݕo���!?A9�	��@mO�b��ٿ�����@II���3@�o4���!?rO�$�W�@mO�b��ٿ�����@II���3@�o4���!?rO�$�W�@mO�b��ٿ�����@II���3@�o4���!?rO�$�W�@���;��ٿ��;�`�@�z���3@Pdi��!?$ZQ��V�@���;��ٿ��;�`�@�z���3@Pdi��!?$ZQ��V�@��aF�ٿ��⁡��@b�PSE�3@��r���!?��pW�(�@��aF�ٿ��⁡��@b�PSE�3@��r���!?��pW�(�@��aF�ٿ��⁡��@b�PSE�3@��r���!?��pW�(�@!t��ٿ$5��@,��	�3@�|R���!?M NJ�6�@��H�Q�ٿ�v*=f��@�q�=M�3@�K���!?�n���@��H�Q�ٿ�v*=f��@�q�=M�3@�K���!?�n���@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@��'��ٿFw�W�@@=p��3@q嵾�!?���p�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@�D�#�ٿ}�9���@q�"��3@�^2��!?]w_�7�@���ٿ��/#�@�Tb���3@v Ϋΐ!?ք��z��@���ٿ��/#�@�Tb���3@v Ϋΐ!?ք��z��@.�W�ٿW$qJG�@�k��V�3@�|� ��!?۶T��~�@.�W�ٿW$qJG�@�k��V�3@�|� ��!?۶T��~�@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@�{X:��ٿ��@H�}�3@:��v�!?�p�,l��@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@rz"y.�ٿ��C��@�*Ar�3@� ��]�!?�eؠnh�@g��ʞ�ٿ��0����@�4W�B�3@Dr��!?�����)�@g��ʞ�ٿ��0����@�4W�B�3@Dr��!?�����)�@g��ʞ�ٿ��0����@�4W�B�3@Dr��!?�����)�@M�W%�ٿ����g�@]����3@������!?�')���@M�W%�ٿ����g�@]����3@������!?�')���@M�W%�ٿ����g�@]����3@������!?�')���@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@=`�K�ٿ�����j�@�Ơ�z�3@l���Ȑ!?}'�{�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@���o��ٿ܄!K���@*~�R��3@˂:��!?
:��R�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@X�:���ٿqq�=^�@��{iM�3@4݆�m�!?+k��v�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@��#Y�ٿ1�̣���@��@���3@12�K��!?�B�~�@����ٿ>El����@�h����3@s*Ӑ!?\ী��@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@N�+��ٿ�=����@<7�q�3@�QZJ��!?Hg[ם:�@����ٿ�%�Kd��@zA���3@`îӋ�!?�)y7��@
�uh�ٿ��+���@M�c��3@p�(��!?��>Jj��@
�uh�ٿ��+���@M�c��3@p�(��!?��>Jj��@Mq��Z�ٿ�[��@�#`��3@�
���!?x�wj3��@39yNǝٿ s|���@�ϴ��3@[�$硐!?����=�@39yNǝٿ s|���@�ϴ��3@[�$硐!?����=�@39yNǝٿ s|���@�ϴ��3@[�$硐!?����=�@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@�
��ݞٿ�ɶm_��@��W�p4@	��!?H��g���@e%���ٿ��?�s�@ϰ����3@�����!?�ՌY,��@�^����ٿk'���4�@��&(�3@'Хlg�!?��	����@�Ar�>�ٿ��?��@s[Hr��3@��]^�!?�O��@�Ar�>�ٿ��?��@s[Hr��3@��]^�!?�O��@�Ar�>�ٿ��?��@s[Hr��3@��]^�!?�O��@�!�)�ٿ��F�A�@]͹A>�3@��|�!?��3�D�@�!�)�ٿ��F�A�@]͹A>�3@��|�!?��3�D�@�!�)�ٿ��F�A�@]͹A>�3@��|�!?��3�D�@��E�ٿ��ѓ��@�����3@�h<w��!?|5P����@��E�ٿ��ѓ��@�����3@�h<w��!?|5P����@��E�ٿ��ѓ��@�����3@�h<w��!?|5P����@��E�ٿ��ѓ��@�����3@�h<w��!?|5P����@�K �7�ٿW��.g�@Y*�2�3@_�Vפ�!?i�-��@�K �7�ٿW��.g�@Y*�2�3@_�Vפ�!?i�-��@���s��ٿ��2:��@8����3@�Q����!?�E%[���@���s��ٿ��2:��@8����3@�Q����!?�E%[���@���s��ٿ��2:��@8����3@�Q����!?�E%[���@�UcK�ٿ�αz��@x�l�.�3@�z�G��!?d�M����@��~��ٿ7�E�@�@��_�3@w�['�!?ě4X�
�@�@]�ٿ9x����@8M-���3@��>s��!?W�w�G��@�@]�ٿ9x����@8M-���3@��>s��!?W�w�G��@ī���ٿ`c�g9<�@#\5@~�3@�����!?��H(�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@>�mťٿ�l����@�����3@�����!?C\�?�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@o�R���ٿZ&ZʌC�@&���3@�L�H��!?m��1�`�@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��g�_�ٿ�����@����3@��=Z�!?�~����@��A��ٿL̾N5��@$|]�^�3@)���!?I*�L��@"f�+B�ٿ�#`��9�@JG����3@W�F�А!?��0J��@"f�+B�ٿ�#`��9�@JG����3@W�F�А!?��0J��@"f�+B�ٿ�#`��9�@JG����3@W�F�А!?��0J��@F���ٿ�8�v�@��ݫ�3@�t����!?s'r��{�@��2-�ٿg�:B�6�@@ɕ�R�3@#�`���!?uBDZU�@��g���ٿ�k�9�@\�3�N�3@�dd�א!?1N�7�2�@��g���ٿ�k�9�@\�3�N�3@�dd�א!?1N�7�2�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@b�kTy�ٿ��H�*�@�\���3@��k���!?�Z^�":�@�	䜢ٿk�����@lT�F��3@*�2��!?�Z�`���@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@Z���*�ٿ�x3�O`�@2ӄ��3@܅+���!?�@K����@ۣ�a8�ٿ�����R�@�ɤN��3@iEn��!?lc�/���@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@��銞�ٿ���S�@� H���3@��|���!?-�m>l�@���0-�ٿbΫ����@)Q����3@��А!?
r�$ʩ�@�u����ٿ-:}�}�@�*�`��3@�qRܐ!?+�J`]�@�u����ٿ-:}�}�@�*�`��3@�qRܐ!?+�J`]�@�u����ٿ-:}�}�@�*�`��3@�qRܐ!?+�J`]�@�u����ٿ-:}�}�@�*�`��3@�qRܐ!?+�J`]�@~Jj��ٿ7he+��@F�B:�3@&#`�А!?'�]�F�@~Jj��ٿ7he+��@F�B:�3@&#`�А!?'�]�F�@a)��͡ٿ/9/� �@.$����3@�j
��!?itrkא�@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��t�:�ٿ��g��@��;���3@m���ǐ!?� �zG��@��Ff�ٿJ.�\3m�@�"�Q�3@m_ƶ�!?���SR�@��Ff�ٿJ.�\3m�@�"�Q�3@m_ƶ�!?���SR�@��'�ٿ������@�o��3@~�2�y�!?�Z�����@��'�ٿ������@�o��3@~�2�y�!?�Z�����@��'�ٿ������@�o��3@~�2�y�!?�Z�����@��'�ٿ������@�o��3@~�2�y�!?�Z�����@��'�ٿ������@�o��3@~�2�y�!?�Z�����@��!(:�ٿ\��{� �@�kE�s�3@�˖���!?o_ ���@�S�.�ٿ#ұc�@ ���3@m�wlѐ!?wG���T�@�S�.�ٿ#ұc�@ ���3@m�wlѐ!?wG���T�@�S�.�ٿ#ұc�@ ���3@m�wlѐ!?wG���T�@�S�.�ٿ#ұc�@ ���3@m�wlѐ!?wG���T�@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@)�S��ٿ@�ؑ�_�@yv$x�3@Z��Dא!?:����@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@������ٿ��H4=��@���Q��3@pnL��!?*������@��?ϟٿ%) �x��@zmB7��3@L*P�͐!?h1��f�@��?ϟٿ%) �x��@zmB7��3@L*P�͐!?h1��f�@��?ϟٿ%) �x��@zmB7��3@L*P�͐!?h1��f�@��?ϟٿ%) �x��@zmB7��3@L*P�͐!?h1��f�@��3u�ٿ��ܑR~�@�x�h�3@�G���!?���.�@��x��ٿn�eJ��@
�gn��3@��!W��!?��`��@��x��ٿn�eJ��@
�gn��3@��!W��!?��`��@�A�םٿ�a���@I�Uh�3@��X\�!?�P����@�A�םٿ�a���@I�Uh�3@��X\�!?�P����@O���ٿ���~�Y�@%Cܔ!�3@�\^i�!?�[�Y���@4���¥ٿ)D�7z�@g9b��3@�5�D�!?mҸ�6�@4���¥ٿ)D�7z�@g9b��3@�5�D�!?mҸ�6�@����ٿW���e�@�����3@Щ_���!?rw]���@����ٿW���e�@�����3@Щ_���!?rw]���@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@0Zv�ٿ�5��Z�@FSwM�3@�WI��!?���ˮ�@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@p|o8O�ٿ����W�@��1�T�3@\׻]��!?�/�]��@�I!<�ٿ{!"�b�@�����3@H���ِ!?����ۣ�@�آ�4�ٿX-�h�@�=Jd
�3@
q�vƐ!?�7y	��@�آ�4�ٿX-�h�@�=Jd
�3@
q�vƐ!?�7y	��@�آ�4�ٿX-�h�@�=Jd
�3@
q�vƐ!?�7y	��@ގ��d�ٿ�[	��@	����3@S<�4��!?�2�O��@ގ��d�ٿ�[	��@	����3@S<�4��!?�2�O��@ގ��d�ٿ�[	��@	����3@S<�4��!?�2�O��@ގ��d�ٿ�[	��@	����3@S<�4��!?�2�O��@{�b���ٿ��n���@0�n��3@gh涝�!?����Z�@{�b���ٿ��n���@0�n��3@gh涝�!?����Z�@{�b���ٿ��n���@0�n��3@gh涝�!?����Z�@{�b���ٿ��n���@0�n��3@gh涝�!?����Z�@{�b���ٿ��n���@0�n��3@gh涝�!?����Z�@ڥ��P�ٿ�7�k�@�Y��l�3@|[����!?/���N�@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@3�EQ��ٿʕ���@7�ճ�3@����!?�M�F���@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@�6���ٿ;�"	K��@�Kҧ�3@R�桐!?���[�@l�[ 9�ٿf��()��@������3@�n5@ؐ!?�-zI�M�@��\��ٿT�_��@�[�1�4@M���!?J� ;v�@���8��ٿ�>w_�^�@�T�8��3@���!?�����@���8��ٿ�>w_�^�@�T�8��3@���!?�����@���8��ٿ�>w_�^�@�T�8��3@���!?�����@~�a~0�ٿ/5#{��@NQ�5�3@=&'sӐ!?B@��{X�@īXx!�ٿ��� �@Ǟ�6��3@~�;�!?��ե���@īXx!�ٿ��� �@Ǟ�6��3@~�;�!?��ե���@īXx!�ٿ��� �@Ǟ�6��3@~�;�!?��ե���@e���Сٿ���+�@e�((��3@@����!?����]�@e���Сٿ���+�@e�((��3@@����!?����]�@e���Сٿ���+�@e�((��3@@����!?����]�@e���Сٿ���+�@e�((��3@@����!?����]�@e���Сٿ���+�@e�((��3@@����!?����]�@e���Сٿ���+�@e�((��3@@����!?����]�@�����ٿ�Ҙ	=�@������3@�Bِ!?��6-"��@�����ٿ�Ҙ	=�@������3@�Bِ!?��6-"��@�k�Y4�ٿ��vy���@D�tk�3@/��ǐ!?����@�k�Y4�ٿ��vy���@D�tk�3@/��ǐ!?����@�k�Y4�ٿ��vy���@D�tk�3@/��ǐ!?����@�k�Y4�ٿ��vy���@D�tk�3@/��ǐ!?����@<����ٿO�qTɫ�@̧8�3@N�u�R�!?�KB�{�@����Q�ٿ��w�U��@���m�3@��R�L�!?)�/��@����Q�ٿ��w�U��@���m�3@��R�L�!?)�/��@����Q�ٿ��w�U��@���m�3@��R�L�!?)�/��@�f��1�ٿ������@q�+�t�3@�L^�^�!?:���@�f��1�ٿ������@q�+�t�3@�L^�^�!?:���@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@U���ٿ���1\�@U
�+�3@w�Q᷐!?3*	��@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@���g�ٿ�!9���@�d���3@)��?��!?��I�@]ς�֙ٿc���m�@O�Lf�3@�fR$��!?Y�ǥ�6�@]ς�֙ٿc���m�@O�Lf�3@�fR$��!?Y�ǥ�6�@]ς�֙ٿc���m�@O�Lf�3@�fR$��!?Y�ǥ�6�@�⺤!�ٿ?rL4���@ �V�Q�3@�b��!�!?�5���@�⺤!�ٿ?rL4���@ �V�Q�3@�b��!�!?�5���@�⺤!�ٿ?rL4���@ �V�Q�3@�b��!�!?�5���@�⺤!�ٿ?rL4���@ �V�Q�3@�b��!�!?�5���@�⺤!�ٿ?rL4���@ �V�Q�3@�b��!�!?�5���@Ԍu��ٿ�܋͊9�@�|T��3@;ͫ	�!?�t9V�@��o��ٿ0�k@��@��>p�3@k.`���!?N��fI��@��o��ٿ0�k@��@��>p�3@k.`���!?N��fI��@��o��ٿ0�k@��@��>p�3@k.`���!?N��fI��@��o��ٿ0�k@��@��>p�3@k.`���!?N��fI��@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@:Nl��ٿ�`\k��@~��\Y�3@N����!?.'�޻�@�v
.&�ٿ1I�Ý�@���"��3@-(�3ސ!?�Z�����@�v
.&�ٿ1I�Ý�@���"��3@-(�3ސ!?�Z�����@�v
.&�ٿ1I�Ý�@���"��3@-(�3ސ!?�Z�����@�v
.&�ٿ1I�Ý�@���"��3@-(�3ސ!?�Z�����@�v
.&�ٿ1I�Ý�@���"��3@-(�3ސ!?�Z�����@?� �A�ٿ�����@g(H���3@���.�!?��I\M��@?� �A�ٿ�����@g(H���3@���.�!?��I\M��@?� �A�ٿ�����@g(H���3@���.�!?��I\M��@?� �A�ٿ�����@g(H���3@���.�!?��I\M��@ܬY���ٿ�Tk���@��� w�3@�W�5:�!?#�mIX}�@ܬY���ٿ�Tk���@��� w�3@�W�5:�!?#�mIX}�@4����ٿ�.*_�@d�C���3@��o�5�!?�����@4����ٿ�.*_�@d�C���3@��o�5�!?�����@4����ٿ�.*_�@d�C���3@��o�5�!?�����@4����ٿ�.*_�@d�C���3@��o�5�!?�����@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@nNKi�ٿ����SJ�@9�p��3@�H��J�!?�m+�E��@{"���ٿh�jM*�@x�S���3@�&;�!?~$�YӍ�@{"���ٿh�jM*�@x�S���3@�&;�!?~$�YӍ�@{"���ٿh�jM*�@x�S���3@�&;�!?~$�YӍ�@{"���ٿh�jM*�@x�S���3@�&;�!?~$�YӍ�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@k�l�ٿ�[$�S�@���3@/���!?S��ү�@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@>"�Ԡٿ�N�g��@7x%d��3@IpQ,��!?U� ����@Mr�۔�ٿ�1M�!��@� ��)�3@�Du��!?ȶ�f��@Mr�۔�ٿ�1M�!��@� ��)�3@�Du��!?ȶ�f��@Mr�۔�ٿ�1M�!��@� ��)�3@�Du��!?ȶ�f��@Mr�۔�ٿ�1M�!��@� ��)�3@�Du��!?ȶ�f��@龟ٿs�Ay�@�@r�����3@Lt��k�!?�!�{@r�@龟ٿs�Ay�@�@r�����3@Lt��k�!?�!�{@r�@龟ٿs�Ay�@�@r�����3@Lt��k�!?�!�{@r�@龟ٿs�Ay�@�@r�����3@Lt��k�!?�!�{@r�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@���n�ٿ�	_����@�	ZT.�3@.�};��!?dl��-\�@�az=,�ٿ���G�@�����3@j���!?�|�Q��@�az=,�ٿ���G�@�����3@j���!?�|�Q��@�az=,�ٿ���G�@�����3@j���!?�|�Q��@��eo��ٿ�ux���@(C���3@J*��/�!?*(\�	�@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@=��Z�ٿO�L��@U��3@�6�?��!?�kM���@8���/�ٿR�����@A�HF��3@<��!?�~�!�@8���/�ٿR�����@A�HF��3@<��!?�~�!�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�f�-��ٿ�	�m�A�@���I��3@�;��!?�8ŉ�&�@�Xu��ٿ�p/U(��@a���3@+���!?�m�g�_�@�Xu��ٿ�p/U(��@a���3@+���!?�m�g�_�@�&-g5�ٿ�iCT�8�@�>o3�3@���!?�(Y���@�&-g5�ٿ�iCT�8�@�>o3�3@���!?�(Y���@D�$��ٿ��0�/V�@���2�3@��y��!?*U��g�@D�$��ٿ��0�/V�@���2�3@��y��!?*U��g�@D�$��ٿ��0�/V�@���2�3@��y��!?*U��g�@D�$��ٿ��0�/V�@���2�3@��y��!?*U��g�@�$�-��ٿ IHC��@�Y���3@)��̴�!?�|(���@��U�ٿ��l3�@oٞ�3@��Ǝ��!?�u��w�@��U�ٿ��l3�@oٞ�3@��Ǝ��!?�u��w�@��U�ٿ��l3�@oٞ�3@��Ǝ��!?�u��w�@��U�ٿ��l3�@oٞ�3@��Ǝ��!?�u��w�@�)�s�ٿ{���ae�@�U��3@9��;r�!?;���>��@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@W�����ٿh��>Q�@��z�3@��WJn�!?���x �@��w�L�ٿa��F�@^����3@��v��!?�8+G�@��w�L�ٿa��F�@^����3@��v��!?�8+G�@��b�
�ٿ���X�@X޵�3@y!	6��!?��kF��@��b�
�ٿ���X�@X޵�3@y!	6��!?��kF��@��b�
�ٿ���X�@X޵�3@y!	6��!?��kF��@��b�
�ٿ���X�@X޵�3@y!	6��!?��kF��@��b�
�ٿ���X�@X޵�3@y!	6��!?��kF��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@Bf.l�ٿ���B��@�}��i�3@�"���!?r9�Y��@9s�Dq�ٿw��d��@��s��3@�zci��!?��"���@9s�Dq�ٿw��d��@��s��3@�zci��!?��"���@���}��ٿ����߽�@�Ӎ��3@�E���!?������@���}��ٿ����߽�@�Ӎ��3@�E���!?������@u��զٿN�M��R�@��7q��3@ʛdƐ!?���q�-�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@G��ٿ�T��Ϻ�@��b�3@L��<��!?���[�!�@��P#��ٿ���nC�@{XA���3@�Tԏ�!?t���
��@��P#��ٿ���nC�@{XA���3@�Tԏ�!?t���
��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@/��y��ٿ�g�?��@A5���3@��A��!? ��~��@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@#	���ٿ�F �"�@�0���3@T�cʐ!?�j�H7�@˖a���ٿ���:F�@P�����3@��v�!?�V��@˖a���ٿ���:F�@P�����3@��v�!?�V��@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@9�ҙ�ٿ��eK�(�@���9�3@{r�ǐ!?_I1ac�@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@QZ=���ٿ����;��@��p�=�3@+K<}��!?�o�Ɲ��@F����ٿ���O>k�@���~0�3@�~{ސ!?�;�"F��@F����ٿ���O>k�@���~0�3@�~{ސ!?�;�"F��@F����ٿ���O>k�@���~0�3@�~{ސ!?�;�"F��@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@��xdT�ٿ�Gg84��@�&.=�3@nn7�!?~��];[�@�-�^�ٿ�y���@�,�K�3@��G�ؐ!?�v �N�@�-�^�ٿ�y���@�,�K�3@��G�ؐ!?�v �N�@|��py�ٿ���^�@D�
3�3@h(Ր!?EX&À��@|��py�ٿ���^�@D�
3�3@h(Ր!?EX&À��@|��py�ٿ���^�@D�
3�3@h(Ր!?EX&À��@|��py�ٿ���^�@D�
3�3@h(Ր!?EX&À��@|��py�ٿ���^�@D�
3�3@h(Ր!?EX&À��@�y-��ٿg\8�be�@�V�<N�3@�#w쬐!?Vi�oU�@�y-��ٿg\8�be�@�V�<N�3@�#w쬐!?Vi�oU�@�y-��ٿg\8�be�@�V�<N�3@�#w쬐!?Vi�oU�@�y-��ٿg\8�be�@�V�<N�3@�#w쬐!?Vi�oU�@�y-��ٿg\8�be�@�V�<N�3@�#w쬐!?Vi�oU�@)c����ٿ*���<�@�AB��3@z��iΐ!?�lA!��@)c����ٿ*���<�@�AB��3@z��iΐ!?�lA!��@)c����ٿ*���<�@�AB��3@z��iΐ!?�lA!��@�|��!�ٿ�)@�L��@����3@��Cʐ!?6_sz��@#F=^ȡٿ\Ͱ���@���,�3@P�vOא!?�����@#F=^ȡٿ\Ͱ���@���,�3@P�vOא!?�����@#F=^ȡٿ\Ͱ���@���,�3@P�vOא!?�����@#F=^ȡٿ\Ͱ���@���,�3@P�vOא!?�����@�g�ӦٿN�]"�@τ�^N�3@Q����!?]�R����@�g�ӦٿN�]"�@τ�^N�3@Q����!?]�R����@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@юڌo�ٿ~��1��@��@�e�3@�PY�!?�Ё���@�����ٿ�$�����@���,��3@���Ӑ!?;�~���@�����ٿ�$�����@���,��3@���Ӑ!?;�~���@�*_4��ٿ��Ė���@�euC�3@�=Yx�!?�r����@�*_4��ٿ��Ė���@�euC�3@�=Yx�!?�r����@�*_4��ٿ��Ė���@�euC�3@�=Yx�!?�r����@�*_4��ٿ��Ė���@�euC�3@�=Yx�!?�r����@�*_4��ٿ��Ė���@�euC�3@�=Yx�!?�r����@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@����-�ٿ5?��}�@e�g��3@��Ԑ!?"F��|	�@W�Q��ٿXZ�t�@��9�.�3@9Ad_��!?I&tx��@W�Q��ٿXZ�t�@��9�.�3@9Ad_��!?I&tx��@W�Q��ٿXZ�t�@��9�.�3@9Ad_��!?I&tx��@W�Q��ٿXZ�t�@��9�.�3@9Ad_��!?I&tx��@1~Ԓ,�ٿY��{��@�� �3@h�m���!?�<QX�k�@1~Ԓ,�ٿY��{��@�� �3@h�m���!?�<QX�k�@1~Ԓ,�ٿY��{��@�� �3@h�m���!?�<QX�k�@1~Ԓ,�ٿY��{��@�� �3@h�m���!?�<QX�k�@�Bk��ٿV�����@&�X-�3@z���ː!?'��'��@�Bk��ٿV�����@&�X-�3@z���ː!?'��'��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�Q��ٿ��b���@�.*�g�3@�(�i��!?����6��@�N��ٞٿm-���@�!���3@�����!?�mf�v��@r��O�ٿ��s���@�!���3@/��!?#5�M&k�@r��O�ٿ��s���@�!���3@/��!?#5�M&k�@�*�W|�ٿ��c|���@z-Ņ�3@Vǯ��!?�X���h�@$��ٿM�տ%�@^�;b��3@���V��!?�2�{��@$��ٿM�տ%�@^�;b��3@���V��!?�2�{��@$��ٿM�տ%�@^�;b��3@���V��!?�2�{��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@뻼"h�ٿ�˴���@�ւ�3@"�x6�!?)�3N��@?2m\Ǘٿ�n;����@���o�3@�ػ���!?�b���@?2m\Ǘٿ�n;����@���o�3@�ػ���!?�b���@?2m\Ǘٿ�n;����@���o�3@�ػ���!?�b���@!�u�Иٿ��i����@�l��3@����!?17�T��@!�u�Иٿ��i����@�l��3@����!?17�T��@!�u�Иٿ��i����@�l��3@����!?17�T��@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@o=�6�ٿ_�ܺ�i�@�5R�&�3@��.�e�!?�J���@:���ڤٿ��e�v��@��k�3@0�Fؐ!?^�F�)�@:���ڤٿ��e�v��@��k�3@0�Fؐ!?^�F�)�@:���ڤٿ��e�v��@��k�3@0�Fؐ!?^�F�)�@:���ڤٿ��e�v��@��k�3@0�Fؐ!?^�F�)�@��]�ٿ��A'z��@��Ȼ�3@Z�褏�!?]�TX��@�{q$�ٿ��p�P�@�����3@q���8�!?-�g �@�����ٿnv���@Q0����3@>
X��!?��rs�@�����ٿnv���@Q0����3@>
X��!?��rs�@>r���ٿ,e�#�k�@�Z��3@x���!?W�W0�P�@�����ٿ���v�@@�>�g�3@��m���!?�V$n���@�����ٿ���v�@@�>�g�3@��m���!?�V$n���@�����ٿ���v�@@�>�g�3@��m���!?�V$n���@��.��ٿ��MKZ�@@z���3@:�\��!?��'�@\��Z�ٿ�����,�@�[p�3@��6�!?a��B��@\��Z�ٿ�����,�@�[p�3@��6�!?a��B��@\��Z�ٿ�����,�@�[p�3@��6�!?a��B��@��B*�ٿ�`s(m�@�H}Ej�3@�;���!?qnx�,�@��B*�ٿ�`s(m�@�H}Ej�3@�;���!?qnx�,�@��B*�ٿ�`s(m�@�H}Ej�3@�;���!?qnx�,�@��B*�ٿ�`s(m�@�H}Ej�3@�;���!?qnx�,�@��B*�ٿ�`s(m�@�H}Ej�3@�;���!?qnx�,�@]Yb`'�ٿ���On�@{�C�3@�R�	�!?��@]Yb`'�ٿ���On�@{�C�3@�R�	�!?��@]Yb`'�ٿ���On�@{�C�3@�R�	�!?��@]Yb`'�ٿ���On�@{�C�3@�R�	�!?��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@ ��4'�ٿ�-�	���@A�0��3@�3*��!?�r˾Q��@oeQŠٿ5�K�!y�@�O�7�3@�6�4֐!??�d��V�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@t��ٿ mb�r�@!p|D��3@lr9�!?����ߪ�@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@���ٿ�Pz�{��@�lDC��3@�Mw<�!?�1�#s��@kk�r��ٿ�J�j�@!���3@ilA}��!?=�m-Y��@kk�r��ٿ�J�j�@!���3@ilA}��!?=�m-Y��@.n�u'�ٿdek���@?fP��3@:Gڸ��!?�j����@.n�u'�ٿdek���@?fP��3@:Gڸ��!?�j����@.n�u'�ٿdek���@?fP��3@:Gڸ��!?�j����@.n�u'�ٿdek���@?fP��3@:Gڸ��!?�j����@�R���ٿ)oe����@,��-�3@Uy��!?��@�Y�@�R���ٿ)oe����@,��-�3@Uy��!?��@�Y�@�R���ٿ)oe����@,��-�3@Uy��!?��@�Y�@
���ٿ�~	�%�@�h��3@�P����!?'�"G�%�@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@=in��ٿ�g8�#�@�C����3@R;�-ΐ!?�t�b��@u^�T�ٿ��!\G�@�f�c��3@(�qM��!?�o�l$�@u^�T�ٿ��!\G�@�f�c��3@(�qM��!?�o�l$�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@��:�a�ٿ�2%���@�]i^�3@�m]�!?�Z{�Ѥ�@vvd��ٿ݉f�h��@���d��3@�ĿEc�!?�/����@vvd��ٿ݉f�h��@���d��3@�ĿEc�!?�/����@vvd��ٿ݉f�h��@���d��3@�ĿEc�!?�/����@vvd��ٿ݉f�h��@���d��3@�ĿEc�!?�/����@�����ٿ��@:��@������3@&�3d�!?��`�"�@�����ٿ��@:��@������3@&�3d�!?��`�"�@�����ٿ��@:��@������3@&�3d�!?��`�"�@�����ٿ��@:��@������3@&�3d�!?��`�"�@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@ƙ@u�ٿ,�~p���@��V��3@a�X��!?'�꣨��@H5�	<�ٿ�5ʩ\5�@_��2�3@$&����!?g���U�@�5O�ٿ��A'o�@� ���3@x�Pä�!?(���=�@BR��M�ٿYd �j�@��o��3@聶~��!?SvM���@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@o]5M�ٿ�-�&�@0���	�3@{_,��!?�/����@�:@D��ٿwWi��d�@��j!�3@M���V�!?E��g�"�@�:@D��ٿwWi��d�@��j!�3@M���V�!?E��g�"�@�:@D��ٿwWi��d�@��j!�3@M���V�!?E��g�"�@��\���ٿ@�?L��@R�
���3@�A%!?@5��@��\���ٿ@�?L��@R�
���3@�A%!?@5��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@˒�mn�ٿ$k�b��@
q��7�3@�����!?Zd��@_D��|�ٿ4{܀l��@��D\��3@;�yǐ!?;�*��@_D��|�ٿ4{܀l��@��D\��3@;�yǐ!?;�*��@_D��|�ٿ4{܀l��@��D\��3@;�yǐ!?;�*��@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@��R<w�ٿ���H�@���ԙ�3@2% �!?�<�$���@���| �ٿ:�(��@�2��3@��/��!?IPI�>��@��[��ٿmKI�}�@���Fp�3@71I���!?������@26G�`�ٿ��SYu��@�qX��3@���)_�!?WU���@�)��ٿ!�X��I�@0:�#�3@ ��^�!?�9�R,��@�)��ٿ!�X��I�@0:�#�3@ ��^�!?�9�R,��@