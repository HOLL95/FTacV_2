�NUMPY v {'descr': '<f8', 'fortran_order': False, 'shape': (3, 10000, 5), }                                                   
������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@"�V�ٿ�������@=�( 4@��JJ[�!?�xϩ4A�@�Vvb�ٿRe�����@�W� 4@-=wtH�!?�Xý4A�@Te�|d�ٿT ��@�'�a 4@��+$<�!?	�v�4A�@Te�|d�ٿT ��@�'�a 4@��+$<�!?	�v�4A�@Te�|d�ٿT ��@�'�a 4@��+$<�!?	�v�4A�@�.#��ٿ�.m ��@�IW� 4@���=�!?�
4y4A�@�.#��ٿ�.m ��@�IW� 4@���=�!?�
4y4A�@��`y�ٿ�˖ ��@��h� 4@ )�!?��
�4A�@�9S�q�ٿ�H� ��@e14 4@:8ѐ!?�FO�4A�@H��gb�ٿ�Gl ��@= �  4@ra>�!?1�n{4A�@H��gb�ٿ�Gl ��@= �  4@ra>�!?1�n{4A�@��b�ٿ�U ��@�`Z� 4@����!?�Y��4A�@��b�ٿ�U ��@�`Z� 4@����!?�Y��4A�@Řx\�ٿbB� ��@B�a 4@�Zm�!?�<4A�@Řx\�ٿbB� ��@B�a 4@�Zm�!?�<4A�@Řx\�ٿbB� ��@B�a 4@�Zm�!?�<4A�@Řx\�ٿbB� ��@B�a 4@�Zm�!?�<4A�@3+��X�ٿ�� ��@�7�� 4@	g��!?!,m�4A�@����N�ٿn�� ��@���� 4@*�����!?e�՘4A�@����N�ٿn�� ��@���� 4@*�����!?e�՘4A�@����N�ٿn�� ��@���� 4@*�����!?e�՘4A�@6?|.e�ٿ�j] ��@�dv� 4@�i�5>�!?=�N�4A�@6?|.e�ٿ�j] ��@�dv� 4@�i�5>�!?=�N�4A�@6?|.e�ٿ�j] ��@�dv� 4@�i�5>�!?=�N�4A�@6?|.e�ٿ�j] ��@�dv� 4@�i�5>�!?=�N�4A�@6?|.e�ٿ�j] ��@�dv� 4@�i�5>�!?=�N�4A�@c�	�g�ٿ�� ��@it� 4@���=8�!?𼜢4A�@c�	�g�ٿ�� ��@it� 4@���=8�!?𼜢4A�@�R��i�ٿ�� ��@f0� 4@�$���!?�k�4A�@�R��i�ٿ�� ��@f0� 4@�$���!?�k�4A�@�p�n�ٿNLA ��@d?�� 4@�J����!?��̶4A�@�p�n�ٿNLA ��@d?�� 4@�J����!?��̶4A�@�p�n�ٿNLA ��@d?�� 4@�J����!?��̶4A�@yB$�d�ٿ�� ��@
T؜ 4@fiUL��!?��#�4A�@yB$�d�ٿ�� ��@
T؜ 4@fiUL��!?��#�4A�@g���e�ٿa5` ��@��� 4@g�'Dя!?Kj�4A�@g���e�ٿa5` ��@��� 4@g�'Dя!?Kj�4A�@g���e�ٿa5` ��@��� 4@g�'Dя!?Kj�4A�@����k�ٿ5Z� ��@9�^/ 4@�|z�j�!?yq�4A�@�le�ٿ��z ��@礸 4@i�1�!?�3�4A�@����g�ٿ�	�# ��@�䕴 4@V�����!?d�4A�@����g�ٿ�	�# ��@�䕴 4@V�����!?d�4A�@a,�zi�ٿ��B ��@5"�4 4@�;".�!?;<j�4A�@a,�zi�ٿ��B ��@5"�4 4@�;".�!?;<j�4A�@��.�v�ٿ�� ��@;[
  4@��^`y�!?�S��4A�@��.�v�ٿ�� ��@;[
  4@��^`y�!?�S��4A�@��.�v�ٿ�� ��@;[
  4@��^`y�!?�S��4A�@��.�v�ٿ�� ��@;[
  4@��^`y�!?�S��4A�@��.�v�ٿ�� ��@;[
  4@��^`y�!?�S��4A�@����{�ٿ�� ��@)�_� 4@M~ߖx�!?s�Ӿ4A�@����{�ٿ�E*$ ��@���� 4@����!?��"�4A�@�w$�~�ٿ�! ��@K���  4@�<!d�!?��(�4A�@�w$�~�ٿ�! ��@K���  4@�<!d�!?��(�4A�@�w$�~�ٿ�! ��@K���  4@�<!d�!?��(�4A�@�w$�~�ٿ�! ��@K���  4@�<!d�!?��(�4A�@A�3w�ٿ3�F ��@�:G� 4@
-5�F�!?%�>�4A�@�E��o�ٿ$� ��@��V 4@��0�!?���4A�@#`��j�ٿ!n� ��@�	V� 4@�vn�f�!?��[�4A�@#`��j�ٿ!n� ��@�	V� 4@�vn�f�!?��[�4A�@#`��j�ٿ!n� ��@�	V� 4@�vn�f�!?��[�4A�@#`��j�ٿ!n� ��@�	V� 4@�vn�f�!?��[�4A�@#`��j�ٿ!n� ��@�	V� 4@�vn�f�!?��[�4A�@�!ņj�ٿzȇ ��@Z�K 4@�s��_�!?x|~�4A�@� $'j�ٿS��
 ��@'�q@ 4@G��|�!?l]d�4A�@�|<�k�ٿGֲ ��@��3G 4@��e��!?
L6�4A�@�|<�k�ٿGֲ ��@��3G 4@��e��!?
L6�4A�@�|<�k�ٿGֲ ��@��3G 4@��e��!?
L6�4A�@4>�l�ٿ�NI ��@;	�� 4@ώ�g)�!?�'��4A�@4>�l�ٿ�NI ��@;	�� 4@ώ�g)�!?�'��4A�@4>�l�ٿ�NI ��@;	�� 4@ώ�g)�!?�'��4A�@4>�l�ٿ�NI ��@;	�� 4@ώ�g)�!?�'��4A�@4>�l�ٿ�NI ��@;	�� 4@ώ�g)�!?�'��4A�@��o�n�ٿ��Z����@Eh� 4@�)L��!?Y���4A�@��o�n�ٿ��Z����@Eh� 4@�)L��!?Y���4A�@��o�n�ٿ��Z����@Eh� 4@�)L��!?Y���4A�@���uq�ٿ�B�����@P�� 4@���'��!?����4A�@3�q�ٿ�������@jA@� 4@~�%�-�!?nP�4A�@5[E�n�ٿ�Կ  ��@�C$� 4@�`��!?�^��4A�@5[E�n�ٿ�Կ  ��@�C$� 4@�`��!?�^��4A�@5[E�n�ٿ�Կ  ��@�C$� 4@�`��!?�^��4A�@�mS^l�ٿ������@��(` 4@�,Ɇ��!?��£4A�@���5m�ٿ燎����@�*Z�  4@�뒐!?�)�4A�@���5m�ٿ燎����@�*Z�  4@�뒐!?�)�4A�@�o�ٿ������@juc& 4@݆�!?�6�4A�@�o�ٿ������@juc& 4@݆�!?�6�4A�@�o�ٿ������@juc& 4@݆�!?�6�4A�@��"o�ٿ������@\�) 4@.3�.�!?QA�4A�@C+Pdl�ٿƽ�����@�/� 4@�V/�d�!?nr��4A�@y�E<l�ٿ��I����@��~ 4@�!�DX�!?%��4A�@y�E<l�ٿ��I����@��~ 4@�!�DX�!?%��4A�@�%"m�ٿ�������@+ ��  4@Bn�<�!?��4A�@|��l�ٿ�q����@����  4@� Q勐!?x�ͻ4A�@
d Br�ٿ�'$����@`g�  4@D�Lgf�!?�ű�4A�@{��t�ٿ}T����@�oo  4@4!��!?�Vղ4A�@��/�q�ٿ�������@}�z  4@����!?�ch�4A�@"|�0m�ٿaN����@{� 4@��_Fɏ!?:��4A�@"|�0m�ٿaN����@{� 4@��_Fɏ!?:��4A�@lŮm�ٿ������@�{,�  4@��&J�!?��4A�@lŮm�ٿ������@�{,�  4@��&J�!?��4A�@�9�i�ٿ{&�����@����  4@��D�)�!?i���4A�@m�(g�ٿ�&!����@pR 4@Ɠ���!?�g�4A�@ ^�g�ٿ�$�����@ul�1 4@OEq�a�!?�#�4A�@��Ͼg�ٿ�{�����@U�  4@KV=u��!?e~*�4A�@��Ͼg�ٿ�{�����@U�  4@KV=u��!?e~*�4A�@��Ͼg�ٿ�{�����@U�  4@KV=u��!?e~*�4A�@��1�d�ٿ:�E����@dA�  4@��V~k�!?�\̲4A�@��1�d�ٿ:�E����@dA�  4@��V~k�!?�\̲4A�@�Z��c�ٿy������@pߥu  4@[�D���!?�NY�4A�@�Z��c�ٿy������@pߥu  4@[�D���!?�NY�4A�@!+Kg�ٿ�$�����@�-�f  4@�����!?r�l�4A�@!+Kg�ٿ�$�����@�-�f  4@�����!?r�l�4A�@!+Kg�ٿ�$�����@�-�f  4@�����!?r�l�4A�@m�LIh�ٿy�����@*o ���3@�O���!?q�4A�@C h�ٿ��c����@�ʦ���3@ȼ4k�!?ۛ�4A�@]a��g�ٿ������@��$���3@:0�::�!?�积4A�@]a��g�ٿ������@��$���3@:0�::�!?�积4A�@]a��g�ٿ������@��$���3@:0�::�!?�积4A�@�L��i�ٿ�m����@�����3@�w�!?���4A�@�L��i�ٿ�m����@�����3@�w�!?���4A�@sy$`f�ٿ������@�1!  4@P����!?��:�4A�@�:g�ٿreD����@w
�  4@�үr%�!?e��4A�@�:g�ٿreD����@w
�  4@�үr%�!?e��4A�@�:g�ٿreD����@w
�  4@�үr%�!?e��4A�@�:g�ٿreD����@w
�  4@�үr%�!?e��4A�@��ʟk�ٿۃi����@BB  4@m�m�$�!?��ޱ4A�@�� �m�ٿ������@D8t���3@�´;�!?�Hd�4A�@�� �m�ٿ������@D8t���3@�´;�!?�Hd�4A�@6Vco�ٿO@�����@U���3@�AerJ�!?g7X�4A�@6Vco�ٿO@�����@U���3@�AerJ�!?g7X�4A�@����o�ٿ�LM����@���c  4@d�r���!?�s�4A�@r\9�m�ٿ*������@l�����3@�6�!?�>��4A�@�DU<k�ٿix~����@R b���3@���`ۏ!?=���4A�@�8��m�ٿK������@�Gt���3@3*%�ݏ!?jMg�4A�@7C{Zk�ٿ�ke����@99����3@Fҭ�!?yȑ�4A�@7C{Zk�ٿ�ke����@99����3@Fҭ�!?yȑ�4A�@�ntan�ٿ0������@��y���3@τt|��!?��&�4A�@��m�ٿl�M����@8�����3@��A��!?yZ�4A�@r
�k�ٿ�������@� ^���3@f3ǳ)�!?�ŭ4A�@r
�k�ٿ�������@� ^���3@f3ǳ)�!?�ŭ4A�@r
�k�ٿ�������@� ^���3@f3ǳ)�!?�ŭ4A�@r
�k�ٿ�������@� ^���3@f3ǳ)�!?�ŭ4A�@r
�k�ٿ�������@� ^���3@f3ǳ)�!?�ŭ4A�@֫j�ٿ/�Y����@55���3@*ĢgB�!?��4A�@��t7m�ٿ��`����@3iG��3@��!�_�!?=x��4A�@��t7m�ٿ��`����@3iG��3@��!�_�!?=x��4A�@��t7m�ٿ��`����@3iG��3@��!�_�!?=x��4A�@��l�ٿ�<�����@������3@�h<�!?�K��4A�@���$p�ٿ�^�����@��Ƕ��3@�G�.�!?ἲ4A�@��~Sp�ٿj����@J�����3@� z�u�!?�+�4A�@��~Sp�ٿj����@J�����3@� z�u�!?�+�4A�@ v:Ur�ٿg�j����@��g,��3@s�.ك�!?�u��4A�@�Fo,r�ٿF`+����@�x���3@�зF�!?�y�4A�@�Y�u�ٿ~������@��]���3@-����!?��M�4A�@���v�ٿv������@�B�@��3@���NS�!?���4A�@q:�su�ٿ�������@�	����3@��2q�!?t'��4A�@q:�su�ٿ�������@�	����3@��2q�!?t'��4A�@�pV`s�ٿp�����@�M�E��3@D6Ӽ��!?}ت4A�@�!��r�ٿ|,p����@��=��3@�)�8n�!?|�]�4A�@�]�t�ٿ�������@��\���3@��]�Y�!?�J�4A�@̢t�ٿ!K"����@�f}���3@�4s�B�!?]cӭ4A�@̢t�ٿ!K"����@�f}���3@�4s�B�!?]cӭ4A�@��As�ٿ;�W����@2�d���3@���_�!?�_�4A�@��As�ٿ;�W����@2�d���3@���_�!?�_�4A�@��x�ٿ�j����@��P��3@u�g�!?�Sͯ4A�@��x�ٿ�j����@��P��3@u�g�!?�Sͯ4A�@��Q�{�ٿϟ����@ҟS���3@E����!?
jG�4A�@��Q�{�ٿϟ����@ҟS���3@E����!?
jG�4A�@��Q�{�ٿϟ����@ҟS���3@E����!?
jG�4A�@�8�Zz�ٿV������@\ ���3@� ��!?W���4A�@�-_t�ٿ�qS����@d����3@�R�0�!?�	ޭ4A�@��0u�ٿ_D����@�5W��3@���!�!?+�(�4A�@O�&�t�ٿB�����@�<�y��3@�5��A�!?>�n�4A�@F��v�ٿ�~=����@S'���3@�v���!?�`$�4A�@K)�nu�ٿ�0-����@ʇ�  4@�h%�!?/��4A�@K)�nu�ٿ�0-����@ʇ�  4@�h%�!?/��4A�@Ղ��v�ٿq"|����@�#  4@��\��!?z%��4A�@ӾV�z�ٿ�"����@N����3@��#�!?��,�4A�@ӾV�z�ٿ�"����@N����3@��#�!?��,�4A�@���|�ٿ�»����@o+���3@�f]�!?���4A�@m�`��ٿ�L�����@d�����3@Ql3`^�!?�=�4A�@������ٿ� ����@
�����3@�$��!?rG|�4A�@������ٿ� ����@
�����3@�$��!?rG|�4A�@������ٿ� ����@
�����3@�$��!?rG|�4A�@S�r��ٿ��S����@�5t��3@��$�!?ִ�4A�@�CH�~�ٿ������@��<��3@˳(��!?���4A�@�CH�~�ٿ������@��<��3@˳(��!?���4A�@�CH�~�ٿ������@��<��3@˳(��!?���4A�@cR��z�ٿ��*����@�*z��3@��tx��!?�Qݞ4A�@��w~�ٿd������@����3@�����!?!��4A�@��K��ٿ�������@j��u��3@��Z՚�!?��}�4A�@��K��ٿ�������@j��u��3@��Z՚�!?��}�4A�@C����ٿBAl����@RG��3@,ˆ^��!?����4A�@$��y��ٿv�����@�l���3@G𑅊�!?g<��4A�@8�2#�ٿ�}�����@�-���3@z�9�s�!?|�W�4A�@�P5^�ٿ������@�*��3@�<��t�!?� a�4A�@i>7ɀ�ٿc)r����@�z8_��3@�V�3Q�!?���4A�@���2��ٿ�wG����@������3@�@��:�!? �4A�@�����ٿct�����@݀���3@���QN�!?��4A�@�ny�ٿ�(y����@�"\���3@1]�'u�!?g@�4A�@HyP���ٿ�����@��P���3@"�&ߪ�!?{�X�4A�@�_F�z�ٿ������@l㡄��3@\�ٗ��!?ci��4A�@N7Fw�ٿƘ�����@��+u��3@�^�z�!?�{C�4A�@N7Fw�ٿƘ�����@��+u��3@�^�z�!?�{C�4A�@l�x�ٿ������@4�����3@52�t�!?��i�4A�@�7_u�ٿ%�����@=��  4@��D�5�!?h�I�4A�@�]�t�ٿ������@������3@5Y	k[�!?J���4A�@�v�q�ٿ5�x����@�r���3@���S`�!?$�4A�@z�tEp�ٿ������@�5A  4@�"��!?(�ӱ4A�@��m�ٿR�����@��&�  4@g��!?��=�4A�@.'7�c�ٿgH����@&U� 4@����!?��3�4A�@��	i�ٿFOp����@W{���3@��	��!?�&��4A�@�n3�e�ٿ�{�����@"5C  4@�KUl�!?~e�4A�@]v̚g�ٿr������@:�'  4@�l�W��!?�
��4A�@]v̚g�ٿr������@:�'  4@�l�W��!?�
��4A�@{�<l�ٿt�O����@pֵ���3@4贔��!?(ݨ�4A�@R��Yv�ٿ������@ֻt��3@[���!?�M��4A�@*Vn�x�ٿk�'����@�3c���3@f�@Z��!?_��4A�@��_�z�ٿ7).����@�����3@���oǐ!?ؖ��4A�@��_�z�ٿ7).����@�����3@���oǐ!?ؖ��4A�@��_�z�ٿ7).����@�����3@���oǐ!?ؖ��4A�@��_�z�ٿ7).����@�����3@���oǐ!?ؖ��4A�@61EZy�ٿW�o����@{vm��3@�>dʐ!?vƪ4A�@!i.��ٿ�D�����@�wc^��3@�[	א!?YV^�4A�@M�)b��ٿ�������@�c��3@�n4]�!?�v��4A�@J,�+��ٿ������@�+�R��3@KZ&Q��!?�|��4A�@�iC���ٿ
�����@�xPI��3@�m{���!?�1�4A�@�����ٿ�������@�� ���3@S:w)��!?�O�4A�@�<٣��ٿ%}�����@��r��3@���&S�!?P��4A�@�<٣��ٿ%}�����@��r��3@���&S�!?P��4A�@�<٣��ٿ%}�����@��r��3@���&S�!?P��4A�@%9����ٿ�
�����@���x��3@��QV�!?�3)�4A�@�5���ٿS�����@h����3@�h(;�!?7���4A�@�����ٿmO3����@��~��3@7��Y9�!?~*�4A�@n3R(��ٿSL(����@�)T��3@�G';4�!?�S��4A�@n3R(��ٿSL(����@�)T��3@�G';4�!?�S��4A�@0k����ٿ��+����@�'q��3@�H�;&�!?B+f�4A�@�l�ͣ�ٿt����@cB����3@���uH�!?n��4A�@�O���ٿ�������@݇���3@A�{0|�!?�P�4A�@��絙ٿŴ����@y�č��3@G�1u�!?�i�4A�@�*����ٿJ�����@^���3@��uk��!?�*�4A�@^oj��ٿ'`M����@١,��3@6����!?d�,4A�@:}��әٿ�{����@�fde��3@$�b:6�!?�K�o4A�@�+Sl��ٿN������@��2���3@,b�+�!?�K�Q4A�@�
{��ٿ`�&����@	�� ��3@��P�!?B�_<4A�@��!�ٿ������@phGf��3@���!?4aWa4A�@�Ģ�ٿ_2����@N�O���3@�V��!?�LD]4A�@�Ģ�ٿ_2����@N�O���3@�V��!?�LD]4A�@�Ģ�ٿ_2����@N�O���3@�V��!?�LD]4A�@�5-ҙٿ�c�����@!�Y���3@a�<�q�!?ڤt4A�@�5-ҙٿ�c�����@!�Y���3@a�<�q�!?ڤt4A�@��2k��ٿDF�����@@^����3@C�x�k�!?�ɛ4A�@��|��ٿ��[����@��D���3@���k�!?�"��4A�@��|��ٿ��[����@��D���3@���k�!?�"��4A�@��|��ٿ��[����@��D���3@���k�!?�"��4A�@]�;Ou�ٿ)<����@��-M��3@c�Î(�!?�+��4A�@�{�V(�ٿr' ��@.u' 4@c���g�!?���4A�@�&��ٿ�' ��@7�fu 4@w��yf�!?EZ"�4A�@Ee8��ٿ"��1 ��@�z	 4@�u�dC�!?��#5A�@Ee8��ٿ"��1 ��@�z	 4@�u�dC�!?��#5A�@j��<�ٿ�X0M ��@�$w 4@�p\�o�!?A�]u5A�@�g�ٿ]�M ��@�ģ" 4@�*]iU�!?�HN�5A�@�g�ٿ]�M ��@�ģ" 4@�*]iU�!?�HN�5A�@R���ٿ��a ��@t  4@^�z��!?�bD�5A�@�����ٿ�� ��@mu�r 4@��JM�!?�.�05A�@���V<�ٿ��Z ��@Y��� 4@ �b+�!?;m�s5A�@A��J�ٿ"��	 ��@�=�� 4@��u5�!?���5A�@]r�Øٿ_\n	 ��@`)? 4@2p).m�!?�5A�@��Fm�ٿȦth ��@Ó�� 4@`�a	�!?�I�5A�@��2ʗٿ�ŅE ��@�;7@ 4@Pԗ,�!?�3e�5A�@��2ʗٿ�ŅE ��@�;7@ 4@Pԗ,�!?�3e�5A�@�|a�ٿ��$� ��@O��% 4@�z�	#�!?�z��6A�@�|a�ٿ��$� ��@O��% 4@�z�	#�!?�z��6A�@�f��Z�ٿ��X� ��@C���  4@�e
.�!?�#�6A�@����ٿA�=B ��@�LiD 4@��םw�!?���%6A�@�����ٿ)0gp ��@1�" 4@or歯�!?H]l�6A�@s�	�ٿK�4� ��@Z_��' 4@*Q�bm�!?x��7A�@��0r�ٿ��g� ��@�0lv! 4@?M�J�!?a|�6A�@�y��N�ٿx��O ��@��fE 4@�|�B�!?6KY6A�@�ҳB�ٿW�@ ��@��@� 4@z��u�!?@��6A�@1��ٿ����@��g 4@q%c�{�!?��05A�@�a��ښٿ`�&����@#��h��3@��!?�Fs�3A�@ ߜ���ٿK��h���@��p��3@���D�!?q1@83A�@a�M�ٿ��* ��@��=  4@ґ�!?2��5A�@a�M�ٿ��* ��@��=  4@ґ�!?2��5A�@<��5�ٿ�S� ��@���	 4@k���1�!?^�8s5A�@������ٿq�j. ��@I�� 4@qM9�*�!?�O��5A�@��#a(�ٿ�'Y ��@42� 4@K�_D%�!?H*6A�@Ͻ�ׄ�ٿw� ��@es'� 4@���!?�J;5A�@����ٿݐ!X ��@�O 4@�ٴE�!?bFָ5A�@ܝ��ٿ{�- ��@e; 4@��톐!?�҈�5A�@ܝ��ٿ{�- ��@e; 4@��톐!?�҈�5A�@t�o���ٿ8������@x^s� 4@5̈́�`�!?7n�5A�@�U����ٿ�H����@Pf� 4@�b��s�!?@˞5A�@�gI���ٿ0����@0��� 4@�Nl��!?k�m$5A�@�gI���ٿ0����@0��� 4@�Nl��!?k�m$5A�@��S�c�ٿ�<X���@�r���3@9M|͋�!?᭺4A�@��S�c�ٿ�<X���@�r���3@9M|͋�!?᭺4A�@��S�c�ٿ�<X���@�r���3@9M|͋�!?᭺4A�@�Ms��ٿJ��Y���@Vw���3@������!?�j�3A�@QҚٿ�` ��@K]����3@���G�!?Z+-�3A�@l{u�ǜٿs�b����@G�����3@.�ي�!?���2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�RTRڜٿ�%V}���@�9��3@�2��9�!?Av�2A�@�Fծ.�ٿ?;���@���/��3@�����!?hΓ�1A�@����ٿ]�����@U�2M��3@Y�!v�!?/ĉv/A�@����ٿ]�����@U�2M��3@Y�!v�!?/ĉv/A�@6�]��ٿ�7�����@�܌
 4@t�.e�!?&̶�5A�@b���ٿ������@xKW� 4@�S�}�!?u��g5A�@b���ٿ������@xKW� 4@�S�}�!?u��g5A�@H ��p�ٿ�5$� ��@��Y�E 4@As���!?����8A�@�kf��ٿ��^� ��@u���= 4@$=�P-�!? V8A�@�kf��ٿ��^� ��@u���= 4@$=�P-�!? V8A�@ϰ�ݫ�ٿ���6 ��@��1 4@xA�<{�!?��V6A�@'y"�ٿ35�g ��@e�R  4@����U�!?P;�6A�@'y"�ٿ35�g ��@e�R  4@����U�!?P;�6A�@� !�Ùٿ��{����@��
���3@�M4�/�!?�TM4A�@� !�Ùٿ��{����@��
���3@�M4�/�!?�TM4A�@0��� �ٿ���U ��@z�ܿ  4@���7�!?�̭6A�@0��� �ٿ���U ��@z�ܿ  4@���7�!?�̭6A�@��\)�ٿX��Q ��@NLc�- 4@���C�!?i8�7A�@��\)�ٿX��Q ��@NLc�- 4@���C�!?i8�7A�@+ՠ��ٿ0�LR ��@�pb{ 4@���=�!?�bgr6A�@����K�ٿ�m����@%�d� 4@�վ��!?퉬I5A�@j
�FŘٿ(������@j�7  4@�[�'+�!?�҇�4A�@j
�FŘٿ(������@j�7  4@�[�'+�!?�҇�4A�@j
�FŘٿ(������@j�7  4@�[�'+�!?�҇�4A�@�����ٿ�k?����@�ZX��3@5��5g�!?��o�3A�@��+�>�ٿ�\����@6�K�
 4@��|���!?�k��5A�@��+�>�ٿ�\����@6�K�
 4@��|���!?�k��5A�@��+�>�ٿ�\����@6�K�
 4@��|���!?�k��5A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@�Ms�j�ٿw� ��@�{vC 4@�-VC�!?Jd��8A�@.��G�ٿ�l����@��(���3@��)ᑐ!?0Ǯ�3A�@���L^�ٿ/+�����@C΀p��3@������!?p.2A�@x��ٿvl5w���@!�����3@/C��!?�`�X2A�@x��ٿvl5w���@!�����3@/C��!?�`�X2A�@�
�J�ٿ6�T����@Uy����3@� ���!?j��3A�@�
�J�ٿ6�T����@Uy����3@� ���!?j��3A�@�
�J�ٿ6�T����@Uy����3@� ���!?j��3A�@ؾ�M]�ٿ�k� ��@0�' 4@�����!?�t7A�@G@�V�ٿz�����@cy���3@!5i&=�!?Ŷ�3A�@G@�V�ٿz�����@cy���3@!5i&=�!?Ŷ�3A�@jדG�ٿ��R��@)Ru�1 4@7�^�N�!?�
}^7A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@�[^r��ٿ3�J����@�~_e��3@8a�c3�!?�L�4A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@}���ٿ?�W� ��@�U:� 4@V.0h�!?6��5A�@�~ O͚ٿ�������@>wy���3@-[�<�!?x*��3A�@60��̗ٿP�/! ��@|�^3 4@���a��!?�˭�5A�@60��̗ٿP�/! ��@|�^3 4@���a��!?�˭�5A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@��a��ٿ�@r���@�4��3@��ƈ4�!?���=4A�@~N��"�ٿҴJ ��@�д� 4@⮼���!?�v396A�@~N��"�ٿҴJ ��@�д� 4@⮼���!?�v396A�@~N��"�ٿҴJ ��@�д� 4@⮼���!?�v396A�@�c���ٿ��@ ��@�q�0 4@���-�!?_�I�4A�@�c���ٿ��@ ��@�q�0 4@���-�!?_�I�4A�@�c���ٿ��@ ��@�q�0 4@���-�!?_�I�4A�@�c���ٿ��@ ��@�q�0 4@���-�!?_�I�4A�@�c���ٿ��@ ��@�q�0 4@���-�!?_�I�4A�@��&��ٿ�}����@xQ���3@�>z^�!?���H4A�@��&��ٿ�}����@xQ���3@�>z^�!?���H4A�@��&��ٿ�}����@xQ���3@�>z^�!?���H4A�@pE�n��ٿ��� ��@�8" 4@/�/�w�!?AY�s6A�@pE�n��ٿ��� ��@�8" 4@/�/�w�!?AY�s6A�@�\cE��ٿj�j��@oM�F= 4@�
3K�!?����7A�@/�G$:�ٿ�ə��@�ÿ�Z 4@��Lہ�!?BA�8A�@/�G$:�ٿ�ə��@�ÿ�Z 4@��Lہ�!?BA�8A�@�dH�3�ٿ�4L���@����x 4@�c�bR�!?pJ�9A�@�dH�3�ٿ�4L���@����x 4@�c�bR�!?pJ�9A�@�dH�3�ٿ�4L���@����x 4@�c�bR�!?pJ�9A�@��o��ٿO$C ��@*�����3@��w#�!?A�#4A�@��o��ٿO$C ��@*�����3@��w#�!?A�#4A�@��o��ٿO$C ��@*�����3@��w#�!?A�#4A�@��o��ٿO$C ��@*�����3@��w#�!?A�#4A�@:Q3z�ٿ[�����@�i4���3@���W�!?Ȣ�q2A�@:Q3z�ٿ[�����@�i4���3@���W�!?Ȣ�q2A�@:Q3z�ٿ[�����@�i4���3@���W�!?Ȣ�q2A�@:Q3z�ٿ[�����@�i4���3@���W�!?Ȣ�q2A�@��BeA�ٿ8�U���@f����3@�� �!?��XT4A�@��BeA�ٿ8�U���@f����3@�� �!?��XT4A�@�:ߓu�ٿ��yP���@H>� 4@�+����!?�H�6A�@�:ߓu�ٿ��yP���@H>� 4@�+����!?�H�6A�@�Ě��ٿ�*���@�UQ 4@��P�(�!?΅�9A�@�Ě��ٿ�*���@�UQ 4@��P�(�!?΅�9A�@�����ٿ��[���@�g��< 4@��ץ��!?�w�x:A�@�է��ٿS�����@����R 4@�l��W�!?H)�<A�@ ?�/�ٿ1G@���@"�� 4@��3(�!?�Z*�8A�@ ?�/�ٿ1G@���@"�� 4@��3(�!?�Z*�8A�@ ?�/�ٿ1G@���@"�� 4@��3(�!?�Z*�8A�@ ?�/�ٿ1G@���@"�� 4@��3(�!?�Z*�8A�@ ?�/�ٿ1G@���@"�� 4@��3(�!?�Z*�8A�@l2�ߏٿ�_�����@�$�{. 4@���ߏ!?���5=A�@l2�ߏٿ�_�����@�$�{. 4@���ߏ!?���5=A�@l2�ߏٿ�_�����@�$�{. 4@���ߏ!?���5=A�@l2�ߏٿ�_�����@�$�{. 4@���ߏ!?���5=A�@��$S�ٿ�}i����@% x�& 4@��$��!?�k��=A�@��$S�ٿ�}i����@% x�& 4@��$��!?�k��=A�@��$S�ٿ�}i����@% x�& 4@��$��!?�k��=A�@��$S�ٿ�}i����@% x�& 4@��$��!?�k��=A�@�O;�c�ٿ������@�	��3@\Ǟ��!?U^��5A�@�O;�c�ٿ������@�	��3@\Ǟ��!?U^��5A�@�y�̚ٿ������@���.��3@��×ݏ!?Icn�5A�@�y�̚ٿ������@���.��3@��×ݏ!?Icn�5A�@P��k�ٿ�����@�5K8��3@KQ�P7�!?���0A�@P��k�ٿ�����@�5K8��3@KQ�P7�!?���0A�@P��k�ٿ�����@�5K8��3@KQ�P7�!?���0A�@P��k�ٿ�����@�5K8��3@KQ�P7�!?���0A�@C�>�p�ٿ�$t����@v��Hz�3@:^��!?��e3A�@C�>�p�ٿ�$t����@v��Hz�3@:^��!?��e3A�@C�>�p�ٿ�$t����@v��Hz�3@:^��!?��e3A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@�l�ٿ��Y����@w�ń��3@����*�!?1��9A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@���z�ٿ�ϥ���@+0w%��3@���1�!?	���8A�@	��qǝٿ��-��@嘵G��3@��2F�!?���Q1A�@����ٿt����@�w���3@ �A��!?��б;A�@����ٿt����@�w���3@ �A��!?��б;A�@����ٿt����@�w���3@ �A��!?��б;A�@����ٿt����@�w���3@ �A��!?��б;A�@�U�b�ٿ[RN���@�����3@�v8:ُ!?�p��7A�@2��o�ٿZ���@�>a7�3@��$��!?i�E�7A�@2��o�ٿZ���@�>a7�3@��$��!?i�E�7A�@.�bY�ٿzw����@�.��3@w����!?��g�;A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@e(z��ٿ)��V��@Y�=��3@��S�+�!?(�Q<A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@9�9&�ٿw޶���@�bdQ�3@S�m7�!?�d=�5A�@�Q��V�ٿ������@s���t�3@`��1�!?;���6A�@|W�W�ٿҊS���@�\|`�3@��_}�!?M��:A�@��צu�ٿxG'R���@Ǚ��A�3@3h���!?x�M27A�@A��(̏ٿؐjه�@�'k[��3@��x���!?y�-�BA�@\@Y�.�ٿ�%k���@%9�/��3@��o��!?���(;A�@ �Kp��ٿ\�Q����@������3@�P��!?�d�1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@��O�ٿgS�T	��@���Y 4@�K�0�!?��1A�@����ٿ̬i���@R0��3@t7�>/�!?�[�.:A�@����ٿ̬i���@R0��3@t7�>/�!?�[�.:A�@����ٿ̬i���@R0��3@t7�>/�!?�[�.:A�@�QAӔ�ٿӲ����@h9 4@�j#vS�!?���/A�@�4�9�ٿC]����@>�n�h 4@���M�!?D�.A�@�4�9�ٿC]����@>�n�h 4@���M�!?D�.A�@�4�9�ٿC]����@>�n�h 4@���M�!?D�.A�@�4�9�ٿC]����@>�n�h 4@���M�!?D�.A�@�>+3�ٿ5���@��Qo�3@:�COZ�!?�Fx=A�@�>+3�ٿ5���@��Qo�3@:�COZ�!?�Fx=A�@Ů�q��ٿ\�oz���@�鵘�3@�Á�l�!?�M��<A�@��⿓ٿ�A`(��@��S�e 4@Z~l��!?d��3A�@��⿓ٿ�A`(��@��S�e 4@Z~l��!?d��3A�@��⿓ٿ�A`(��@��S�e 4@Z~l��!?d��3A�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�(�O��ٿh��݇�@�~=��3@�h�k�!?%y~8AA�@�B$<Ǒٿ�L����@~M�# 4@�*�!?��6�:A�@�B$<Ǒٿ�L����@~M�# 4@�*�!?��6�:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@ռHꯕٿ湩���@��й�3@B�G�(�!?8��m:A�@�`��^�ٿYY����@ad����3@`���!?��<6A�@�`��^�ٿYY����@ad����3@`���!?��<6A�@�Z����ٿ��ڇ�@w^�/��3@m��&�!?���a>A�@�Z����ٿ��ڇ�@w^�/��3@m��&�!?���a>A�@'+7A�ٿB��`���@�TO�_�3@vEM�:�!?��>1A�@'+7A�ٿB��`���@�TO�_�3@vEM�:�!?��>1A�@'+7A�ٿB��`���@�TO�_�3@vEM�:�!?��>1A�@���!�ٿ�	\����@8�)L�3@ �-�/�!?�8�/A�@���!�ٿ�	\����@8�)L�3@ �-�/�!?�8�/A�@���!�ٿ�	\����@8�)L�3@ �-�/�!?�8�/A�@�Ч��ٿo����@���Ȕ 4@��~�;�!?^��N2A�@�Ч��ٿo����@���Ȕ 4@��~�;�!?^��N2A�@i��pA�ٿwM���@�."J��3@Ș8G��!?�X|8A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@��", �ٿeHM���@u��k4@>#(�!?M�.0A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@�l�m�ٿ���@��@L	!k�4@e��\�!?�W�k%A�@\v<x�ٿ�&��X��@Å؜�4@�ٍ�g�!?��IA�@\v<x�ٿ�&��X��@Å؜�4@�ٍ�g�!?��IA�@\v<x�ٿ�&��X��@Å؜�4@�ٍ�g�!?��IA�@\v<x�ٿ�&��X��@Å؜�4@�ٍ�g�!?��IA�@v�dm)�ٿG�Τ��@+���4@�$5k�!?VFlA�@ԅb��ٿ�㋩��@H�&��4@�ډ�y�!?JB�}A�@ԅb��ٿ�㋩��@H�&��4@�ډ�y�!?JB�}A�@�}��ٿҲ6����@���2�4@���ux�!?*�ϵA�@�}��ٿҲ6����@���2�4@���ux�!?*�ϵA�@�I�=�ٿ4zM�)��@G9OB�4@� ��s�!?��<�'A�@�n`:͙ٿ=��nx��@1�7��4@+��ß�!?�qjA�@�n`:͙ٿ=��nx��@1�7��4@+��ß�!?�qjA�@�n`:͙ٿ=��nx��@1�7��4@+��ß�!?�qjA�@�n`:͙ٿ=��nx��@1�7��4@+��ß�!?�qjA�@��Nfk�ٿ�����@ɘ���3@���<��!?���Q2A�@�J�-.�ٿO�����@rO(��3@Ǔh�=�!?,"��FA�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@^	�X�ٿ��/Rׇ�@ ��3:�3@6�xU�!?�b�8A�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���ٿ�o�@��@!� ��3@k�т_�!?Jj,�XA�@���^�ٿ$���@����3@�u��\�!?��wA�@���^�ٿ$���@����3@�u��\�!?��wA�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�O��ٿ/X�iz��@�:�D�3@�AM�!?E}��A�@�\����ٿ�
{>��@���Y�3@�A�[�!?E<��A�@�\����ٿ�
{>��@���Y�3@�A�[�!?E<��A�@�\����ٿ�
{>��@���Y�3@�A�[�!?E<��A�@�\����ٿ�
{>��@���Y�3@�A�[�!?E<��A�@�c�%��ٿ���&ۅ�@�Qw���3@T*>�d�!?Q]�m�A�@�c�%��ٿ���&ۅ�@�Qw���3@T*>�d�!?Q]�m�A�@�c�%��ٿ���&ۅ�@�Qw���3@T*>�d�!?Q]�m�A�@ Nat��ٿ� l��@]��+
�3@�?+��!?s�D�A�@ Nat��ٿ� l��@]��+
�3@�?+��!?s�D�A�@ Nat��ٿ� l��@]��+
�3@�?+��!?s�D�A�@�ߤ��ٿtP�^N��@��vi�4@`�!��!?Æ�pA�@�ߤ��ٿtP�^N��@��vi�4@`�!��!?Æ�pA�@�ߤ��ٿtP�^N��@��vi�4@`�!��!?Æ�pA�@�����ٿ�9����@���M��3@�Z�+��!?N�`A�@�����ٿ�9����@���M��3@�Z�+��!?N�`A�@�����ٿ�9����@���M��3@�Z�+��!?N�`A�@�����ٿ�9����@���M��3@�Z�+��!?N�`A�@�����ٿ�9����@���M��3@�Z�+��!?N�`A�@b@��7�ٿ_�EĆ�@ї����3@�kg�ʐ!?�wB^A�@b@��7�ٿ_�EĆ�@ї����3@�kg�ʐ!?�wB^A�@b@��7�ٿ_�EĆ�@ї����3@�kg�ʐ!?�wB^A�@b@��7�ٿ_�EĆ�@ї����3@�kg�ʐ!?�wB^A�@n��DC�ٿ��ڀA��@�]4���3@��q��!?;���/A�@n��DC�ٿ��ڀA��@�]4���3@��q��!?;���/A�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@^_����ٿ�@��@yx�"�3@�=; �!?Ǧ.yA�@cњٿ�W,eR��@�(����3@@&�̻�!?��|uA�@cњٿ�W,eR��@�(����3@@&�̻�!?��|uA�@̚UU�ٿ6�l���@8JiOI4@�"U=^�!?��A�@̚UU�ٿ6�l���@8JiOI4@�"U=^�!?��A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�fG�ٿ�V�p��@zh�p�3@�\��!?�&�`;A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@�d�ѓٿ��L��@5M���3@C��!1�!?��ʋ\A�@���uǖٿ�]�6X��@u��N�3@�Ƙ���!?�-��BA�@���uǖٿ�]�6X��@u��N�3@�Ƙ���!?�-��BA�@���uǖٿ�]�6X��@u��N�3@�Ƙ���!?�-��BA�@���uǖٿ�]�6X��@u��N�3@�Ƙ���!?�-��BA�@�d�Z��ٿ¦��_��@t���3@��L��!?�
te�A�@��D�ٚٿ���}}��@�P�3@@$��2�!?�鏞�A�@��D�ٚٿ���}}��@�P�3@@$��2�!?�鏞�A�@�W�J�ٿ���#��@Jc2��3@�z?�!?s�sxaA�@�W�J�ٿ���#��@Jc2��3@�z?�!?s�sxaA�@�W�J�ٿ���#��@Jc2��3@�z?�!?s�sxaA�@�W�J�ٿ���#��@Jc2��3@�z?�!?s�sxaA�@�W�J�ٿ���#��@Jc2��3@�z?�!?s�sxaA�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@3i�R4�ٿ0�Ĉ�@d�=4@��Aa?�!?3$�#
A�@.��+�ٿG.KZ���@�k���3@qŻ�!?B�xtA�@.��+�ٿG.KZ���@�k���3@qŻ�!?B�xtA�@.��+�ٿG.KZ���@�k���3@qŻ�!?B�xtA�@yr��F�ٿS�҇��@ro��e4@��)��!?Wl�l@A�@yr��F�ٿS�҇��@ro��e4@��)��!?Wl�l@A�@yr��F�ٿS�҇��@ro��e4@��)��!?Wl�l@A�@yr��F�ٿS�҇��@ro��e4@��)��!?Wl�l@A�@yr��F�ٿS�҇��@ro��e4@��)��!?Wl�l@A�@�jNg�ٿ��~��@�e��[4@ǟ���!?C�t�@�@�jNg�ٿ��~��@�e��[4@ǟ���!?C�t�@�@���=j�ٿq���@��OX4 4@Yw@�!?�2��A�@�wⰝٿ�}|���@�*���3@�GsT�!?LTO�#A�@�wⰝٿ�}|���@�*���3@�GsT�!?LTO�#A�@�wⰝٿ�}|���@�*���3@�GsT�!?LTO�#A�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@ye��ݚٿ��W����@��P�-�3@j�U��!?����AA�@e-�=śٿ��Cn��@=��$�3@�cu��!?G�PA�@Ey�xÚٿ{Wˢ��@JSP�4@)��H�!?m��A�@��ː�ٿ� �ׇ�@ R�	��3@�g#�3�!?��
�OA�@��ː�ٿ� �ׇ�@ R�	��3@�g#�3�!?��
�OA�@��ː�ٿ� �ׇ�@ R�	��3@�g#�3�!?��
�OA�@���-��ٿxU:c��@uAĭ'�3@����H�!?;4
QA�@���-��ٿxU:c��@uAĭ'�3@����H�!?;4
QA�@�[�'�ٿtN=o>��@�|Z��3@��2�!?�恞A�@�[�'�ٿtN=o>��@�|Z��3@��2�!?�恞A�@�[�'�ٿtN=o>��@�|Z��3@��2�!?�恞A�@��}H�ٿ16��W��@�(��3@q?M��!?��>��A�@��}H�ٿ16��W��@�(��3@q?M��!?��>��A�@�p����ٿ>_�`]��@�0�N�3@�-7ː!??G!2{A�@�p����ٿ>_�`]��@�0�N�3@�-7ː!??G!2{A�@�p����ٿ>_�`]��@�0�N�3@�-7ː!??G!2{A�@�p����ٿ>_�`]��@�0�N�3@�-7ː!??G!2{A�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@�Fdxr�ٿq�yV���@���9�3@��ʐ��!?u�e�uA�@m]�ٿ��z���@@��<��3@��L 8�!?bc8�A�@�
?V;�ٿ�	1W��@ۺ�T�3@L��Tv�!?�OD�_A�@�
?V;�ٿ�	1W��@ۺ�T�3@L��Tv�!?�OD�_A�@�
?V;�ٿ�	1W��@ۺ�T�3@L��Tv�!?�OD�_A�@$
{�_�ٿ����H��@��%�4@6�8�!?��A�@$
{�_�ٿ����H��@��%�4@6�8�!?��A�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@I���ʙٿ/�1���@��C�4@}XL�b�!?��dS�@�@�-�f��ٿ�k\	���@�v>��3@�yY�!?���T=A�@Z!\Ɛٿ���Cw��@���yT�3@D�FT�!?�e�ۿA�@Z!\Ɛٿ���Cw��@���yT�3@D�FT�!?�e�ۿA�@Z!\Ɛٿ���Cw��@���yT�3@D�FT�!?�e�ۿA�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@|E,��ٿҼ�����@��k��4@-�s��!?�	�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@�w�3�ٿ�8p�X��@U�w���3@8�e�M�!?���(�A�@��&�ٿ;�oiU��@�	���3@y�Y�Q�!?&X�A�@��&�ٿ;�oiU��@�	���3@y�Y�Q�!?&X�A�@��&�ٿ;�oiU��@�	���3@y�Y�Q�!?&X�A�@��&�ٿ;�oiU��@�	���3@y�Y�Q�!?&X�A�@��&�ٿ;�oiU��@�	���3@y�Y�Q�!?&X�A�@�_OMΗٿ������@M��p�3@`y}4�!?��\�kB�@�_OMΗٿ������@M��p�3@`y}4�!?��\�kB�@�_OMΗٿ������@M��p�3@`y}4�!?��\�kB�@�_OMΗٿ������@M��p�3@`y}4�!?��\�kB�@�_OMΗٿ������@M��p�3@`y}4�!?��\�kB�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@#�mk��ٿ�Pʭ��@�ܭ��3@:�����!?�~|��B�@"/��̒ٿه�]݅�@�km���3@��V�!?�A�9�B�@"/��̒ٿه�]݅�@�km���3@��V�!?�A�9�B�@"/��̒ٿه�]݅�@�km���3@��V�!?�A�9�B�@�2I1D�ٿʖw��@7�@H�
4@s����!?!��A�@�2I1D�ٿʖw��@7�@H�
4@s����!?!��A�@�2I1D�ٿʖw��@7�@H�
4@s����!?!��A�@���hӟٿ�"�����@(�^��3@B(]z׏!?F���'B�@���hӟٿ�"�����@(�^��3@B(]z׏!?F���'B�@�ӝ��ٿ�e��Ն�@(α��3@� �2ŏ!?��~�)B�@�ӝ��ٿ�e��Ն�@(α��3@� �2ŏ!?��~�)B�@�ӝ��ٿ�e��Ն�@(α��3@� �2ŏ!?��~�)B�@�ӝ��ٿ�e��Ն�@(α��3@� �2ŏ!?��~�)B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@�Xר��ٿ{3��g��@>ɑ��3@m��(�!?����>B�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@����Ǘٿ�e;�|��@�Ө �3@Z��u�!?�!DmA�@K$f�ٿ�[�J��@�K�=�3@�w[Y��!?�~>A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��K�Q�ٿn�(hl��@V����3@����!?�Gk�A�@��ҥT�ٿ`X�ۇ�@R�6�v�3@P���!?Y��?A�@^�s��ٿޔ?����@"�R��3@%$V�X�!?-�:|LA�@^�s��ٿޔ?����@"�R��3@%$V�X�!?-�:|LA�@��o��ٿI���{��@�h���3@�;�À�!? O�ULA�@��o��ٿI���{��@�h���3@�;�À�!? O�ULA�@е��ٖٿƖ$�W��@�,��3@����!?Ir�;pA�@е��ٖٿƖ$�W��@�,��3@����!?Ir�;pA�@е��ٖٿƖ$�W��@�,��3@����!?Ir�;pA�@е��ٖٿƖ$�W��@�,��3@����!?Ir�;pA�@е��ٖٿƖ$�W��@�,��3@����!?Ir�;pA�@��ܹ�ٿ�~q�H��@�AR��4@*?�rp�!?��Ӵ=A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@ѱڌ�ٿ�1ٛ\��@!vL��3@K��w�!?�;���A�@���a8�ٿyq|v̅�@:X���3@�߃�f�!?��]B�@���a8�ٿyq|v̅�@:X���3@�߃�f�!?��]B�@��F�ٿ�����@��đ��3@�9�O�!?�vJ�B�@��F�ٿ�����@��đ��3@�9�O�!?�vJ�B�@��F�ٿ�����@��đ��3@�9�O�!?�vJ�B�@��F�ٿ�����@��đ��3@�9�O�!?�vJ�B�@4�)ݑ�ٿ[�ʆ�@����3@K&�q�!?�c�8�A�@4�)ݑ�ٿ[�ʆ�@����3@K&�q�!?�c�8�A�@4�)ݑ�ٿ[�ʆ�@����3@K&�q�!?�c�8�A�@4�)ݑ�ٿ[�ʆ�@����3@K&�q�!?�c�8�A�@ �����ٿ�|�L}��@K�� 4@s��!?����A�@ �����ٿ�|�L}��@K�� 4@s��!?����A�@ �����ٿ�|�L}��@K�� 4@s��!?����A�@ل:�g�ٿë���@��&�9�3@U}k���!?�ӈ9�A�@�D���ٿ0�w"{��@ѓ�44@l���!?2�x[(A�@�U�mx�ٿ��D>��@��T�4@j*�D4�!?K
n|AC�@�U�mx�ٿ��D>��@��T�4@j*�D4�!?K
n|AC�@�U�mx�ٿ��D>��@��T�4@j*�D4�!?K
n|AC�@PZҌٿ��
��@� m�u4@����!?q���vC�@PZҌٿ��
��@� m�u4@����!?q���vC�@PZҌٿ��
��@� m�u4@����!?q���vC�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@���>&�ٿ��ѨL��@��M���3@�B!�!?DP�� C�@%ŭ}�ٿ�J����@��ܯ�	4@��t Y�!?��m�hD�@%ŭ}�ٿ�J����@��ܯ�	4@��t Y�!?��m�hD�@x��="�ٿËx����@�vNX�	4@����!?�w�ʸE�@x��="�ٿËx����@�vNX�	4@����!?�w�ʸE�@x��="�ٿËx����@�vNX�	4@����!?�w�ʸE�@x��="�ٿËx����@�vNX�	4@����!?�w�ʸE�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@������ٿM��p���@Yl�h�4@+�!�ԏ!?p��G�@h���>�ٿ�ͰD"��@Mn��3@�Z�Q��!?����C�@~yze�ٿ���=��@�i
�3@E����!?���8C�@~yze�ٿ���=��@�i
�3@E����!?���8C�@~yze�ٿ���=��@�i
�3@E����!?���8C�@� ���ٿ!)Y���@�N$�V4@1�_�,�!?W,*G�@� ���ٿ!)Y���@�N$�V4@1�_�,�!?W,*G�@� ���ٿ!)Y���@�N$�V4@1�_�,�!?W,*G�@� ���ٿ!)Y���@�N$�V4@1�_�,�!?W,*G�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@����ٿ;�E���@yE:y�4@ö���!?�Mz�"J�@�O� ȘٿC������@a%��3@<A�~�!?C�bQF�@�O� ȘٿC������@a%��3@<A�~�!?C�bQF�@y���ٿ+{�L��@�mR���3@ʅw�\�!?>����J�@~a��ٿ@�E���@�k��4@���!?�
_'H�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@t����ٿ������@�^�( �3@���c/�!?�CN��B�@����M�ٿ`�L�u��@�A;��3@� �*�!?B^R�8�@O� ��ٿ��,���@����3@�ҍ4�!?\6h�8�@O� ��ٿ��,���@����3@�ҍ4�!?\6h�8�@O� ��ٿ��,���@����3@�ҍ4�!?\6h�8�@O� ��ٿ��,���@����3@�ҍ4�!?\6h�8�@Q5�$`�ٿ��b���@��܊d�3@(�+<�!?$���IC�@Q5�$`�ٿ��b���@��܊d�3@(�+<�!?$���IC�@��1��ٿ�|	q}��@FJ�f��3@?��6�!?7!j�Z4�@��1��ٿ�|	q}��@FJ�f��3@?��6�!?7!j�Z4�@9�Ma�ٿ�K9��@+����3@m�T��!?����;�@M����ٿ�t]���@B�1��3@y�t�!?%�0ȴ<�@M����ٿ�t]���@B�1��3@y�t�!?%�0ȴ<�@M����ٿ�t]���@B�1��3@y�t�!?%�0ȴ<�@M����ٿ�t]���@B�1��3@y�t�!?%�0ȴ<�@M����ٿ�t]���@B�1��3@y�t�!?%�0ȴ<�@3o���ٿ-��T��@,�M���3@?Q��!?� �X7�@htj�ٿ��+�҇�@��b��3@t�k��!?��!TA�@htj�ٿ��+�҇�@��b��3@t�k��!?��!TA�@�"Q.�ٿ�$f���@�$0�T�3@��RR�!?h^uk@�@�"Q.�ٿ�$f���@�$0�T�3@��RR�!?h^uk@�@� ����ٿ� C�X��@�O)��4@g��&��!?9z?P�@� ����ٿ� C�X��@�O)��4@g��&��!?9z?P�@� ����ٿ� C�X��@�O)��4@g��&��!?9z?P�@� ����ٿ� C�X��@�O)��4@g��&��!?9z?P�@� ����ٿ� C�X��@�O)��4@g��&��!?9z?P�@���y�ٿ󌨷݁�@�vj���3@�W�"-�!?Ĥ�&L�@���y�ٿ󌨷݁�@�vj���3@�W�"-�!?Ĥ�&L�@���y�ٿ󌨷݁�@�vj���3@�W�"-�!?Ĥ�&L�@���y�ٿ󌨷݁�@�vj���3@�W�"-�!?Ĥ�&L�@���y�ٿ󌨷݁�@�vj���3@�W�"-�!?Ĥ�&L�@Pn�w`�ٿ�B��]��@9'��q�3@c�D�r�!?�^P�O�@Pn�w`�ٿ�B��]��@9'��q�3@c�D�r�!?�^P�O�@Pn�w`�ٿ�B��]��@9'��q�3@c�D�r�!?�^P�O�@Pn�w`�ٿ�B��]��@9'��q�3@c�D�r�!?�^P�O�@Pn�w`�ٿ�B��]��@9'��q�3@c�D�r�!?�^P�O�@�Vv�#�ٿw�J�8��@V���h�3@�ޠ�ҏ!?��x��2�@߅�俒ٿ��>)��@稖d,4@��-�!?��,�@߅�俒ٿ��>)��@稖d,4@��-�!?��,�@߅�俒ٿ��>)��@稖d,4@��-�!?��,�@߅�俒ٿ��>)��@稖d,4@��-�!?��,�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@/�J�ٿXz%�E��@�ը��3@sh�,�!?�7=�@��.��ٿx��F��@[Ri�@�3@z�:�!?7�^/��@��.��ٿx��F��@[Ri�@�3@z�:�!?7�^/��@��.��ٿx��F��@[Ri�@�3@z�:�!?7�^/��@��.��ٿx��F��@[Ri�@�3@z�:�!?7�^/��@�;�e�ٿ5$�Ԩ�@f|�Va�3@�A����!?�o����@�k�ٿ�eQ���@u26�
4@;�+�!?�;�F_�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@u9x��ٿ��i��@1(�z�3@�S�� �!?h6G0�(�@T8��ʖٿ���ܖ�@"����4@�+��l�!?hSp$�@T8��ʖٿ���ܖ�@"����4@�+��l�!?hSp$�@T8��ʖٿ���ܖ�@"����4@�+��l�!?hSp$�@T8��ʖٿ���ܖ�@"����4@�+��l�!?hSp$�@9��Ǖٿ���ˬ�@`ڇ��4@��#c�!?���~��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@�]L9��ٿI�����@\���4@�"F�!?.�z��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@蘡�i�ٿ/3����@9��C4@p�jt=�!?��3$��@ף���ٿ)�?1���@hv���4@�X�z�!?�v�ۖ��@ף���ٿ)�?1���@hv���4@�X�z�!?�v�ۖ��@ף���ٿ)�?1���@hv���4@�X�z�!?�v�ۖ��@��`�ٿ	�/���@�+td^�3@�_��!?�4�Q��@��`�ٿ	�/���@�+td^�3@�_��!?�4�Q��@��`�ٿ	�/���@�+td^�3@�_��!?�4�Q��@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@���HP�ٿa��j��@��b���3@W�1���!?1�ŭ�W�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@�jeJp�ٿAer��f�@�ۇ�r�3@�7?M��!?UO���c�@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@0��<��ٿ^(+��9�@L�9�m	4@����a�!?�uͱĵ@�R���ٿ6����@��y��3@���!?%���@�Le��ٿ��PPI�@��Q�"4@����m�!?�'ߥ馵@�Le��ٿ��PPI�@��Q�"4@����m�!?�'ߥ馵@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@?]ܴ�ٿQ�e1s��@C���4@nA`:t�!?�ѻm4+�@�/���ٿO�T,�`�@
�g�4@�'�]�!?�W��w�@�/���ٿO�T,�`�@
�g�4@�'�]�!?�W��w�@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@W�4\t�ٿċɻ@�@��NI?4@L�RR�!?��%_���@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���I�ٿ���sR�@��4��3@a5�J~�!?y�)�?��@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@���g�ٿ�~�y�@8�%�4@�Q	X�!?
ҳ��?�@g�����ٿ��z���@x9�R�4@^"��!?O"#Z�@g�����ٿ��z���@x9�R�4@^"��!?O"#Z�@���m��ٿq��X�-�@�|I�4@ʯĂ�!?�., ��@���m��ٿq��X�-�@�|I�4@ʯĂ�!?�., ��@���m��ٿq��X�-�@�|I�4@ʯĂ�!?�., ��@���m��ٿq��X�-�@�|I�4@ʯĂ�!?�., ��@�ԩ�g�ٿu�F��T�@�=���3@cL�R�!?�q�%{��@�ԩ�g�ٿu�F��T�@�=���3@cL�R�!?�q�%{��@�ԩ�g�ٿu�F��T�@�=���3@cL�R�!?�q�%{��@�ԩ�g�ٿu�F��T�@�=���3@cL�R�!?�q�%{��@U�\��ٿ�B���\�@!�k��3@u�.-��!??7��}�@U�\��ٿ�B���\�@!�k��3@u�.-��!??7��}�@U�\��ٿ�B���\�@!�k��3@u�.-��!??7��}�@U�\��ٿ�B���\�@!�k��3@u�.-��!??7��}�@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�=n�Y�ٿ�!S¾.�@̏ZQ��3@<��n�!?0���fٵ@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@�$^>��ٿr�Z�h�@zu@��3@3��T�!?�z��^�@� �֜ٿ6,�W��@�*^A5�3@͟L�G�!?>�C�@� �֜ٿ6,�W��@�*^A5�3@͟L�G�!?>�C�@� �֜ٿ6,�W��@�*^A5�3@͟L�G�!?>�C�@�Un��ٿy����@����u�3@,"k�m�!?�����@��7k=�ٿ���'54�@����3@̸󃗐!?L�OL�յ@��7k=�ٿ���'54�@����3@̸󃗐!?L�OL�յ@��7k=�ٿ���'54�@����3@̸󃗐!?L�OL�յ@��7k=�ٿ���'54�@����3@̸󃗐!?L�OL�յ@��7k=�ٿ���'54�@����3@̸󃗐!?L�OL�յ@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@CjR�7�ٿ'��M�@���d��3@_`�!?-�l��@K�;^.�ٿ��<(:_�@�����3@H��X}�!?��hn\t�@K�;^.�ٿ��<(:_�@�����3@H��X}�!?��hn\t�@G��M�ٿ4�E��@�ϟ�`�3@<8��<�!?��M^x�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@	`~��ٿ��e����@��w�3@<�4E9�!?�d��m�@�%�ːٿ��3�f1�@� ���3@,��Y�!?I
N�%޵@�%�ːٿ��3�f1�@� ���3@,��Y�!?I
N�%޵@�%�ːٿ��3�f1�@� ���3@,��Y�!?I
N�%޵@�%�ːٿ��3�f1�@� ���3@,��Y�!?I
N�%޵@�%�ːٿ��3�f1�@� ���3@,��Y�!?I
N�%޵@�X��w�ٿ�PmZ�@�tZwl�3@�fD�!�!?�c+�@�X��w�ٿ�PmZ�@�tZwl�3@�fD�!�!?�c+�@�X��w�ٿ�PmZ�@�tZwl�3@�fD�!�!?�c+�@�X��w�ٿ�PmZ�@�tZwl�3@�fD�!�!?�c+�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�鸑̘ٿ�n9?��@2Yz���3@ؔn;=�!?�����1�@�6{�ٿ04��'�@�Y���3@I�

�!?���Aߵ@�6{�ٿ04��'�@�Y���3@I�

�!?���Aߵ@��p��ٿR�=ϙ�@�1��3@` B�Y�!?�Ny/�@��p��ٿR�=ϙ�@�1��3@` B�Y�!?�Ny/�@=��r��ٿ?��r�@��y3�3@g.�0�!?Q�@>L�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@�@�A�ٿ�&2��@�#G 4@��|Ү�!?+36�@�@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@q��\�ٿ!�{�^M�@���4�3@V�����!?�I@C��@
��D��ٿ�7��E�@�c��3@�)&6z�!?M�N���@
��D��ٿ�7��E�@�c��3@�)&6z�!?M�N���@
��D��ٿ�7��E�@�c��3@�)&6z�!?M�N���@
��D��ٿ�7��E�@�c��3@�)&6z�!?M�N���@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�h�#�ٿ��� ���@`'X���3@�
�l�!?�U�;�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@�@��ٿ��쓉�@�8-�C�3@d��.��!?�'��$�@���9��ٿk#�ŕI�@�B$���3@|��v��!?� ��ů�@���9��ٿk#�ŕI�@�B$���3@|��v��!?� ��ů�@��o��ٿ����@�53 4@q�vY��!?t�|A�@��o��ٿ����@�53 4@q�vY��!?t�|A�@��o��ٿ����@�53 4@q�vY��!?t�|A�@��o��ٿ����@�53 4@q�vY��!?t�|A�@��o��ٿ����@�53 4@q�vY��!?t�|A�@��o��ٿ����@�53 4@q�vY��!?t�|A�@���ٿW�4��-�@�l��3@�!Di��!?d�!��@�HP
�ٿ��VEW�@�/��#�3@�Ġ�{�!?�F8� ��@�HP
�ٿ��VEW�@�/��#�3@�Ġ�{�!?�F8� ��@�HP
�ٿ��VEW�@�/��#�3@�Ġ�{�!?�F8� ��@�HP
�ٿ��VEW�@�/��#�3@�Ġ�{�!?�F8� ��@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�?���ٿRVK��^�@ƣ��I�3@~!2��!?�&_w�@�k��ٿCIvPo�@B@q� 4@�=�#a�!?!��˅`�@�0���ٿ5��0G�@ӽ��C4@�]4̐!?��F�w��@�0���ٿ5��0G�@ӽ��C4@�]4̐!?��F�w��@�0���ٿ5��0G�@ӽ��C4@�]4̐!?��F�w��@��p�ٿG8��@���L4@�xϐ!?���8�	�@��p�ٿG8��@���L4@�xϐ!?���8�	�@��p�ٿG8��@���L4@�xϐ!?���8�	�@8�~��ٿ������@4�d��	4@��"�t�!?ҋPU�=�@8�~��ٿ������@4�d��	4@��"�t�!?ҋPU�=�@���#�ٿ�"i���@�j�ܦ4@��M�'�!?��%o��@���#�ٿ�"i���@�j�ܦ4@��M�'�!?��%o��@���#�ٿ�"i���@�j�ܦ4@��M�'�!?��%o��@���#�ٿ�"i���@�j�ܦ4@��M�'�!?��%o��@���#�ٿ�"i���@�j�ܦ4@��M�'�!?��%o��@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�1��ۑٿ�F�n�@o�=���3@�,���!?感yVS�@�c�Յ�ٿ!����@��3�q�3@��I�!?]���(�@�c�Յ�ٿ!����@��3�q�3@��I�!?]���(�@�c�Յ�ٿ!����@��3�q�3@��I�!?]���(�@�c�Յ�ٿ!����@��3�q�3@��I�!?]���(�@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@v��愜ٿ��|����@YY��^�3@$�ƌ��!?���� �@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@�d_��ٿ}[��C�@0
��)�3@ߑ��!?�eL���@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@gh�e�ٿk�h��L�@;��+ �3@[
�T=�!?����H��@)x� %�ٿz@ zG�@�W�@��3@&�:��!?���L���@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@'��x��ٿj���*�@�"!I�4@3�
���!?�c)v��@��!ݑٿmy��@<,��3@���_�!?��8tB�@��!ݑٿmy��@<,��3@���_�!?��8tB�@��!ݑٿmy��@<,��3@���_�!?��8tB�@��!ݑٿmy��@<,��3@���_�!?��8tB�@��!ݑٿmy��@<,��3@���_�!?��8tB�@��S�җٿ����@�nBv�3@�H5�!?�T���@��S�җٿ����@�nBv�3@�H5�!?�T���@��S�җٿ����@�nBv�3@�H5�!?�T���@�1�ޑ�ٿc�]C�@�9�Q4@Y��>0�!?d�T8V�@�1�ޑ�ٿc�]C�@�9�Q4@Y��>0�!?d�T8V�@�6�2��ٿ��K�@|��i�3@����`�!?���D�@�WY,�ٿ�����+�@o�C��3@��zy`�!?�~Iل��@�WY,�ٿ�����+�@o�C��3@��zy`�!?�~Iل��@�WY,�ٿ�����+�@o�C��3@��zy`�!?�~Iل��@�WY,�ٿ�����+�@o�C��3@��zy`�!?�~Iل��@�WY,�ٿ�����+�@o�C��3@��zy`�!?�~Iل��@Վ�4r�ٿ����V�@����e4@��Vm%�!?0����@Վ�4r�ٿ����V�@����e4@��Vm%�!?0����@ ��Xƒٿ�]~�	�@c}��3@��C�!?�l*�lL�@v���K�ٿ=��Z��@6ӻ[�3@ G:�_�!?���"�@v���K�ٿ=��Z��@6ӻ[�3@ G:�_�!?���"�@.�C+��ٿ���~���@ȯ���3@VJ��!?����k��@.�C+��ٿ���~���@ȯ���3@VJ��!?����k��@.�C+��ٿ���~���@ȯ���3@VJ��!?����k��@.�C+��ٿ���~���@ȯ���3@VJ��!?����k��@4ԿC��ٿ��m��@�>e�Z�3@f�y
�!?��.W���@m�*�\�ٿ������@�����3@���\�!?-j 2�,�@m�*�\�ٿ������@�����3@���\�!?-j 2�,�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@t�uxޘٿ��k�=��@i(���3@��#y�!?��(�@��̗ٿ��h
�D�@��V��3@B�B�!?��/���@;�I�ߚٿ�h���F�@񯔶d�3@o��/�!?����@s8�C�ٿ9J��V,�@y��Š�3@N�c�!?�oM��@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@bSw^�ٿϬ �E�@�|�[E4@����u�!?�����@���px�ٿia��V�@��a��3@o��A�!?����"��@��*O�ٿ�9&�<�@9�Z��3@Q�_�?�!?�K�mQ��@��*O�ٿ�9&�<�@9�Z��3@Q�_�?�!?�K�mQ��@��*O�ٿ�9&�<�@9�Z��3@Q�_�?�!?�K�mQ��@��*O�ٿ�9&�<�@9�Z��3@Q�_�?�!?�K�mQ��@��*O�ٿ�9&�<�@9�Z��3@Q�_�?�!?�K�mQ��@�L�R�ٿ1 BRF_�@c,f4@R�TD��!?��\p��@�L�R�ٿ1 BRF_�@c,f4@R�TD��!?��\p��@�م �ٿ�;]��^�@v뼠��3@�2��(�!?��r]�@�م �ٿ�;]��^�@v뼠��3@�2��(�!?��r]�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@�[iЎ�ٿgF9;�8�@��=��3@ՙC��!?���~�@Vsr��ٿg�l-�@��dI��3@,��!?��b���@Vsr��ٿg�l-�@��dI��3@,��!?��b���@$#��ٿ2л��Z�@�SM�4@�N]7�!?�U��@���5�ٿt
�g�L�@��a��3@�&_�;�!?���@���5�ٿt
�g�L�@��a��3@�&_�;�!?���@���5�ٿt
�g�L�@��a��3@�&_�;�!?���@���5�ٿt
�g�L�@��a��3@�&_�;�!?���@���5�ٿt
�g�L�@��a��3@�&_�;�!?���@��~/��ٿ��2<�@'���3@b��2
�!?��Gk��@��~/��ٿ��2<�@'���3@b��2
�!?��Gk��@��~/��ٿ��2<�@'���3@b��2
�!?��Gk��@���ٿ��ޗn�@ry(�3@�!��!?���J?�@����a�ٿ��fQ�s�@��y!x�3@��:�`�!?橥1/��@����a�ٿ��fQ�s�@��y!x�3@��:�`�!?橥1/��@ߜ �&�ٿ$]�oܟ�@̳~z�3@T��oE�!?�����@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�Z��ٿ��r�V��@�6!�(�3@�����!?VaW~C�@�4R��ٿ�i�:�L�@6[I��3@�%E
��!?�5w+0l�@�4R��ٿ�i�:�L�@6[I��3@�%E
��!?�5w+0l�@�4R��ٿ�i�:�L�@6[I��3@�%E
��!?�5w+0l�@���n�ٿR%�HbI�@�����3@�12&�!?�P�e�:�@F�GC:�ٿ�*K����@/?B��4@��vV�!?4/�a��@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@ui.U�ٿ܄�ܗ%�@�����3@�*��g�!?3�b]�!�@��V ?�ٿ��^\�@�>/v��3@�C縶�!?O�2�r|�@��V ?�ٿ��^\�@�>/v��3@�C縶�!?O�2�r|�@��V ?�ٿ��^\�@�>/v��3@�C縶�!?O�2�r|�@:�4"�ٿۛ���@MC�d4@b�|���!?�#]{�}�@±��ٿ�>�����@B��{�3@���$�!?r�� ��@±��ٿ�>�����@B��{�3@���$�!?r�� ��@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@dQ��ҙٿ�ײk;��@ų��4@���!?Zg����@)���ٿ�;Br��@J�����3@M��	�!?�����~�@�F�<�ٿ�s�$��@��_S 4@˯j�!?ݗ�ƍ��@�F�<�ٿ�s�$��@��_S 4@˯j�!?ݗ�ƍ��@�8(*E�ٿ4��|�E�@��y� 4@\���!?�q>s��@�8(*E�ٿ4��|�E�@��y� 4@\���!?�q>s��@�8(*E�ٿ4��|�E�@��y� 4@\���!?�q>s��@�8(*E�ٿ4��|�E�@��y� 4@\���!?�q>s��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@��?˚ٿ��!�v��@������3@c�p��!?!a ߾��@����ٿ�pK��L�@�Q1v�4@%r��~�!?�%�2�@����ٿ�pK��L�@�Q1v�4@%r��~�!?�%�2�@����ٿ�pK��L�@�Q1v�4@%r��~�!?�%�2�@���j��ٿ=��`�@��SW4@���%G�!?�2Vq�@���j��ٿ=��`�@��SW4@���%G�!?�2Vq�@���j��ٿ=��`�@��SW4@���%G�!?�2Vq�@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@��y�ٿ_�sn�/�@�T@�v�3@��J?6�!?�����@U�^�ٿj�z�r3�@֧@��4@J�)0�!?��GdTҴ@U�^�ٿj�z�r3�@֧@��4@J�)0�!?��GdTҴ@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@%�F�ٿ�y���>�@�Z�h��3@_b��!?�����2�@�l��z�ٿ����n��@s�ۛ��3@�{7��!?|��[Go�@��%4�ٿ���n��@�8d���3@�����!?�^]�+@�@��%4�ٿ���n��@�8d���3@�����!?�^]�+@�@��%4�ٿ���n��@�8d���3@�����!?�^]�+@�@�r��Ǜٿ?�#i��@����4@ �M��!?d^\[��@�-���ٿDo�2�@�Tar4@�2U�8�!?��~̪��@�-���ٿDo�2�@�Tar4@�2U�8�!?��~̪��@�-���ٿDo�2�@�Tar4@�2U�8�!?��~̪��@�-���ٿDo�2�@�Tar4@�2U�8�!?��~̪��@�-���ٿDo�2�@�Tar4@�2U�8�!?��~̪��@D6X�N�ٿ�ە]?�@���4@S��4��!?LH�QW��@D6X�N�ٿ�ە]?�@���4@S��4��!?LH�QW��@D6X�N�ٿ�ە]?�@���4@S��4��!?LH�QW��@=?K���ٿt���^�@��G��3@��so'�!?�����@=?K���ٿt���^�@��G��3@��so'�!?�����@=?K���ٿt���^�@��G��3@��so'�!?�����@=?K���ٿt���^�@��G��3@��so'�!?�����@�C4M7�ٿNs|ߒ�@�%�B�3@W$�xO�!?Oէq^Ǵ@�C4M7�ٿNs|ߒ�@�%�B�3@W$�xO�!?Oէq^Ǵ@�C4M7�ٿNs|ߒ�@�%�B�3@W$�xO�!?Oէq^Ǵ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@��=d��ٿ(���H�@"ս/�3@����{�!?e�c�nѴ@�o/�ٿ�3�Y���@T�����3@���3�!?�[���ǵ@�o/�ٿ�3�Y���@T�����3@���3�!?�[���ǵ@�o/�ٿ�3�Y���@T�����3@���3�!?�[���ǵ@�o/�ٿ�3�Y���@T�����3@���3�!?�[���ǵ@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@�D�lu�ٿ�����@~Kn�Z�3@����!?� Q@C.�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@nh�ڛٿx�%#���@���v��3@1�N�+�!?���t)�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@�^�6&�ٿs�4ɴm�@�Ny��4@$g�y�!?��	�X�@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@���ᆖٿ�_���q�@n*���3@�Ɇw�!?�!���@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@�Ar8�ٿH��u�@�P��
�3@�D�9T�!?A�����@֡����ٿQ�4KI�@�����3@�4�&.�!?]ī���@֡����ٿQ�4KI�@�����3@�4�&.�!?]ī���@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@5Eg��ٿ�D+)��@�
�3@���5�!?2�n3��@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@z���ٿ}SC1��@�ҹ*��3@�d��C�!?��g@%q�@��]�J�ٿBbP���@��d
"�3@�l:�Y�!?���`#v�@��]�J�ٿBbP���@��d
"�3@�l:�Y�!?���`#v�@��]�J�ٿBbP���@��d
"�3@�l:�Y�!?���`#v�@��]�J�ٿBbP���@��d
"�3@�l:�Y�!?���`#v�@��]�J�ٿBbP���@��d
"�3@�l:�Y�!?���`#v�@6��ٿ���zq��@��Y���3@�n�
�!?�����@��M��ٿ6 �ٗ�@H���3@5��"��!?h$dj'��@'�3���ٿMx���g�@q`�3@��L���!?;1����@'�3���ٿMx���g�@q`�3@��L���!?;1����@'�3���ٿMx���g�@q`�3@��L���!?;1����@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@�`��ːٿj����s�@�E���3@_���!?Ø�	�@S�Q&g�ٿ��$1��@T�j��3@B�#��!?K����@S�Q&g�ٿ��$1��@T�j��3@B�#��!?K����@S�Q&g�ٿ��$1��@T�j��3@B�#��!?K����@S�Q&g�ٿ��$1��@T�j��3@B�#��!?K����@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@ ��{�ٿ�{���@��Mx��3@cۥ��!?��� #�@��.���ٿC�@RM��@��`=W�3@C��.�!?���d�@��.���ٿC�@RM��@��`=W�3@C��.�!?���d�@��.���ٿC�@RM��@��`=W�3@C��.�!?���d�@��.���ٿC�@RM��@��`=W�3@C��.�!?���d�@��.���ٿC�@RM��@��`=W�3@C��.�!?���d�@κ��R�ٿX�L9�@W��j��3@�$H�?�!?2��0��@κ��R�ٿX�L9�@W��j��3@�$H�?�!?2��0��@κ��R�ٿX�L9�@W��j��3@�$H�?�!?2��0��@κ��R�ٿX�L9�@W��j��3@�$H�?�!?2��0��@κ��R�ٿX�L9�@W��j��3@�$H�?�!?2��0��@:ﶴj�ٿ��<g��@yT��3@��V�Ϗ!?U2�T�3�@:ﶴj�ٿ��<g��@yT��3@��V�Ϗ!?U2�T�3�@:ﶴj�ٿ��<g��@yT��3@��V�Ϗ!?U2�T�3�@��~_q�ٿ�4�;��@:H�r��3@��mT��!? ����(�@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@�h8ц�ٿ�D�E��@d�?��3@�E9��!?�9�Y���@��#gt�ٿM�յn�@iw]@�3@�֧��!?W|xì�@?�C��ٿ�[�}n�@�+L��3@���ߏ!?ڒ #��@?�C��ٿ�[�}n�@�+L��3@���ߏ!?ڒ #��@?�C��ٿ�[�}n�@�+L��3@���ߏ!?ڒ #��@I5iy�ٿa�߲��@Ĵ����3@ܭ$�܏!?*0h�B�@I5iy�ٿa�߲��@Ĵ����3@ܭ$�܏!?*0h�B�@I5iy�ٿa�߲��@Ĵ����3@ܭ$�܏!?*0h�B�@ޗ��ٿ�ߗ%M�@���<�3@D����!?l��79�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@��Q�ٿ`9�Vu�@�zF/, 4@~E�T�!?�i��&�@�S5�E�ٿ���@��lƟ4@0<��!?qEb�@�S5�E�ٿ���@��lƟ4@0<��!?qEb�@�S5�E�ٿ���@��lƟ4@0<��!?qEb�@v�4 �ٿ�7��@A��%9�3@�/g��!?��3ʗ�@v�4 �ٿ�7��@A��%9�3@�/g��!?��3ʗ�@v�4 �ٿ�7��@A��%9�3@�/g��!?��3ʗ�@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@�0��ٿAG�n��@�j��F�3@�?���!?�E�V��@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@��V��ٿ��8]�@{!q�7�3@_�/�`�!?����ȴ@3/�^r�ٿ�	��1N�@f�jp��3@.yq���!?��,P]�@3/�^r�ٿ�	��1N�@f�jp��3@.yq���!?��,P]�@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@N����ٿ竸��e�@/�����3@sչ1|�!?��]p��@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@.����ٿ(�3Z�p�@��А��3@�N��!?e��4_�@�霎ٿ��Y
��@�DxW��3@cb8v��!?���9�@�霎ٿ��Y
��@�DxW��3@cb8v��!?���9�@�霎ٿ��Y
��@�DxW��3@cb8v��!?���9�@�霎ٿ��Y
��@�DxW��3@cb8v��!?���9�@�霎ٿ��Y
��@�DxW��3@cb8v��!?���9�@e�9E�ٿ����@�����3@�D�d�!?Ϝ;���@e�9E�ٿ����@�����3@�D�d�!?Ϝ;���@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@>�h?q�ٿʉ��@�@Z��y�3@o�Gdj�!?�~IW��@���z��ٿ���e�@ON{y�3@�
�^�!?A���+�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@�28��ٿ颞��@�����3@�kЙ��!?�?Z�F�@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@_/>4��ٿ������@2�_�3@&o��l�!?�&��@~IBa��ٿj�YIџ�@
�~�3@�Ś�h�!?�����K�@~IBa��ٿj�YIџ�@
�~�3@�Ś�h�!?�����K�@n�4��ٿ�,�:?�@'��L��3@�7D�!?�ub+�`�@n�4��ٿ�,�:?�@'��L��3@�7D�!?�ub+�`�@n�4��ٿ�,�:?�@'��L��3@�7D�!?�ub+�`�@n�4��ٿ�,�:?�@'��L��3@�7D�!?�ub+�`�@8�%Z�ٿ���mT��@�j���3@I�{�(�!?��ʙ�@8�%Z�ٿ���mT��@�j���3@I�{�(�!?��ʙ�@8�%Z�ٿ���mT��@�j���3@I�{�(�!?��ʙ�@8�%Z�ٿ���mT��@�j���3@I�{�(�!?��ʙ�@8�%Z�ٿ���mT��@�j���3@I�{�(�!?��ʙ�@ʹW�Ǖٿs8����@fx�%��3@I���*�!?PM`O�@ʹW�Ǖٿs8����@fx�%��3@I���*�!?PM`O�@ʹW�Ǖٿs8����@fx�%��3@I���*�!?PM`O�@��ʴ�ٿw^<x��@F�y$��3@S�L�!?f��3���@��ʴ�ٿw^<x��@F�y$��3@S�L�!?f��3���@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@Dϵ���ٿ��N���@� �B�3@oő"i�!?g�o��a�@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@�>&���ٿ�z��[\�@�]��3@֨15�!?��n��@��"�՘ٿ
?��?��@�c)�3@��:�!?G-ye��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@���ٿLd�s1��@ϧ�X��3@�����!?s��?��@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@��`�:�ٿ�q�|��@�-�E�3@aO�'�!?����r�@nf���ٿW�
�E�@��v���3@���{�!?�+e��A�@�M;S�ٿ{�|����@���`'�3@�㐔�!?��67t�@�M;S�ٿ{�|����@���`'�3@�㐔�!?��67t�@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@9t(DI�ٿ�dS1�@BRʣ�3@����y�!?�Iq�{ʹ@�b�ٿV�ﰜ��@��))�3@T�J�!?���O�״@�b�ٿV�ﰜ��@��))�3@T�J�!?���O�״@�b�ٿV�ﰜ��@��))�3@T�J�!?���O�״@A\�v��ٿ�尔��@�|�*�3@��9P�!?�{.N۴@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@#����ٿ��WXҷ�@"�ARr4@�x.M�!?��6"�<�@�v����ٿ�����`�@.��w-4@���L0�!?�x��/�@�v����ٿ�����`�@.��w-4@���L0�!?�x��/�@�v����ٿ�����`�@.��w-4@���L0�!?�x��/�@�	�l�ٿ�dwE�V�@I9�%c�3@ٗ�(�!?�dy��@�	�l�ٿ�dwE�V�@I9�%c�3@ٗ�(�!?�dy��@�	�l�ٿ�dwE�V�@I9�%c�3@ٗ�(�!?�dy��@�8��ٿ�<2*1��@]���3@X�]jO�!?u���`=�@�8��ٿ�<2*1��@]���3@X�]jO�!?u���`=�@�8��ٿ�<2*1��@]���3@X�]jO�!?u���`=�@�8��ٿ�<2*1��@]���3@X�]jO�!?u���`=�@�8��ٿ�<2*1��@]���3@X�]jO�!?u���`=�@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@m�[a�ٿU��9R�@�Vn�3@�!���!?Dz�<��@.}�� �ٿ��?ךz�@�{W��3@͋�m�!?D�O�n״@�:!o��ٿ��~�[�@����o�3@�f�V�!?����,�@�:!o��ٿ��~�[�@����o�3@�f�V�!?����,�@�:!o��ٿ��~�[�@����o�3@�f�V�!?����,�@�:!o��ٿ��~�[�@����o�3@�f�V�!?����,�@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@���ٿEV��t �@����3@rMW�!?�Iw
7��@����ٿ"��Ϧ��@e_N��3@�k94�!?:~f�@����ٿ"��Ϧ��@e_N��3@�k94�!?:~f�@����ٿ"��Ϧ��@e_N��3@�k94�!?:~f�@!K)H��ٿz$�%���@��Ӻa�3@<6��!?����x,�@���ٿ���(���@��Ⱥ��3@^W���!?<k���@��l�ٿ(�Nv���@n�^=��3@��@��!?���>��@��l�ٿ(�Nv���@n�^=��3@��@��!?���>��@��l�ٿ(�Nv���@n�^=��3@��@��!?���>��@��l�ٿ(�Nv���@n�^=��3@��@��!?���>��@�~{w7�ٿ�?m����@�o��3@xT��!?���k��@�~{w7�ٿ�?m����@�o��3@xT��!?���k��@C-+D�ٿS��f(�@29���3@������!?v�w��@C-+D�ٿS��f(�@29���3@������!?v�w��@C-+D�ٿS��f(�@29���3@������!?v�w��@~�Ms{�ٿ�H}�ߔ�@'uǫS�3@i�J��!?J�,���@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@����ٿļN�ū�@��6��3@�� ���!?P��X�@�E+��ٿ�(���@A�l��3@z�;o�!?�#��@�E+��ٿ�(���@A�l��3@z�;o�!?�#��@X�F���ٿ?i����@?3;��3@%����!?%Ş�_�@!j!/�ٿ���y��@gv��3@��;�z�!?q$g�@!j!/�ٿ���y��@gv��3@��;�z�!?q$g�@)�ٿ��r:���@�׺H��3@�k��4�!?�[��]�@)�ٿ��r:���@�׺H��3@�k��4�!?�[��]�@)�ٿ��r:���@�׺H��3@�k��4�!?�[��]�@E��@G�ٿ�F�oNS�@�x�� 4@����3�!?��6���@E��@G�ٿ�F�oNS�@�x�� 4@����3�!?��6���@E��@G�ٿ�F�oNS�@�x�� 4@����3�!?��6���@E��@G�ٿ�F�oNS�@�x�� 4@����3�!?��6���@�	t��ٿ��U�;��@Kz���3@д��o�!?����r��@�	t��ٿ��U�;��@Kz���3@д��o�!?����r��@�	t��ٿ��U�;��@Kz���3@д��o�!?����r��@�	t��ٿ��U�;��@Kz���3@д��o�!?����r��@�	t��ٿ��U�;��@Kz���3@д��o�!?����r��@��c�ٿ����@-6qh�3@�Јp��!?�~�mj�@��c�ٿ����@-6qh�3@�Јp��!?�~�mj�@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@w��F�ٿ����@�]�İ�3@=��;�!?�T���@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@F?p6��ٿ?(�I ��@EY�3@J�Z�!?�/��L�@���SR�ٿ�J�
|�@�H����3@��[�!?4�ˤ�δ@���SR�ٿ�J�
|�@�H����3@��[�!?4�ˤ�δ@���SR�ٿ�J�
|�@�H����3@��[�!?4�ˤ�δ@���SR�ٿ�J�
|�@�H����3@��[�!?4�ˤ�δ@5�_�ٿ)A�K �@z����3@�N��~�!?���dv�@5�_�ٿ)A�K �@z����3@�N��~�!?���dv�@Z�6�ٿ2��{���@��V�4@���TW�!?^�����@Z�6�ٿ2��{���@��V�4@���TW�!?^�����@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@� c�L�ٿ��?-�<�@lFIrv4@)}�j��!?H�w#m�@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���K��ٿ����y��@.���3@Y���_�!?�4�r��@���~X�ٿڗ�;'�@��W��3@B���G�!?��'����@���~X�ٿڗ�;'�@��W��3@B���G�!?��'����@��P6�ٿ,{qњٿ@r�KuD�3@f�����!?]/�0C��@��P6�ٿ,{qњٿ@r�KuD�3@f�����!?]/�0C��@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@޵��x�ٿw��g�+�@�eϏ�3@���Pn�!?gG�T�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@o�c�ٿ7dߌ��@���յ�3@D�w�!?�Y4]}�@��N�N�ٿ��$"�$�@��6�Z�3@�5��6�!?"YUd_�@��N�N�ٿ��$"�$�@��6�Z�3@�5��6�!?"YUd_�@��N�N�ٿ��$"�$�@��6�Z�3@�5��6�!?"YUd_�@��N�N�ٿ��$"�$�@��6�Z�3@�5��6�!?"YUd_�@�Y�\�ٿ8��u��@ث���3@��k�a�!?���~.��@|�M��ٿt���>�@�1��8�3@�5�"z�!?6Fy��@� ���ٿ��2?O��@���4@���!?%�#!�Ŵ@� ���ٿ��2?O��@���4@���!?%�#!�Ŵ@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@�k�sёٿg��$���@UG�G��3@?WǊ�!?Oq���9�@���C��ٿm��,�@�v���3@p�t�g�!?.4�6�[�@���C��ٿm��,�@�v���3@p�t�g�!?.4�6�[�@���C��ٿm��,�@�v���3@p�t�g�!?.4�6�[�@��7^��ٿ�g���@�.���3@�d��3�!?z߬1	�@��7^��ٿ�g���@�.���3@�d��3�!?z߬1	�@��7^��ٿ�g���@�.���3@�d��3�!?z߬1	�@��7^��ٿ�g���@�.���3@�d��3�!?z߬1	�@��7^��ٿ�g���@�.���3@�d��3�!?z߬1	�@�_݉�ٿPQ!�_��@����3@'N<`r�!?W��,��@�_݉�ٿPQ!�_��@����3@'N<`r�!?W��,��@�_݉�ٿPQ!�_��@����3@'N<`r�!?W��,��@�_݉�ٿPQ!�_��@����3@'N<`r�!?W��,��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�0s��ٿ��;��@��o9��3@@}f���!?�Y֝��@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@�61&��ٿk�j�Gc�@�����3@�޼N�!?�/H�0�@b���ۚٿ ���M\�@�����3@�u?�d�!?d���@b���ۚٿ ���M\�@�����3@�u?�d�!?d���@b���ۚٿ ���M\�@�����3@�u?�d�!?d���@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@������ٿ�`���@Zg@
��3@�=�;�!?��N��@���\��ٿ/ �7@"�@j�p�4@��PV�!?m�Q���@E�(yӟٿ�oq_���@��"@Q 4@�>$z�!??�����@E�(yӟٿ�oq_���@��"@Q 4@�>$z�!??�����@E�(yӟٿ�oq_���@��"@Q 4@�>$z�!??�����@���	�ٿ�H*%�|�@!�5HB
4@�Ӳ�\�!?�OD���@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@n�fc��ٿ��r�+��@㔼L��3@���B�!?{�,!��@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@[	����ٿ��@
h��@�lA�3@����U�!?��h9丵@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@���7�ٿWgU�2��@u��>S�3@���W�!?ח�c��@j"v�`�ٿ�Ɂ��@k��O�3@�vH�!?w�tu�ѵ@̡3"��ٿ"�!b�w�@�����3@�� �/�!?q��#��@̡3"��ٿ"�!b�w�@�����3@�� �/�!?q��#��@̡3"��ٿ"�!b�w�@�����3@�� �/�!?q��#��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@�T,! �ٿ��=�@�s�� 4@�j�R��!?��d&��@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@Cl�G�ٿ�H���@��ϱ��3@
��}�!?���|`w�@�c��$�ٿ��y����@�VmUQ�3@�8�
I�!?졛�V�@�c��$�ٿ��y����@�VmUQ�3@�8�
I�!?졛�V�@�c��$�ٿ��y����@�VmUQ�3@�8�
I�!?졛�V�@�c��$�ٿ��y����@�VmUQ�3@�8�
I�!?졛�V�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@�� ��ٿ ŮF��@�J��3@5m�[�!?�H>��p�@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@P��<f�ٿ&n~�(�@����L�3@Z�!?�VA�ٵ@�����ٿ�Hn�Z��@W�*y�3@׮�%�!?	�?		�@�����ٿ�Hn�Z��@W�*y�3@׮�%�!?	�?		�@�����ٿ�Hn�Z��@W�*y�3@׮�%�!?	�?		�@U���ٿi�1j
�@�2S���3@�gd,�!?���Г�@����ٿ�2��%��@��sg��3@�_�oC�!?�_�A��@����ٿ�2��%��@��sg��3@�_�oC�!?�_�A��@���>�ٿV���@�Ju���3@%J��i�!?0��Jp-�@���>�ٿV���@�Ju���3@%J��i�!?0��Jp-�@���>�ٿV���@�Ju���3@%J��i�!?0��Jp-�@���>�ٿV���@�Ju���3@%J��i�!?0��Jp-�@���>�ٿV���@�Ju���3@%J��i�!?0��Jp-�@(<�7�ٿ�G��'�@��*���3@�%���!?��1 ���@(<�7�ٿ�G��'�@��*���3@�%���!?��1 ���@(<�7�ٿ�G��'�@��*���3@�%���!?��1 ���@�����ٿ��:t"��@FJ�&�3@6��W�!?��2��+�@�����ٿ��:t"��@FJ�&�3@6��W�!?��2��+�@�����ٿ��:t"��@FJ�&�3@6��W�!?��2��+�@�����ٿ��:t"��@FJ�&�3@6��W�!?��2��+�@�&ĝ��ٿ苨d�@��#��3@�kt��!?������@�&ĝ��ٿ苨d�@��#��3@�kt��!?������@�&ĝ��ٿ苨d�@��#��3@�kt��!?������@�&ĝ��ٿ苨d�@��#��3@�kt��!?������@�&ĝ��ٿ苨d�@��#��3@�kt��!?������@�5=̗ٿIg�����@8I���3@�`V���!?{F\5��@�5=̗ٿIg�����@8I���3@�`V���!?{F\5��@��T�/�ٿ�#$���@
���3@};�]G�!?i"a�K�@��T�/�ٿ�#$���@
���3@};�]G�!?i"a�K�@��T�/�ٿ�#$���@
���3@};�]G�!?i"a�K�@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@Kꟍ�ٿ"ĩ��{�@m|.�d�3@���eP�!?��0����@�/�'�ٿx:�����@@��+��3@֖w�!?�u1E�@�/�'�ٿx:�����@@��+��3@֖w�!?�u1E�@�/�'�ٿx:�����@@��+��3@֖w�!?�u1E�@�/�'�ٿx:�����@@��+��3@֖w�!?�u1E�@�/�'�ٿx:�����@@��+��3@֖w�!?�u1E�@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@�G|p��ٿ�K�wQ��@(],K�3@�>�q�!?�1�E�ִ@^7�
�ٿv�|��@�&�8�3@��2;�!?��R.h�@#?j�H�ٿ[����@��`��3@��ɏ!?#-*��@#?j�H�ٿ[����@��`��3@��ɏ!?#-*��@�Z����ٿ���5b|�@�:���3@Z]�z�!?g���@�Z����ٿ���5b|�@�:���3@Z]�z�!?g���@�Z����ٿ���5b|�@�:���3@Z]�z�!?g���@�Z����ٿ���5b|�@�:���3@Z]�z�!?g���@�Z����ٿ���5b|�@�:���3@Z]�z�!?g���@��P�d�ٿ10((�q�@�����3@��O��!?j�״@��P�d�ٿ10((�q�@�����3@��O��!?j�״@�v����ٿ��G|v��@����3@=�*Q�!?R�L1W��@�v����ٿ��G|v��@����3@=�*Q�!?R�L1W��@�t�䯘ٿ*~�^�N�@k�e�!�3@���n�!?��'�g�@�t�䯘ٿ*~�^�N�@k�e�!�3@���n�!?��'�g�@�_�4V�ٿ�/�w@|�@��?�3@F�'wˏ!?�x��=�@�_�4V�ٿ�/�w@|�@��?�3@F�'wˏ!?�x��=�@�_�4V�ٿ�/�w@|�@��?�3@F�'wˏ!?�x��=�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@�h'���ٿP��n���@���^d�3@�~f��!?}��һ�@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@ �L�S�ٿߔ�&��@B~�3��3@�&��M�!?�	�ް��@�[�5�ٿ����h �@��c�3@?+�R�!?jkךP��@�[�5�ٿ����h �@��c�3@?+�R�!?jkךP��@�[�5�ٿ����h �@��c�3@?+�R�!?jkךP��@�[�5�ٿ����h �@��c�3@?+�R�!?jkךP��@�[�5�ٿ����h �@��c�3@?+�R�!?jkךP��@�N��ٿ���pw�@81���3@H�Q��!?λ�%j/�@�N��ٿ���pw�@81���3@H�Q��!?λ�%j/�@����ٿ��,��@������3@�jHM�!?9�,L%�@b�__ژٿ?��T��@혝�]�3@^�?#�!?�G�M�h�@b�__ژٿ?��T��@혝�]�3@^�?#�!?�G�M�h�@b�__ژٿ?��T��@혝�]�3@^�?#�!?�G�M�h�@b�__ژٿ?��T��@혝�]�3@^�?#�!?�G�M�h�@�aS㞓ٿ�xށ���@h��,�3@�礙J�!?���}�@�aS㞓ٿ�xށ���@h��,�3@�礙J�!?���}�@�aS㞓ٿ�xށ���@h��,�3@�礙J�!?���}�@�aS㞓ٿ�xށ���@h��,�3@�礙J�!?���}�@�����ٿ�A�8̛�@�{<�`�3@�w8�!?���x=��@�����ٿ�A�8̛�@�{<�`�3@�w8�!?���x=��@+��M�ٿ�P8/@�@ݭ0^��3@��`�!?C�?��@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@|�����ٿp�Hxv�@#,����3@�_W@T�!?��?���@�%�?�ٿ������@
��K��3@���n�!?f��f�0�@��Kњٿc����@ʭ�*z�3@��ͽl�!?/=�e	�@��Kњٿc����@ʭ�*z�3@��ͽl�!?/=�e	�@��Kњٿc����@ʭ�*z�3@��ͽl�!?/=�e	�@��Kњٿc����@ʭ�*z�3@��ͽl�!?/=�e	�@"ِ�Q�ٿ���T��@�	���3@�?�!?-$�tI�@"ِ�Q�ٿ���T��@�	���3@�?�!?-$�tI�@"ِ�Q�ٿ���T��@�	���3@�?�!?-$�tI�@"ِ�Q�ٿ���T��@�	���3@�?�!?-$�tI�@"ِ�Q�ٿ���T��@�	���3@�?�!?-$�tI�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@E�0���ٿ)bo,���@��p���3@�a.4�!?���l[�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@��qC�ٿ֋���@��3}��3@��}�B�!?����lB�@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�E��.�ٿ�x/u�$�@���J�3@�/�!?v=���Ӵ@�[��ٿ��y�@݁;]��3@���F�!?t���s��@�[��ٿ��y�@݁;]��3@���F�!?t���s��@�[��ٿ��y�@݁;]��3@���F�!?t���s��@,J��ٖٿt����@���7�3@=�c�!?G��o�z�@,J��ٖٿt����@���7�3@=�c�!?G��o�z�@,J��ٖٿt����@���7�3@=�c�!?G��o�z�@,J��ٖٿt����@���7�3@=�c�!?G��o�z�@,J��ٖٿt����@���7�3@=�c�!?G��o�z�@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@<�̙�ٿ�BT̬
�@&���3@���d �!?��-����@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@Ӟ�u�ٿ�Y�����@J�p�4�3@̥���!?c!�
%�@E�*>�ٿ���"�@����3@��
�!?) 9I��@E�*>�ٿ���"�@����3@��
�!?) 9I��@E�*>�ٿ���"�@����3@��
�!?) 9I��@E�*>�ٿ���"�@����3@��
�!?) 9I��@E�*>�ٿ���"�@����3@��
�!?) 9I��@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@�.��R�ٿi3?�>��@Q�|��3@�t� [�!?5����@{+��ٿgzycn)�@<f_(&�3@���)�!?���!dd�@{+��ٿgzycn)�@<f_(&�3@���)�!?���!dd�@��5�o�ٿf({�)�@lX����3@l��]�!?�����2�@��5�o�ٿf({�)�@lX����3@l��]�!?�����2�@��5�o�ٿf({�)�@lX����3@l��]�!?�����2�@��5�o�ٿf({�)�@lX����3@l��]�!?�����2�@ԗRhޘٿ����@��@��Y�4@>D�s��!?��R:�@ԗRhޘٿ����@��@��Y�4@>D�s��!?��R:�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@��-�ٿT�0Ӈ�@N��9�4@w��g�!?zڣY0�@�TԘ��ٿf|����@#�T�4@k��V�!?�B�h)�@�TԘ��ٿf|����@#�T�4@k��V�!?�B�h)�@�TԘ��ٿf|����@#�T�4@k��V�!?�B�h)�@�TԘ��ٿf|����@#�T�4@k��V�!?�B�h)�@!��BݕٿR�����@/�C;�3@-�0�!?D�E�[�@!��BݕٿR�����@/�C;�3@-�0�!?D�E�[�@���e$�ٿËv:�@~�$ױ�3@I��ri�!?Hi��,�@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@dO￝�ٿ�wQm��@;z���3@� �IG�!?lH�N���@��P��ٿ�`;���@<�g<4@ub��e�!?��?Ŵ@��P��ٿ�`;���@<�g<4@ub��e�!?��?Ŵ@��P��ٿ�`;���@<�g<4@ub��e�!?��?Ŵ@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@;�GL��ٿ��I�@�ri���3@&��F�!?��Ui �@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@s!`��ٿ�ܪ�U��@�Q �3@��V�!?���J+�@+_y)��ٿ�$�a���@ZK�5��3@��!f�!?�\G�ش@Q��.Ɠٿ�/�=�/�@�}\-�3@���X��!?��8V6�@Q��.Ɠٿ�/�=�/�@�}\-�3@���X��!?��8V6�@Q��.Ɠٿ�/�=�/�@�}\-�3@���X��!?��8V6�@Q��.Ɠٿ�/�=�/�@�}\-�3@���X��!?��8V6�@Q��.Ɠٿ�/�=�/�@�}\-�3@���X��!?��8V6�@���h�ٿ6Wp�S�@9�'���3@P��Az�!?z;��@���h�ٿ6Wp�S�@9�'���3@P��Az�!?z;��@���h�ٿ6Wp�S�@9�'���3@P��Az�!?z;��@���h�ٿ6Wp�S�@9�'���3@P��Az�!?z;��@���h�ٿ6Wp�S�@9�'���3@P��Az�!?z;��@��M�ٿzP؃���@]���3@�u׌Z�!?w�c;qݴ@��M�ٿzP؃���@]���3@�u׌Z�!?w�c;qݴ@�;�Ęٿ�h\��W�@�4����3@e2FQ�!?$�bF��@�;�Ęٿ�h\��W�@�4����3@e2FQ�!?$�bF��@�;�Ęٿ�h\��W�@�4����3@e2FQ�!?$�bF��@1=c��ٿ�.�e�@�q�M�3@[	?�!?x=�&l��@��8K�ٿ�3��@�����3@Y,�Ef�!?�8�})�@��8K�ٿ�3��@�����3@Y,�Ef�!?�8�})�@ν��#�ٿtKB����@�]14@�q�v��!?8�wϩ�@ν��#�ٿtKB����@�]14@�q�v��!?8�wϩ�@ν��#�ٿtKB����@�]14@�q�v��!?8�wϩ�@ν��#�ٿtKB����@�]14@�q�v��!?8�wϩ�@��4s�ٿF��A�@k c�4@W�/��!?�F��]��@��4s�ٿF��A�@k c�4@W�/��!?�F��]��@��4s�ٿF��A�@k c�4@W�/��!?�F��]��@��4s�ٿF��A�@k c�4@W�/��!?�F��]��@��4s�ٿF��A�@k c�4@W�/��!?�F��]��@�d"ϳ�ٿva���@�(H�� 4@0&`���!?H��=���@�d"ϳ�ٿva���@�(H�� 4@0&`���!?H��=���@�d"ϳ�ٿva���@�(H�� 4@0&`���!?H��=���@��>��ٿk9%�"�@ge�6�4@mX�U��!?��B���@��>��ٿk9%�"�@ge�6�4@mX�U��!?��B���@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@(���P�ٿ�!�(y��@2g��3@�l|B)�!?6�@��@�Nșٿ,:J��@���P�3@%L�.�!?����͏�@�Nșٿ,:J��@���P�3@%L�.�!?����͏�@���%��ٿ�Ù"a_�@�D+ ��3@�W:J2�!?::-���@���%��ٿ�Ù"a_�@�D+ ��3@�W:J2�!?::-���@���%��ٿ�Ù"a_�@�D+ ��3@�W:J2�!?::-���@���%��ٿ�Ù"a_�@�D+ ��3@�W:J2�!?::-���@t��3�ٿ��_��^�@���F�3@Ȗ�md�!?"�<l�@"�w%;�ٿ]�Ex��@��(�}�3@n��G�!?�R�\p�@"�w%;�ٿ]�Ex��@��(�}�3@n��G�!?�R�\p�@�ww61�ٿ��G���@{z�@v�3@=�p��!?ASVq�@�ww61�ٿ��G���@{z�@v�3@=�p��!?ASVq�@�ww61�ٿ��G���@{z�@v�3@=�p��!?ASVq�@>uf��ٿ���~�@��s�3@�c39�!?�bV�
�@啈=�ٿ��zO��@�؉!4@�bz�0�!?�Z��˴@啈=�ٿ��zO��@�؉!4@�bz�0�!?�Z��˴@�#��ٿys�����@��@��3@����c�!?e�$۪�@B� ���ٿ(D(��@Q�>��3@P��e�!?m�V�	�@��蛷�ٿ\ *?�g�@[�0��3@�rl5��!?P-�h��@bpp��ٿ{Cˠ��@ks8Z� 4@=	m�!?<׎�짴@�Ԥ��ٿ�MS����@��|z	4@������!?��=��@�Ԥ��ٿ�MS����@��|z	4@������!?��=��@�Ԥ��ٿ�MS����@��|z	4@������!?��=��@�Ԥ��ٿ�MS����@��|z	4@������!?��=��@�Ԥ��ٿ�MS����@��|z	4@������!?��=��@;�<�ٿ� C��@I�Lp4�3@�,"ɐ!?�K_����@;�<�ٿ� C��@I�Lp4�3@�,"ɐ!?�K_����@`b㻑ٿ�cδg|�@���J��3@[(�M��!?���\��@`b㻑ٿ�cδg|�@���J��3@[(�M��!?���\��@����Ҍٿ�w|��@�2��|�3@����z�!?�o)��@����Ҍٿ�w|��@�2��|�3@����z�!?�o)��@����Ҍٿ�w|��@�2��|�3@����z�!?�o)��@����Ҍٿ�w|��@�2��|�3@����z�!?�o)��@5Į�ڏٿ]����@A����3@��o�!?� �#|�@5Į�ڏٿ]����@A����3@��o�!?� �#|�@5Į�ڏٿ]����@A����3@��o�!?� �#|�@5Į�ڏٿ]����@A����3@��o�!?� �#|�@5Į�ڏٿ]����@A����3@��o�!?� �#|�@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@~mK�ɓٿ���ߵ��@�R�h4@�i:�&�!?=)���@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@��;]�ٿ������@#��b
4@��N�Z�!?��y*�Y�@�X�m��ٿ�.�}��@��=�4@P_�)c�!?��3�0��@�X�m��ٿ�.�}��@��=�4@P_�)c�!?��3�0��@�X�m��ٿ�.�}��@��=�4@P_�)c�!?��3�0��@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@�9ʺ�ٿ��l���@��舳�3@)��(�!?9,���@��cC�ٿ/u<l��@������3@�DX[t�!?������@s���ٿ�+ji��@`�}T��3@�If9l�!?F�ܝ됴@s���ٿ�+ji��@`�}T��3@�If9l�!?F�ܝ됴@s���ٿ�+ji��@`�}T��3@�If9l�!?F�ܝ됴@W�!�6�ٿ� n,��@������3@���}�!?AX�Ҵ@W�!�6�ٿ� n,��@������3@���}�!?AX�Ҵ@W�!�6�ٿ� n,��@������3@���}�!?AX�Ҵ@>�Ot�ٿ�?vU���@�w���3@��*͏!?zmW.��@>�Ot�ٿ�?vU���@�w���3@��*͏!?zmW.��@>�Ot�ٿ�?vU���@�w���3@��*͏!?zmW.��@���{�ٿ�3 H�@��X��4@��*}�!?�Fnbv��@���{�ٿ�3 H�@��X��4@��*}�!?�Fnbv��@|�-��ٿ�Y����@�A!i��3@��o��!?�]!���@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@���BڝٿN
A���@��t�x�3@�x��2�!?�����@�-��ٿ�A�x�@��ް��3@��7��!?�?:�W��@�U$8c�ٿ��*���@��ܺK�3@T[1��!?K���Sյ@�U$8c�ٿ��*���@��ܺK�3@T[1��!?K���Sյ@�U$8c�ٿ��*���@��ܺK�3@T[1��!?K���Sյ@�8��c�ٿ�g�QSk�@�߰܏�3@E��!?���,�ĵ@�8��c�ٿ�g�QSk�@�߰܏�3@E��!?���,�ĵ@�8��c�ٿ�g�QSk�@�߰܏�3@E��!?���,�ĵ@�8��c�ٿ�g�QSk�@�߰܏�3@E��!?���,�ĵ@����e�ٿ{PNA�@���ܲ�3@�_M�j�!?�1�6��@����e�ٿ{PNA�@���ܲ�3@�_M�j�!?�1�6��@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@�G�䯞ٿVE>��d�@�{���3@�ޑ9�!?�q�í�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@���
ژٿi0��l
�@�N���3@�k�N@�!?��X�c�@诫��ٿ;1�m'_�@��$�3@�����!?n'�4'�@诫��ٿ;1�m'_�@��$�3@�����!?n'�4'�@诫��ٿ;1�m'_�@��$�3@�����!?n'�4'�@诫��ٿ;1�m'_�@��$�3@�����!?n'�4'�@�&0�]�ٿ�0�+L�@l���3@=�/�!?X���ȅ�@Yk!��ٿ'"=�ֽ�@�?�`�3@�uS�9�!?Kt����@r�݌ٿ��8C�@:���3@$�"��!?�ĪY�@r�݌ٿ��8C�@:���3@$�"��!?�ĪY�@��D�ٿ���v��@5����3@���֏!?�Q2Iy�@��D�ٿ���v��@5����3@���֏!?�Q2Iy�@��D�ٿ���v��@5����3@���֏!?�Q2Iy�@��D�ٿ���v��@5����3@���֏!?�Q2Iy�@��D�ٿ���v��@5����3@���֏!?�Q2Iy�@�#�֚ٿ]6��@���Z�3@q��2�!?Ń1�9�@�m�1ޒٿ:���1�@S{��	4@�vi��!?���G��@�m�1ޒٿ:���1�@S{��	4@�vi��!?���G��@|��hq�ٿ�@fh��@�;b��3@�R&��!?f�9�@|��hq�ٿ�@fh��@�;b��3@�R&��!?f�9�@/��J�ٿw��4Ż�@�mЩ�3@��{�<�!?	��f�@/��J�ٿw��4Ż�@�mЩ�3@��{�<�!?	��f�@/��J�ٿw��4Ż�@�mЩ�3@��{�<�!?	��f�@�U`��ٿ؉���@�䐻��3@9�e��!?�1�[��@�U`��ٿ؉���@�䐻��3@9�e��!?�1�[��@g��7݌ٿ�`~��@*^i	��3@j�7P�!?QCQՖM�@B��ߓٿ�Bc�t�@�����3@�� �D�!?������@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@� /飗ٿ�������@'6e��3@���h/�!?�6�-�@	�nZ��ٿF�Ԉ��@�;�� 4@Ɣ� �!?��:hSĴ@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@h2%�~�ٿ^V��A�@�Y7#��3@L_�Q�!?T���ʖ�@���tC�ٿ��/ �)�@�q�3	4@%U�Da�!?q �ߴ@���tC�ٿ��/ �)�@�q�3	4@%U�Da�!?q �ߴ@��+�ٿ�r�#j��@8�����3@��;>�!?]��0�@��+�ٿ�r�#j��@8�����3@��;>�!?]��0�@��+�ٿ�r�#j��@8�����3@��;>�!?]��0�@��+�ٿ�r�#j��@8�����3@��;>�!?]��0�@�6�*�ٿ��a��@c�����3@e]5/�!?:�C1�;�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@���f��ٿ�����@l�GI� 4@����X�!?�ɘ2�@|����ٿ	��k�@\��W|�3@�|��@�!?��k@u�@|����ٿ	��k�@\��W|�3@�|��@�!?��k@u�@|����ٿ	��k�@\��W|�3@�|��@�!?��k@u�@L����ٿ���?��@_�mR��3@�S�;�!?U\B�k�@L����ٿ���?��@_�mR��3@�S�;�!?U\B�k�@L����ٿ���?��@_�mR��3@�S�;�!?U\B�k�@L����ٿ���?��@_�mR��3@�S�;�!?U\B�k�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�C�"��ٿ�Q2%��@�����3@�кj>�!?�T6S�@�k��s�ٿ�Z�_R}�@[���3@9�}AT�!?�'e�c��@�k��s�ٿ�Z�_R}�@[���3@9�}AT�!?�'e�c��@(�3@z�ٿ!HD���@W�!.��3@��6@�!?�%����@(�3@z�ٿ!HD���@W�!.��3@��6@�!?�%����@(�3@z�ٿ!HD���@W�!.��3@��6@�!?�%����@(�3@z�ٿ!HD���@W�!.��3@��6@�!?�%����@(�3@z�ٿ!HD���@W�!.��3@��6@�!?�%����@���_۔ٿ=���^�@F
m�3@�[�!�!?�8�X��@���_۔ٿ=���^�@F
m�3@�[�!�!?�8�X��@���_۔ٿ=���^�@F
m�3@�[�!�!?�8�X��@=dĒٿ��Z�:��@$ƞf��3@q�sGM�!?�����!�@��"�y�ٿ/��6��@�L����3@ZtS�!?�7Z��@P~[���ٿ5�V��8�@}n��3@�VĆ�!?�Z֗�@P~[���ٿ5�V��8�@}n��3@�VĆ�!?�Z֗�@P~[���ٿ5�V��8�@}n��3@�VĆ�!?�Z֗�@P~[���ٿ5�V��8�@}n��3@�VĆ�!?�Z֗�@P~[���ٿ5�V��8�@}n��3@�VĆ�!?�Z֗�@����r�ٿ�HU��1�@�^�|��3@�
��B�!?{TBP�>�@����r�ٿ�HU��1�@�^�|��3@�
��B�!?{TBP�>�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@�̜��ٿ��@��<�6�3@b���_�!?�;�ˀH�@��j�ٿ�)�^qb�@�H
Ǩ�3@2A�C�!?���t��@��j�ٿ�)�^qb�@�H
Ǩ�3@2A�C�!?���t��@��j�ٿ�)�^qb�@�H
Ǩ�3@2A�C�!?���t��@��j�ٿ�)�^qb�@�H
Ǩ�3@2A�C�!?���t��@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@uԈ�ٿ�J�-�@$\�d�3@����!?�����$�@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@y�ٿ�8ѡ�@�.���3@K9=��!?*{��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@��;W�ٿkSq~��@"�z��3@���J�!?��
�z��@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@D��Q�ٿپ}�v�@X&�3��3@Q��Lޏ!?�*�~�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@�U�V�ٿ���yV�@"���;�3@�sfw1�!?_ٹڿ8�@��G�șٿ�bJ����@I�i��3@�\�yk�!?�S��<�@���G��ٿ��TsgT�@ďٿ��3@*%>B�!?��~�@���G��ٿ��TsgT�@ďٿ��3@*%>B�!?��~�@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@����X�ٿ�]鿪��@�����3@Io0�<�!?��Ѫx��@7�rx�ٿ?�%��@1Ք�e�3@�l�\<�!?��6���@7�rx�ٿ?�%��@1Ք�e�3@�l�\<�!?��6���@��ÿB�ٿ�K썈�@U�*y�3@�� FD�!?W��@�oo\�ٿ�g�p3�@Cz�`�3@/hZ�@�!?|;lsʹ@�oo\�ٿ�g�p3�@Cz�`�3@/hZ�@�!?|;lsʹ@�oo\�ٿ�g�p3�@Cz�`�3@/hZ�@�!?|;lsʹ@�����ٿ�m�N��@,��3@�H�E�!?2zb�!L�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@*d�=��ٿ������@�WL�3@{H_�~�!?����)X�@vL�ݝٿPʌ.���@L%����3@)���y�!?V 䧜�@o{���ٿ�び��@l�l���3@�X5	F�!?��'u�V�@o{���ٿ�び��@l�l���3@�X5	F�!?��'u�V�@��u�ٿ���`L�@��M�4@v�Y�!?$OreC��@��u�ٿ���`L�@��M�4@v�Y�!?$OreC��@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@�WT�ٿ���W l�@����\�3@��[m�!?L�V�ƴ@wP�י�ٿ�!�T��@ `�1%�3@��vw�!?���f��@wP�י�ٿ�!�T��@ `�1%�3@��vw�!?���f��@wP�י�ٿ�!�T��@ `�1%�3@��vw�!?���f��@wP�י�ٿ�!�T��@ `�1%�3@��vw�!?���f��@�D�Ϛٿt�8¥�@-�W�`�3@��L��!?�q�~�е@܄l} �ٿnӔx=�@�(���3@F���!?�����@Q����ٿ���si��@_�u
��3@"�0��!?gk$m�Y�@Q����ٿ���si��@_�u
��3@"�0��!?gk$m�Y�@Q����ٿ���si��@_�u
��3@"�0��!?gk$m�Y�@Q����ٿ���si��@_�u
��3@"�0��!?gk$m�Y�@Q����ٿ���si��@_�u
��3@"�0��!?gk$m�Y�@�,��͔ٿ�ˀv���@�Ʋ���3@8zw��!?[����>�@�,��͔ٿ�ˀv���@�Ʋ���3@8zw��!?[����>�@�,��͔ٿ�ˀv���@�Ʋ���3@8zw��!?[����>�@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@���� �ٿ "����@� �
}�3@�5P��!?���	��@�0��v�ٿC��i<�@�ۖ�t�3@ҍ���!?�0v_�ݴ@ �Sұ�ٿ^�\�_��@k��{�3@��0|�!?��� �@ �Sұ�ٿ^�\�_��@k��{�3@��0|�!?��� �@ �Sұ�ٿ^�\�_��@k��{�3@��0|�!?��� �@����3�ٿ ����y�@F�vJ�3@A���O�!?z����@����3�ٿ ����y�@F�vJ�3@A���O�!?z����@+���d�ٿ��):;�@�y2�
�3@�,��N�!?K���.�@+���d�ٿ��):;�@�y2�
�3@�,��N�!?K���.�@+���d�ٿ��):;�@�y2�
�3@�,��N�!?K���.�@���b�ٿ����s�@0o�(4@d�Z=�!?��V#��@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@�Í$�ٿ"RBc4;�@�:Hg 4@�5�+R�!?GO�X�@��c�s�ٿ=���I�@��� 4@�p-B�!?���@��c�s�ٿ=���I�@��� 4@�p-B�!?���@x���ٿr����@��94@%���e�!?O��E�ƴ@x���ٿr����@��94@%���e�!?O��E�ƴ@x���ٿr����@��94@%���e�!?O��E�ƴ@x���ٿr����@��94@%���e�!?O��E�ƴ@x���ٿr����@��94@%���e�!?O��E�ƴ@x���ٿr����@��94@%���e�!?O��E�ƴ@O����ٿ!oz�0��@��Z�3@�$��?�!?~�h���@O����ٿ!oz�0��@��Z�3@�$��?�!?~�h���@O����ٿ!oz�0��@��Z�3@�$��?�!?~�h���@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@�8W0�ٿո�S�@.u"*��3@Y�}
k�!?���S�@ &���ٿ�q�����@3��pm�3@��X�9�!?̠��$Y�@ &���ٿ�q�����@3��pm�3@��X�9�!?̠��$Y�@���k:�ٿ��ϗ���@g���3@�Q8J)�!?���?��@NR'p�ٿd����D�@9�_k��3@O�I��!?2٧z�O�@L���S�ٿ���mr��@�R:���3@�0S�ڏ!?�>�h���@L���S�ٿ���mr��@�R:���3@�0S�ڏ!?�>�h���@�e	ӳ�ٿ������@E�.���3@
�>T�!?��0��j�@�e	ӳ�ٿ������@E�.���3@
�>T�!?��0��j�@�e	ӳ�ٿ������@E�.���3@
�>T�!?��0��j�@�e	ӳ�ٿ������@E�.���3@
�>T�!?��0��j�@�J�Ŭ�ٿ�4����@y��\�3@����.�!?.�H�\�@?���[�ٿS��&�{�@v�!��3@��q���!?�pT ��@?���[�ٿS��&�{�@v�!��3@��q���!?�pT ��@?���[�ٿS��&�{�@v�!��3@��q���!?�pT ��@4�$Jp�ٿ��{���@�M���3@���o��!?!���-�@4�$Jp�ٿ��{���@�M���3@���o��!?!���-�@4�$Jp�ٿ��{���@�M���3@���o��!?!���-�@�ia�ٿ�dm��+�@�}����3@m��uU�!?��Knֵ@�m��ŏٿ݈��U�@���V��3@\~?OW�!?�]'���@�m��ŏٿ݈��U�@���V��3@\~?OW�!?�]'���@�m��ŏٿ݈��U�@���V��3@\~?OW�!?�]'���@�m��ŏٿ݈��U�@���V��3@\~?OW�!?�]'���@�_�p�ٿ�K@�M�@�/A�3@����&�!?��W7>�@��@�!�ٿR��Eq�@�v 4�3@o$�� �!?m��9B#�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@&Ag�ݖٿ�Af}p�@Nsc�G�3@��� ?�!?�� �_�@�׸I��ٿki��K��@�����3@�uo�i�!?Y��/�@���6q�ٿ����.�@l���3@5X8z�!?�Pٓ�6�@���6q�ٿ����.�@l���3@5X8z�!?�Pٓ�6�@R}ݞŗٿf�C�E�@b�9���3@8�H%z�!?�!����@R}ݞŗٿf�C�E�@b�9���3@8�H%z�!?�!����@R}ݞŗٿf�C�E�@b�9���3@8�H%z�!?�!����@���BT�ٿ�߽W���@lx�M^�3@V~�(�!?�$��ެ�@���BT�ٿ�߽W���@lx�M^�3@V~�(�!?�$��ެ�@A	⪰�ٿ�c�%.��@Q��>�3@[��97�!?ֲ��#�@��=\�ٿ�-��X�@S���K�3@@+vw�!?ku��*�@��=\�ٿ�-��X�@S���K�3@@+vw�!?ku��*�@��=\�ٿ�-��X�@S���K�3@@+vw�!?ku��*�@��=\�ٿ�-��X�@S���K�3@@+vw�!?ku��*�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�F|��ٿ	����@� V��3@TN,l�!?eK���>�@�tG� �ٿaU�u.��@�"W��3@�X�E�!?OtC�@�@�tG� �ٿaU�u.��@�"W��3@�X�E�!?OtC�@�@�tG� �ٿaU�u.��@�"W��3@�X�E�!?OtC�@�@�Y��9�ٿ�A��qp�@�nF�z�3@�
.ʏ!?�Y�b}�@�Y��9�ٿ�A��qp�@�nF�z�3@�
.ʏ!?�Y�b}�@�Y��9�ٿ�A��qp�@�nF�z�3@�
.ʏ!?�Y�b}�@�Y��9�ٿ�A��qp�@�nF�z�3@�
.ʏ!?�Y�b}�@�Y��9�ٿ�A��qp�@�nF�z�3@�
.ʏ!?�Y�b}�@u��x�ٿ�3��d��@�ă��3@'i�7ԏ!?|╳��@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�=��ٿ���=�@�.:t�3@�4�ߏ!?���)δ@�:�$�ٿ2��#�@����3@4��u�!?�ꚞ�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@��?M�ٿ;���@"����3@AC(s�!?�I�+|�@ڈ���ٿ S���c�@'��D}�3@I9��n�!?!H@w� �@t!*�p�ٿ�c	;���@!�p��3@o�T5�!?v~���@���f��ٿ��%����@���r�3@�	�p��!?�&=|b��@���f��ٿ��%����@���r�3@�	�p��!?�&=|b��@���f��ٿ��%����@���r�3@�	�p��!?�&=|b��@���f��ٿ��%����@���r�3@�	�p��!?�&=|b��@Jeu�ٿTk4$��@ms�	��3@�ܖ�q�!?5�r�P�@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@²E�*�ٿ��]V��@�PT��3@ýP4��!?�W���@.��F�ٿ<_�����@\��(i�3@Nޱ�	�!?��⭴@.��F�ٿ<_�����@\��(i�3@Nޱ�	�!?��⭴@.��F�ٿ<_�����@\��(i�3@Nޱ�	�!?��⭴@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@�ў��ٿ"�/Na��@��yup�3@b7��P�!?z鍓��@��P��ٿ�iMkS�@~��T�3@R����!?e	qڈ��@��P��ٿ�iMkS�@~��T�3@R����!?e	qڈ��@��	���ٿ���nJ�@8�l���3@g
�F��!?��gH��@��	���ٿ���nJ�@8�l���3@g
�F��!?��gH��@��	���ٿ���nJ�@8�l���3@g
�F��!?��gH��@��	���ٿ���nJ�@8�l���3@g
�F��!?��gH��@��	���ٿ���nJ�@8�l���3@g
�F��!?��gH��@U��zG�ٿ�O���@���Ě�3@qN�9�!?J|xx(�@U��zG�ٿ�O���@���Ě�3@qN�9�!?J|xx(�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@�V[��ٿ�Ֆ?�@r>�.�3@�K{K�!?�^��a�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@V���Öٿ	�m��W�@�M��_�3@��`�!?�S;-�@䥹���ٿ��hP��@}˄���3@��Gzj�!?��Y��@䥹���ٿ��hP��@}˄���3@��Gzj�!?��Y��@䥹���ٿ��hP��@}˄���3@��Gzj�!?��Y��@䥹���ٿ��hP��@}˄���3@��Gzj�!?��Y��@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@
���7�ٿ�=H`�@`1���3@c��9�!?�VkbXm�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�O��q�ٿ���	�$�@�:���3@uⱒm�!?����F�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@�t�2J�ٿ<Þך�@���M�3@�2��W�!?5|5�ar�@��&D�ٿ����O��@S�����3@+�хz�!?����KI�@%��ٿ� }�С�@�{���3@&��א!?
�gB�@W2�?%�ٿ�K�f��@������3@��i͐!?C�N�۴@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@GG�ٿr���Z��@@�ݿ�3@���դ�!?[(մ@c���ٿ�E��+�@2G����3@���!?�=++7,�@c���ٿ�E��+�@2G����3@���!?�=++7,�@c���ٿ�E��+�@2G����3@���!?�=++7,�@c���ٿ�E��+�@2G����3@���!?�=++7,�@�o����ٿ��KF���@?yFi�4@��
%��!?b1���5�@h�x�ٿ���X8�@����4@���\u�!?P��PA2�@h�x�ٿ���X8�@����4@���\u�!?P��PA2�@��eҔٿ����X�@�x�$T�3@_�PUЏ!?e�mM��@��eҔٿ����X�@�x�$T�3@_�PUЏ!?e�mM��@��eҔٿ����X�@�x�$T�3@_�PUЏ!?e�mM��@��eҔٿ����X�@�x�$T�3@_�PUЏ!?e�mM��@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@7�07��ٿ�]C2���@.��Bw�3@�l�dM�!?��o��ѵ@�N���ٿ��eCK��@3�O�3�3@�W��I�!?A*�C=��@�N���ٿ��eCK��@3�O�3�3@�W��I�!?A*�C=��@�N���ٿ��eCK��@3�O�3�3@�W��I�!?A*�C=��@}?4=N�ٿ�QZu��@v�0�3@�:-�D�!?��7����@}?4=N�ٿ�QZu��@v�0�3@�:-�D�!?��7����@}?4=N�ٿ�QZu��@v�0�3@�:-�D�!?��7����@}?4=N�ٿ�QZu��@v�0�3@�:-�D�!?��7����@}?4=N�ٿ�QZu��@v�0�3@�:-�D�!?��7����@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@6���}�ٿ�;i���@y���3@�^�I8�!?�0�>��@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@����@�ٿ��3���@Se���3@9D����!?�>���@���mj�ٿ�a��x�@q�����3@#Q�l��!?6���r�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@���QǗٿ�$,�!n�@�A��b�3@T�"&��!?���ԏ7�@�H�<�ٿR�_��/�@�M!�3@�&��z�!?���8M�@�H�<�ٿR�_��/�@�M!�3@�&��z�!?���8M�@�H�<�ٿR�_��/�@�M!�3@�&��z�!?���8M�@���䛒ٿ�2�E�u�@�=�,��3@6�Ҙ8�!?�� tj��@���䛒ٿ�2�E�u�@�=�,��3@6�Ҙ8�!?�� tj��@���䛒ٿ�2�E�u�@�=�,��3@6�Ҙ8�!?�� tj��@Q���:�ٿeV"�r�@yC�j�3@{�T�H�!?�"$�* �@Q���:�ٿeV"�r�@yC�j�3@{�T�H�!?�"$�* �@Q���:�ٿeV"�r�@yC�j�3@{�T�H�!?�"$�* �@>�̜��ٿ��$ˤ!�@���T�3@ޮ�K�!?��㫴@>�̜��ٿ��$ˤ!�@���T�3@ޮ�K�!?��㫴@>�̜��ٿ��$ˤ!�@���T�3@ޮ�K�!?��㫴@>�̜��ٿ��$ˤ!�@���T�3@ޮ�K�!?��㫴@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@~_��ٿ$9lb��@����X�3@�1��!?TR�9�@�5��ٿ�D&�5��@:��c��3@���n�!?'PB}]t�@a�!� �ٿΪ���*�@���9�3@ ��G�!?�E��s��@a�!� �ٿΪ���*�@���9�3@ ��G�!?�E��s��@a�!� �ٿΪ���*�@���9�3@ ��G�!?�E��s��@���ٿ�TE�]Y�@sD��[�3@GI�A�!?r�b~�g�@���ٿ�TE�]Y�@sD��[�3@GI�A�!?r�b~�g�@���ٿ�TE�]Y�@sD��[�3@GI�A�!?r�b~�g�@(>��ٿw!�?�^�@��Q���3@��x��!?\���@(>��ٿw!�?�^�@��Q���3@��x��!?\���@(>��ٿw!�?�^�@��Q���3@��x��!?\���@(>��ٿw!�?�^�@��Q���3@��x��!?\���@(>��ٿw!�?�^�@��Q���3@��x��!?\���@(>��ٿw!�?�^�@��Q���3@��x��!?\���@��F���ٿ�Z���@�#<��3@�8�<�!?�]�j�h�@��F���ٿ�Z���@�#<��3@�8�<�!?�]�j�h�@�����ٿN�؀��@+𙞒�3@%�� �!?�������@�����ٿN�؀��@+𙞒�3@%�� �!?�������@�����ٿN�؀��@+𙞒�3@%�� �!?�������@�z���ٿ���9�@Q�6�3@?�CǏ!?�ʞ�`W�@`�mB>�ٿ�]��k�@�h��� 4@<�����!?%<�;�@`�mB>�ٿ�]��k�@�h��� 4@<�����!?%<�;�@!;%���ٿE��o�}�@�ې���3@��3�x�!?v��H�H�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@|�,��ٿ�����@��n`N�3@:�<�[�!?��d�@�	d{��ٿ�`͏h��@<�,C�3@oz>k�!?AZµ@��?�ٿM������@<b+m4@,[�V'�!?ܶ����@��?�ٿM������@<b+m4@,[�V'�!?ܶ����@�4����ٿ��þ7�@���D��3@�����!?�[ѳx�@�4����ٿ��þ7�@���D��3@�����!?�[ѳx�@�4����ٿ��þ7�@���D��3@�����!?�[ѳx�@�4����ٿ��þ7�@���D��3@�����!?�[ѳx�@�4����ٿ��þ7�@���D��3@�����!?�[ѳx�@k�+�O�ٿ��"d>w�@�t��3@�a�b�!?+KM���@k�+�O�ٿ��"d>w�@�t��3@�a�b�!?+KM���@k�+�O�ٿ��"d>w�@�t��3@�a�b�!?+KM���@k�+�O�ٿ��"d>w�@�t��3@�a�b�!?+KM���@C�y�3�ٿ���#�@�����3@��G�c�!?��M�6��@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@@�F�ٿ����_.�@�M�15�3@�	uM�!?v���ϵ@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@�+.�ٿ��Z�]�@��C��3@GV
�/�!?'�@P.��@2?�àٿH}Gl�f�@�!*�-�3@*o�d�!?\��<m�@2?�àٿH}Gl�f�@�!*�-�3@*o�d�!?\��<m�@2?�àٿH}Gl�f�@�!*�-�3@*o�d�!?\��<m�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@M;&O�ٿ^�E��^�@nT�y-	4@�=�Q�!?���qG�@��!�ٿ���ޮ��@͓p"4@�龝�!?�=o���@��!�ٿ���ޮ��@͓p"4@�龝�!?�=o���@��6��ٿ"�7#�f�@�!�nn4@�0�,�!?�p�q��@�s�z��ٿ��b�5��@�C�E��3@S��!?xgFD&ֵ@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@Pqղ�ٿq ߵ���@8o���3@�GG\�!?OJ6��@�̿繓ٿ��)����@ǆ}hX�3@0a	�!?V�4C烵@�̿繓ٿ��)����@ǆ}hX�3@0a	�!?V�4C烵@�̿繓ٿ��)����@ǆ}hX�3@0a	�!?V�4C烵@PG�)��ٿxF��}��@?E6�h�3@��{�+�!?�_]g�Ҵ@PG�)��ٿxF��}��@?E6�h�3@��{�+�!?�_]g�Ҵ@�^��ٿ$�� /m�@�/
4@/ؙ=�!?A? ���@�^��ٿ$�� /m�@�/
4@/ؙ=�!?A? ���@�^��ٿ$�� /m�@�/
4@/ؙ=�!?A? ���@�^��ٿ$�� /m�@�/
4@/ؙ=�!?A? ���@����l�ٿ�H_��@�/����3@�}z�ŏ!?B(;���@��� �ٿ4��:T�@W����3@��<���!?C���̵@��� �ٿ4��:T�@W����3@��<���!?C���̵@��� �ٿ4��:T�@W����3@��<���!?C���̵@����ٿ� Gz �@*B<���3@����s�!?�L7�F��@J&�d�ٿ�<���@}?*�3@����!?��H���@J&�d�ٿ�<���@}?*�3@����!?��H���@J&�d�ٿ�<���@}?*�3@����!?��H���@J&�d�ٿ�<���@}?*�3@����!?��H���@J&�d�ٿ�<���@}?*�3@����!?��H���@J&�d�ٿ�<���@}?*�3@����!?��H���@x=����ٿg1�.��@9b�J�3@��0Bv�!?��-��@x=����ٿg1�.��@9b�J�3@��0Bv�!?��-��@x=����ٿg1�.��@9b�J�3@��0Bv�!?��-��@���E�ٿK����@��=0�3@���!?�i%�O��@���E�ٿK����@��=0�3@���!?�i%�O��@���E�ٿK����@��=0�3@���!?�i%�O��@���E�ٿK����@��=0�3@���!?�i%�O��@���E�ٿK����@��=0�3@���!?�i%�O��@�G�V��ٿ�����@#�m��4@��_��!?���Ĵ�@�G�V��ٿ�����@#�m��4@��_��!?���Ĵ�@�G�V��ٿ�����@#�m��4@��_��!?���Ĵ�@�G�V��ٿ�����@#�m��4@��_��!?���Ĵ�@�G�V��ٿ�����@#�m��4@��_��!?���Ĵ�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@�-���ٿ���%�/�@`�lq�3@f��$�!?�qqװ|�@E�W���ٿy3~�-c�@����h�3@��h�!?�ΛjHI�@E�W���ٿy3~�-c�@����h�3@��h�!?�ΛjHI�@E�W���ٿy3~�-c�@����h�3@��h�!?�ΛjHI�@�V��ٿ�1���@��b�[�3@�I�)3�!?(]3���@�)]W��ٿϘ��<��@���j��3@���v�!?��g�<۳@�<S�ٿ P��&�@�}i�K�3@��v<��!?�,w�Z�@�<S�ٿ P��&�@�}i�K�3@��v<��!?�,w�Z�@�<S�ٿ P��&�@�}i�K�3@��v<��!?�,w�Z�@��S��ٿ�F��&|�@H��m�3@����#�!?t�� �3�@��S��ٿ�F��&|�@H��m�3@����#�!?t�� �3�@|�@K�ٿ���@�('�3@�#�J�!?`nNyet�@|�@K�ٿ���@�('�3@�#�J�!?`nNyet�@|�@K�ٿ���@�('�3@�#�J�!?`nNyet�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@9c| H�ٿN�>��x�@<����3@r�wlJ�!?F�]��K�@�<�L��ٿ����j�@����3@���E��!?��b�F$�@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@���1h�ٿt��<'�@�;94@@Up�g�!?�dD����@x�d�ٿ���L��@�S+���3@�=#��!?VI��R�@x�d�ٿ���L��@�S+���3@�=#��!?VI��R�@x���әٿcz����@�<���3@Q)x��!?�4]2�<�@x���әٿcz����@�<���3@Q)x��!?�4]2�<�@x���әٿcz����@�<���3@Q)x��!?�4]2�<�@x���әٿcz����@�<���3@Q)x��!?�4]2�<�@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@��7�N�ٿ7Nm*��@wV�)��3@b?�!?��1��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@ȏ5�ʘٿ����Ũ�@vQ{l�3@EnVֶ�!?�X�Q��@�����ٿ�y�X4��@^)�͘4@��6��!?��)��@�5<�ٿc+d��@��I�4@J�sA �!?ˋ���w�@��=��ٿ�0����@A����3@0S?��!?*��x��@��=��ٿ�0����@A����3@0S?��!?*��x��@��=��ٿ�0����@A����3@0S?��!?*��x��@��=��ٿ�0����@A����3@0S?��!?*��x��@���W��ٿ�N�9��@ьtsJ�3@A����!?]��@���W��ٿ�N�9��@ьtsJ�3@A����!?]��@���:�ٿ;�6ō�@�P�/5�3@ſ�Yz�!?���	d�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@L�*'y�ٿ�*����@-�<��3@��u�@�!?i���h�@�ڋNM�ٿ��y�a��@B���n�3@`�����!?���M�@�ڋNM�ٿ��y�a��@B���n�3@`�����!?���M�@�ڋNM�ٿ��y�a��@B���n�3@`�����!?���M�@�ڋNM�ٿ��y�a��@B���n�3@`�����!?���M�@�ڋNM�ٿ��y�a��@B���n�3@`�����!?���M�@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@˻���ٿ�g���@��D��3@M��!?�'�=۵@��C���ٿ����@Zy��3@t�	
�!?L��&i�@��C���ٿ����@Zy��3@t�	
�!?L��&i�@�2Ie�ٿ�X'�_�@��B���3@�Z��S�!?�N�_�@�2Ie�ٿ�X'�_�@��B���3@�Z��S�!?�N�_�@�2Ie�ٿ�X'�_�@��B���3@�Z��S�!?�N�_�@�2Ie�ٿ�X'�_�@��B���3@�Z��S�!?�N�_�@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@�����ٿ��
��@I?{�3@�4�|Y�!?� ����@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@\+���ٿ��g��{�@nyjo��3@�Ԩ�h�!?�׮�C�@!PI�N�ٿ��#h��@@��a�3@�\]�!?�Z�,�*�@!PI�N�ٿ��#h��@@��a�3@�\]�!?�Z�,�*�@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@�^(�ٿ��2��@I�mzV�3@�����!?\ ����@[��5�ٿ3�9�w�@џUML�3@P���	�!?�w3�(�@[��5�ٿ3�9�w�@џUML�3@P���	�!?�w3�(�@^3df�ٿ=v�	�@W�U�3@����!?�>�WG�@^3df�ٿ=v�	�@W�U�3@����!?�>�WG�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�γE�ٿz����@���I�3@L���z�!?�J��"�@�#�N�ٿ|�Y����@�֒��3@o�An�!?(en@u�@�#�N�ٿ|�Y����@�֒��3@o�An�!?(en@u�@�#�N�ٿ|�Y����@�֒��3@o�An�!?(en@u�@�#�N�ٿ|�Y����@�֒��3@o�An�!?(en@u�@�Bo��ٿ�Ӎ���@c�����3@�y�P�!?�k�$!��@�Bo��ٿ�Ӎ���@c�����3@�y�P�!?�k�$!��@�Bo��ٿ�Ӎ���@c�����3@�y�P�!?�k�$!��@����ٿ
k+b�@������3@ҷ�Rx�!?	�'Ե@����ٿ
k+b�@������3@ҷ�Rx�!?	�'Ե@����ٿ
k+b�@������3@ҷ�Rx�!?	�'Ե@������ٿC�W��K�@�V�S3�3@C��H�!?�*����@�1�;�ٿdV�@���
��3@j�13�!?|ͺ ��@���z�ٿGt�1��@�r�3@��J�,�!?��$��@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@�/	�`�ٿ�c�D�b�@�����3@o���U�!?�>�Yõ@����ٿ��3z4k�@��ȷ.�3@|��u�!?���@��@����ٿ��3z4k�@��ȷ.�3@|��u�!?���@��@����ٿ��3z4k�@��ȷ.�3@|��u�!?���@��@T��U�ٿf�.`	�@��|��3@�Z���!?����Q�@T��U�ٿf�.`	�@��|��3@�Z���!?����Q�@T��U�ٿf�.`	�@��|��3@�Z���!?����Q�@T��U�ٿf�.`	�@��|��3@�Z���!?����Q�@��r �ٿ�v�?z�@=��f��3@}a4s�!?�w�HqI�@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@$�>P�ٿ)�cG���@yIjV�3@��NL8�!?������@����ٿ�C�b���@ �Ԍt�3@�����!?���0���@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�o��ϑٿ btvl�@��Ԏ��3@(��&�!?��IP�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@�����ٿS��ؗ��@M�vP�3@�u'�!?�0=�Δ�@l����ٿY0]���@pj�vK�3@~m�=/�!?���	�@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@D�YO��ٿF́x�@��<lR4@Y.@��!?�;����@�b���ٿP����@P��p"�3@��'G!?]�� |�@���Џ�ٿ��a�@߭��q�3@���R�!?>��s��@���Џ�ٿ��a�@߭��q�3@���R�!?>��s��@����ƕٿ-w=O�@�χ���3@2yoL/�!?v]�t��@����ƕٿ-w=O�@�χ���3@2yoL/�!?v]�t��@��'(f�ٿ�=����@��j�6�3@�f��!?�b��@��'(f�ٿ�=����@��j�6�3@�f��!?�b��@��'(f�ٿ�=����@��j�6�3@�f��!?�b��@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@U]��m�ٿy�ב5��@;̊�$�3@��e �!?t� �#�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@�,M�ٿ��l���@��-�3@g��k�!?���e�@���Ps�ٿ���+���@Ce���3@����!?ł�7��@�ro)Ŏٿh?����@\��U�3@P��!?϶	ƨ�@�ro)Ŏٿh?����@\��U�3@P��!?϶	ƨ�@�ro)Ŏٿh?����@\��U�3@P��!?϶	ƨ�@����@�ٿ�y�!H�@@�#Q� 4@�X�ؐ!?�{����@����@�ٿ�y�!H�@@�#Q� 4@�X�ؐ!?�{����@����@�ٿ�y�!H�@@�#Q� 4@�X�ؐ!?�{����@����@�ٿ�y�!H�@@�#Q� 4@�X�ؐ!?�{����@����@�ٿ�y�!H�@@�#Q� 4@�X�ؐ!?�{����@���u�ٿ�����@���\�4@�����!?�#/���@��G���ٿ*���=�@�ި<4@�꿻w�!?8V}q�@��G���ٿ*���=�@�ި<4@�꿻w�!?8V}q�@��G���ٿ*���=�@�ި<4@�꿻w�!?8V}q�@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@֧����ٿFy@�R�@��)���3@�8٠w�!?��45 �@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@,��ޖٿ�q�����@-�r��3@��u`�!?"ح�ʴ@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@s�����ٿ��0;�s�@_{W�Z�3@R��3I�!?|��E��@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@��2�ٿG>����@�3�e�3@�/��!?�T����@Z�9Z��ٿ�
"Y�@�K��3@��z�!?p�N�q�@1�؅P�ٿR$���@�H	|��3@�Cᇐ!?]1p�p<�@1�؅P�ٿR$���@�H	|��3@�Cᇐ!?]1p�p<�@1�؅P�ٿR$���@�H	|��3@�Cᇐ!?]1p�p<�@1�؅P�ٿR$���@�H	|��3@�Cᇐ!?]1p�p<�@���;��ٿ����)|�@=u�]4@Dۄ?Z�!?����0��@���;��ٿ����)|�@=u�]4@Dۄ?Z�!?����0��@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@K԰��ٿ��u���@r��c�3@�φG�!?�r9�D1�@4]��ٿ�J��:�@cm���3@fLx� �!?��ǭ�@�j_�ٿަo���@h�h�`�3@R]n�!?Nw}��J�@�j_�ٿަo���@h�h�`�3@R]n�!?Nw}��J�@�j_�ٿަo���@h�h�`�3@R]n�!?Nw}��J�@�j_�ٿަo���@h�h�`�3@R]n�!?Nw}��J�@
���p�ٿγ��w��@��%�H�3@�ܧ���!?8�1�@
���p�ٿγ��w��@��%�H�3@�ܧ���!?8�1�@\'�J��ٿ����@�@fZ���4@K4*H�!?n�rm6�@\'�J��ٿ����@�@fZ���4@K4*H�!?n�rm6�@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@,�0~��ٿHG�$v��@`�E �3@��ܜc�!?��a�x��@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@(�C��ٿɃrpV_�@Q��'O�3@2��b�!?�Ԯ+2�@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@ �C$7�ٿ�ٶ65��@��\�3@�4�u��!?��\a���@�C���ٿr s
W�@�!�9�3@lM��!?9U��ܴ@��'�
�ٿ⓲	^�@i�+0�3@����Z�!?����@��1��ٿ$d����@��F:�3@6��Y�!?�{� nȴ@��1��ٿ$d����@��F:�3@6��Y�!?�{� nȴ@��1��ٿ$d����@��F:�3@6��Y�!?�{� nȴ@��1��ٿ$d����@��F:�3@6��Y�!?�{� nȴ@��1��ٿ$d����@��F:�3@6��Y�!?�{� nȴ@����ٿ�E&�ߔ�@��l���3@�֪v�!?�l@�l{�@����ٿ�E&�ߔ�@��l���3@�֪v�!?�l@�l{�@����ٿ�E&�ߔ�@��l���3@�֪v�!?�l@�l{�@2��'�ٿQ��[���@��P���3@��>-�!?��.���@2��'�ٿQ��[���@��P���3@��>-�!?��.���@2��'�ٿQ��[���@��P���3@��>-�!?��.���@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@��@�B�ٿ���g)�@G����3@�9 �<�!?#�<��@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@o,���ٿ�D��@'5����3@\��a�!?�
I7J�@���\�ٿ���ч�@Zg�́�3@��c�"�!?'�@���j̏ٿ�`^��@��p�3@��"*�!?+��K���@���j̏ٿ�`^��@��p�3@��"*�!?+��K���@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@bB�ݝ�ٿ>�G
��@�����3@���C�!?�Q_��1�@��1�ٿOD&7x��@*�^��3@�h�E�!?�ZlM��@��{ͬ�ٿ�ْu��@��sn��3@K�J�x�!?*�t���@��{ͬ�ٿ�ْu��@��sn��3@K�J�x�!?*�t���@��{ͬ�ٿ�ْu��@��sn��3@K�J�x�!?*�t���@��{ͬ�ٿ�ْu��@��sn��3@K�J�x�!?*�t���@k�w�ٿ�M8�ڬ�@����3@V�- ݐ!?Ŷa��^�@؞�j�ٿ�NR��L�@�26���3@k:[��!?�0��@؞�j�ٿ�NR��L�@�26���3@k:[��!?�0��@�}+��ٿj�,��g�@Xǁ)�3@[��7�!?�5/�*�@�}+��ٿj�,��g�@Xǁ)�3@[��7�!?�5/�*�@�}+��ٿj�,��g�@Xǁ)�3@[��7�!?�5/�*�@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@a4��k�ٿ�~�� ��@�L�}��3@��M�r�!?"2.���@�6��(�ٿ��N��@Q�/��3@X1�`��!?�8���@�6��(�ٿ��N��@Q�/��3@X1�`��!?�8���@�6��(�ٿ��N��@Q�/��3@X1�`��!?�8���@v��IR�ٿ�{E52|�@C��M��3@	���!?PN�]�@�����ٿ����3�@��B�r4@���5��!?3vc��@�����ٿ����3�@��B�r4@���5��!?3vc��@�����ٿ����3�@��B�r4@���5��!?3vc��@�����ٿ����3�@��B�r4@���5��!?3vc��@��.��ٿ�v.�z�@�����3@u�p&�!?g��k�@��.��ٿ�v.�z�@�����3@u�p&�!?g��k�@��.��ٿ�v.�z�@�����3@u�p&�!?g��k�@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@�����ٿ�H ���@�m�$��3@Xt��!?\�e�:��@>���ٿ������@)�*c
�3@I84z��!?��2��@>���ٿ������@)�*c
�3@I84z��!?��2��@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@$����ٿ���\H��@��@r�3@�P���!?r:���@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@����ٿ ��Z�@�f�e�3@������!?�J?6 ��@(����ٿ��@RO�@�7��3@9LlzV�!? ����@(����ٿ��@RO�@�7��3@9LlzV�!? ����@(����ٿ��@RO�@�7��3@9LlzV�!? ����@(����ٿ��@RO�@�7��3@9LlzV�!? ����@(����ٿ��@RO�@�7��3@9LlzV�!? ����@(����ٿ��@RO�@�7��3@9LlzV�!? ����@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@u"{��ٿ�(P��@FSao��3@@���1�!?����(��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@c6N�ٿT���/�@�G���3@�3RV�!?�C{��@Ԇ�<��ٿi���O�@��Ւ��3@��S_�!?c��l�@�eb�ٿ���,�@�a[��3@�˧WZ�!?��M�}��@�eb�ٿ���,�@�a[��3@�˧WZ�!?��M�}��@�eb�ٿ���,�@�a[��3@�˧WZ�!?��M�}��@�eb�ٿ���,�@�a[��3@�˧WZ�!?��M�}��@�eb�ٿ���,�@�a[��3@�˧WZ�!?��M�}��@��w.��ٿ����z��@r�h���3@Q5��3�!?�4ˮR%�@��w.��ٿ����z��@r�h���3@Q5��3�!?�4ˮR%�@��w.��ٿ����z��@r�h���3@Q5��3�!?�4ˮR%�@�[mi�ٿI0~�@�>���3@��R��!?Y��VL�@�[mi�ٿI0~�@�>���3@��R��!?Y��VL�@�[mi�ٿI0~�@�>���3@��R��!?Y��VL�@d�5�ƛٿZo]@y\�@~u���3@�{��W�!?����ݴ@d�5�ƛٿZo]@y\�@~u���3@�{��W�!?����ݴ@d�5�ƛٿZo]@y\�@~u���3@�{��W�!?����ݴ@d�5�ƛٿZo]@y\�@~u���3@�{��W�!?����ݴ@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@�{�T��ٿP�J�7<�@=0���3@�0��R�!?I��nd�@)`�r��ٿ���)�>�@��A$}�3@nc/��!?���cܵ@)`�r��ٿ���)�>�@��A$}�3@nc/��!?���cܵ@)`�r��ٿ���)�>�@��A$}�3@nc/��!?���cܵ@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@���c�ٿ���]��@E��*�3@�[�|�!?5�e�@ ���-�ٿJ�2`�5�@y`	���3@|�4O��!?n�p:��@�����ٿ��;�Q�@r�傹�3@��H�]�!?DA׿&J�@�����ٿ��;�Q�@r�傹�3@��H�]�!?DA׿&J�@)��P��ٿ(��>���@Q��#�3@� t㱐!?�ia=�@�g����ٿ�̩����@f ��|�3@�1`�P�!? ���(�@�g����ٿ�̩����@f ��|�3@�1`�P�!? ���(�@�g����ٿ�̩����@f ��|�3@�1`�P�!? ���(�@�g����ٿ�̩����@f ��|�3@�1`�P�!? ���(�@z'U���ٿ��JA�@[����3@�vE>�!?�L��)(�@�PWz�ٿ˗�u���@�M��3@Ә�yZ�!?\��j�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@�FZ�;�ٿ�c���@'T���3@x_���!?�6R~�=�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@`[���ٿJ���@�^�C
�3@z��t�!?8�-!B(�@}x��y�ٿ��p�ڂ�@��'�3@��$㬐!?'Φ=��@}x��y�ٿ��p�ڂ�@��'�3@��$㬐!?'Φ=��@}x��y�ٿ��p�ڂ�@��'�3@��$㬐!?'Φ=��@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@[ذ�Ҝٿ�㪮"�@�C��7�3@q�o.��!?��m-�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@������ٿ�T�Z��@��n�3@��ס'�!?���:�@�(cJ+�ٿ���N�@�o(p�3@cy�!?��ml~8�@�(cJ+�ٿ���N�@�o(p�3@cy�!?��ml~8�@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@��I/�ٿf!_�c�@ g��'�3@��n�w�!?�q�#ش@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@<����ٿM�<%���@Q���3@��,$�!?�EpI��@Kvf1��ٿ\}ar�@�ԛs�3@�K l�!?4��B�@Kvf1��ٿ\}ar�@�ԛs�3@�K l�!?4��B�@�nWm��ٿ�b+�]�@3�?��3@�UP�n�!?}����ʹ@Nϋ�S�ٿ������@c�o�6�3@^2	s�!?n��@Nϋ�S�ٿ������@c�o�6�3@^2	s�!?n��@���ٿ�~��@����3@+�D?�!?�>K�@��Jm*�ٿ�}�M��@Uu�{D�3@��çD�!?B�Ă�@��Jm*�ٿ�}�M��@Uu�{D�3@��çD�!?B�Ă�@��Jm*�ٿ�}�M��@Uu�{D�3@��çD�!?B�Ă�@��Jm*�ٿ�}�M��@Uu�{D�3@��çD�!?B�Ă�@S��w��ٿ� ��6�@!�C@@�3@I
�fo�!?�ԝ\�ʴ@S��w��ٿ� ��6�@!�C@@�3@I
�fo�!?�ԝ\�ʴ@n��nٿ�ki���@����3@٬X��!?bT2LI�@n��nٿ�ki���@����3@٬X��!?bT2LI�@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@종nޖٿ�`�n�@��O� �3@���r��!?�lF濴@���3֕ٿ�B�NE�@&e�	b�3@��,�N�!?P��ө��@{�#4�ٿ�q����@�)�u�3@�]t��!?!Y�ѫ�@{�#4�ٿ�q����@�)�u�3@�]t��!?!Y�ѫ�@{�#4�ٿ�q����@�)�u�3@�]t��!?!Y�ѫ�@{�#4�ٿ�q����@�)�u�3@�]t��!?!Y�ѫ�@�{����ٿr?oc��@�v����3@�߆�s�!?M�r04|�@�{����ٿr?oc��@�v����3@�߆�s�!?M�r04|�@�{����ٿr?oc��@�v����3@�߆�s�!?M�r04|�@�{����ٿr?oc��@�v����3@�߆�s�!?M�r04|�@eD����ٿ;o�OC�@KHa;��3@��X�!?�����@��.�ٿ�"�*��@d�s���3@��d�!?>|�4�@��.�ٿ�"�*��@d�s���3@��d�!?>|�4�@��.�ٿ�"�*��@d�s���3@��d�!?>|�4�@��.�ٿ�"�*��@d�s���3@��d�!?>|�4�@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@:_����ٿ��v'�@}���k�3@��a:�!?>�-��@�mw3��ٿD��m�@��S�x�3@�I
��!?��C?Q��@�mw3��ٿD��m�@��S�x�3@�I
��!?��C?Q��@�mw3��ٿD��m�@��S�x�3@�I
��!?��C?Q��@�mw3��ٿD��m�@��S�x�3@�I
��!?��C?Q��@B=��<�ٿ]��z�w�@�y�So�3@h��b�!?N��;�ô@B=��<�ٿ]��z�w�@�y�So�3@h��b�!?N��;�ô@B=��<�ٿ]��z�w�@�y�So�3@h��b�!?N��;�ô@B=��<�ٿ]��z�w�@�y�So�3@h��b�!?N��;�ô@�;L�S�ٿ�'ҿ܂�@H�
��3@��z[=�!?��^��@�;L�S�ٿ�'ҿ܂�@H�
��3@��z[=�!?��^��@�;L�S�ٿ�'ҿ܂�@H�
��3@��z[=�!?��^��@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@.D�U�ٿ���i�@���ɖ�3@�CߜY�!?�@�(R�@��I�h�ٿ������@q� ,�3@�KA�U�!?�**Y�@��I�h�ٿ������@q� ,�3@�KA�U�!?�**Y�@��I�h�ٿ������@q� ,�3@�KA�U�!?�**Y�@��I�h�ٿ������@q� ,�3@�KA�U�!?�**Y�@��I�h�ٿ������@q� ,�3@�KA�U�!?�**Y�@��J�ٿۨ3����@\����3@�ǲmi�!?�ޥM.2�@��J�ٿۨ3����@\����3@�ǲmi�!?�ޥM.2�@��J�ٿۨ3����@\����3@�ǲmi�!?�ޥM.2�@����ٿ�
��+M�@��.b��3@D#s1O�!?+ɑ�5�@��вg�ٿ2��`��@��7��3@���!?g�W�[�@��вg�ٿ2��`��@��7��3@���!?g�W�[�@_�����ٿ����V�@��R��3@����E�!?�����@R!yX��ٿ��$W�@ȡ)uW�3@Q�Gg�!?8��u1�@R!yX��ٿ��$W�@ȡ)uW�3@Q�Gg�!?8��u1�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@^ޖ��ٿ��#����@�c����3@c���P�!?�Z���R�@�?��ٿ�77���@Z� � 4@Y>M5d�!?�����@�_n�ٿ=�lמ{�@��dś�3@Z7޴%�!?n��	4ص@m�÷�ٿ�+�&��@ȍEn��3@^5ڤi�!?w`�J�@m�÷�ٿ�+�&��@ȍEn��3@^5ڤi�!?w`�J�@m�÷�ٿ�+�&��@ȍEn��3@^5ڤi�!?w`�J�@�]t�ݙٿ��	d[�@������3@�6�h�!?����Eq�@�]t�ݙٿ��	d[�@������3@�6�h�!?����Eq�@�]t�ݙٿ��	d[�@������3@�6�h�!?����Eq�@�]t�ݙٿ��	d[�@������3@�6�h�!?����Eq�@�]t�ݙٿ��	d[�@������3@�6�h�!?����Eq�@(a��C�ٿ��Z�|�@Ǹ�|~�3@���l\�!?H)tQ��@(a��C�ٿ��Z�|�@Ǹ�|~�3@���l\�!?H)tQ��@(a��C�ٿ��Z�|�@Ǹ�|~�3@���l\�!?H)tQ��@(a��C�ٿ��Z�|�@Ǹ�|~�3@���l\�!?H)tQ��@(a��C�ٿ��Z�|�@Ǹ�|~�3@���l\�!?H)tQ��@#�@ "�ٿi�*�w�@N{���3@ܬ�p�!?{|(c��@#�@ "�ٿi�*�w�@N{���3@ܬ�p�!?{|(c��@2���f�ٿ���r�@��v<J�3@YQӰx�!?��[Q�@2���f�ٿ���r�@��v<J�3@YQӰx�!?��[Q�@2���f�ٿ���r�@��v<J�3@YQӰx�!?��[Q�@���*J�ٿ�=�=W�@(�s��3@�+"�Q�!?�I�kI+�@���*J�ٿ�=�=W�@(�s��3@�+"�Q�!?�I�kI+�@Gz��ٿ����&�@������3@����;�!?I�_PJ�@�B�f��ٿ��Z�H�@W+�k4�3@�Z��!?~���~�@�O6z�ٿ���l3�@��M�W�3@����T�!?�By�T�@�a���ٿ�����n�@a�5�3@�G�*�!?�8U|'��@�a���ٿ�����n�@a�5�3@�G�*�!?�8U|'��@�a���ٿ�����n�@a�5�3@�G�*�!?�8U|'��@�a���ٿ�����n�@a�5�3@�G�*�!?�8U|'��@V��>G�ٿ�����@��h�3@��e�x�!?��ݼ��@V��>G�ٿ�����@��h�3@��e�x�!?��ݼ��@)�2�o�ٿ]3��?��@�W����3@�+�j�!?��]�Ю�@)�2�o�ٿ]3��?��@�W����3@�+�j�!?��]�Ю�@)�2�o�ٿ]3��?��@�W����3@�+�j�!?��]�Ю�@)�2�o�ٿ]3��?��@�W����3@�+�j�!?��]�Ю�@)�2�o�ٿ]3��?��@�W����3@�+�j�!?��]�Ю�@��
�ٿ[x-����@����6�3@L ��W�!?��bv�@��
�ٿ[x-����@����6�3@L ��W�!?��bv�@1B}���ٿ{���� �@b�K. �3@I!M�=�!?
.xȅ�@����ٿQka\��@���)$�3@��jA#�!?��dml�@����ٿQka\��@���)$�3@��jA#�!?��dml�@����ٿQka\��@���)$�3@��jA#�!?��dml�@����ٿQka\��@���)$�3@��jA#�!?��dml�@w�+�ٿ�������@i�aY��3@
�@�I�!?ʶ �/��@GNFX�ٿ����@J����3@��B!?�Tl��c�@GNFX�ٿ����@J����3@��B!?�Tl��c�@GNFX�ٿ����@J����3@��B!?�Tl��c�@GNFX�ٿ����@J����3@��B!?�Tl��c�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@�v�/�ٿ-�����@�ɜ�\�3@��z�!?��Y��]�@%l$�S�ٿ�n���@Xކ��3@��"�a�!?0���1�@c�d�ٿ5�X�K��@ɇm��3@���-�!?�d�.��@c�d�ٿ5�X�K��@ɇm��3@���-�!?�d�.��@c�d�ٿ5�X�K��@ɇm��3@���-�!?�d�.��@!��j�ٿ-P~�à�@�RlX��3@ϸ%��!?��v�+��@!��j�ٿ-P~�à�@�RlX��3@ϸ%��!?��v�+��@�W����ٿ+r���?�@��\*�3@�F�!?,7�ZxԵ@�W����ٿ+r���?�@��\*�3@�F�!?,7�ZxԵ@�W����ٿ+r���?�@��\*�3@�F�!?,7�ZxԵ@�W����ٿ+r���?�@��\*�3@�F�!?,7�ZxԵ@����ٿTNt�!�@K{`:/�3@.F�yJ�!?��[�o��@��B-՞ٿ��[���@xs��3@<�08�!?dC��z��@��B-՞ٿ��[���@xs��3@<�08�!?dC��z��@��B-՞ٿ��[���@xs��3@<�08�!?dC��z��@ʌ����ٿ��MK�v�@dˀ�
�3@���@�!?U�tiZ�@ʌ����ٿ��MK�v�@dˀ�
�3@���@�!?U�tiZ�@���G:�ٿ�/��f��@C����3@�g	��!?G�Zϵ@�M�י�ٿH� ���@�����3@C$p�!?�������@�M�י�ٿH� ���@�����3@C$p�!?�������@�M�י�ٿH� ���@�����3@C$p�!?�������@ڣ�Tq�ٿ�48��@������3@+���!?vb9�jW�@ڣ�Tq�ٿ�48��@������3@+���!?vb9�jW�@ڣ�Tq�ٿ�48��@������3@+���!?vb9�jW�@ڣ�Tq�ٿ�48��@������3@+���!?vb9�jW�@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�� ��ٿ���
��@_V��o�3@1*=L~�!?ǢO��@�?�!�ٿ kLm���@��"?D�3@t���{�!?2²�I��@�?�!�ٿ kLm���@��"?D�3@t���{�!?2²�I��@�?�!�ٿ kLm���@��"?D�3@t���{�!?2²�I��@�C�ؚٿ�^ ���@��I��3@��I���!?
�`kq;�@�C�ؚٿ�^ ���@��I��3@��I���!?
�`kq;�@�C�ؚٿ�^ ���@��I��3@��I���!?
�`kq;�@�4漘ٿ��m��@�]��3@΅`;�!?�N)<���@�4漘ٿ��m��@�]��3@΅`;�!?�N)<���@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@�5�d�ٿ��̧���@W��&��3@?.��9�!?
�sQ�,�@Ի�V�ٿ���UD��@-/2Y�3@�h��s�!?t���Q�@Ի�V�ٿ���UD��@-/2Y�3@�h��s�!?t���Q�@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@$�b��ٿ�����@<��S�3@m,P��!?8 ����@�1�|��ٿ��7��k�@���y�3@�{_�!?�hȏ4h�@���0גٿ�X�,)E�@��@�� 4@[1��!?�a詍��@���0גٿ�X�,)E�@��@�� 4@[1��!?�a詍��@�?����ٿN@�^��@��M� 4@����!?�w� ߐ�@�?����ٿN@�^��@��M� 4@����!?�w� ߐ�@uB��ٿ�M�̲�@ڄ�
�3@���|��!?�zMW�@uB��ٿ�M�̲�@ڄ�
�3@���|��!?�zMW�@uB��ٿ�M�̲�@ڄ�
�3@���|��!?�zMW�@;`�Q˔ٿl���h`�@�>d��3@����f�!?D{!.W��@;`�Q˔ٿl���h`�@�>d��3@����f�!?D{!.W��@;`�Q˔ٿl���h`�@�>d��3@����f�!?D{!.W��@�e-=�ٿ�(��&�@���J��3@ő���!?�V�ϵ@�e-=�ٿ�(��&�@���J��3@ő���!?�V�ϵ@�e-=�ٿ�(��&�@���J��3@ő���!?�V�ϵ@m�g ��ٿ'#�`�@����E�3@o�|�ڏ!?�&O2y��@�A~�T�ٿq�Ū!�@6�G��3@�����!?FP��n�@�A~�T�ٿq�Ū!�@6�G��3@�����!?FP��n�@�A~�T�ٿq�Ū!�@6�G��3@�����!?FP��n�@�A~�T�ٿq�Ū!�@6�G��3@�����!?FP��n�@�A~�T�ٿq�Ū!�@6�G��3@�����!?FP��n�@[j4牒ٿi@�
�@�<�)�3@��� �!?����h�@'j7,��ٿO�s���@����1�3@��	��!?8b%G��@'j7,��ٿO�s���@����1�3@��	��!?8b%G��@'j7,��ٿO�s���@����1�3@��	��!?8b%G��@=A���ٿ&�}� �@9�vJM�3@�R�?ۏ!?�`���@=A���ٿ&�}� �@9�vJM�3@�R�?ۏ!?�`���@=A���ٿ&�}� �@9�vJM�3@�R�?ۏ!?�`���@=A���ٿ&�}� �@9�vJM�3@�R�?ۏ!?�`���@֭�٧�ٿC�`�w�@3��i/	4@UD�O�!?��YӼ�@:Q)���ٿ��NO�@��dv	4@���>�!?���u�@�����ٿ���z���@Tg�$g4@��%�!?��{��T�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@�G�	̖ٿ�A�q�}�@����4@��x�S�!?�QL+�1�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@���o��ٿ�|�a�@<O��4@���e�!?�a4^�@�1!L=�ٿ��Ђ6��@mH�i�3@�e�!?������@�1!L=�ٿ��Ђ6��@mH�i�3@�e�!?������@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���e�ٿ�[�'��@�O��U�3@ 2��F�!?��UF�@���ƒٿ%�#�N��@�-����3@��v�!?K.G���@܄;^y�ٿp�NG]�@w���3@�f��Ȑ!?�f%�%�@܄;^y�ٿp�NG]�@w���3@�f��Ȑ!?�f%�%�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@�����ٿǫ"e�@B�bmJ�3@a8�=�!?�7��,�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@��F.��ٿBüȀ��@R��`��3@؍�F�!?�D �`�@�"�ٿ	M>4���@�%ޭ(�3@���O�!?VE{�O�@�"�ٿ	M>4���@�%ޭ(�3@���O�!?VE{�O�@�����ٿ�h���r�@:(�@�3@��(B�!?��#��Ǵ@a�v�t�ٿ�"D�	~�@�G����3@��B,�!?�+4;��@a�v�t�ٿ�"D�	~�@�G����3@��B,�!?�+4;��@D0\uk�ٿ��0H��@@\H�3@�|��%�!?(�SG�L�@Oۗ
8�ٿZxҽ�@b��"�3@n��t�!?�.�"�j�@Oۗ
8�ٿZxҽ�@b��"�3@n��t�!?�.�"�j�@By�g��ٿ��O�͵�@��ߣf�3@5@�G�!?(�\�� �@By�g��ٿ��O�͵�@��ߣf�3@5@�G�!?(�\�� �@.J1v��ٿ���m��@�4x���3@`���!?�J��썴@.J1v��ٿ���m��@�4x���3@`���!?�J��썴@.J1v��ٿ���m��@�4x���3@`���!?�J��썴@.J1v��ٿ���m��@�4x���3@`���!?�J��썴@[a���ٿ�{8�@¼����3@f��}$�!?�'��x2�@[a���ٿ�{8�@¼����3@f��}$�!?�'��x2�@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@88Y���ٿ�ܛ��@>�T��3@�Q-��!?rY����@�Y'�Ҕٿ	�H�c�@-pf��3@rlt%�!?�1��y�@�Y'�Ҕٿ	�H�c�@-pf��3@rlt%�!?�1��y�@�Y'�Ҕٿ	�H�c�@-pf��3@rlt%�!?�1��y�@�Y'�Ҕٿ	�H�c�@-pf��3@rlt%�!?�1��y�@�Y'�Ҕٿ	�H�c�@-pf��3@rlt%�!?�1��y�@>��*�ٿV��vx��@��E0+4@�ly	K�!? ����@>��*�ٿV��vx��@��E0+4@�ly	K�!? ����@>��*�ٿV��vx��@��E0+4@�ly	K�!? ����@>��*�ٿV��vx��@��E0+4@�ly	K�!? ����@�c���ٿ�6|Ӈ:�@$?���3@�|a{�!?`�@�,���ٿ$�����@n3�~�3@���r�!?;�$��@���Z�ٿ2�h����@�9 &�3@�.,6��!?�]��r�@���Z�ٿ2�h����@�9 &�3@�.,6��!?�]��r�@���Z�ٿ2�h����@�9 &�3@�.,6��!?�]��r�@�����ٿ�D䴩�@�Y(S��3@��@~�!?�0͓�@�����ٿ�D䴩�@�Y(S��3@��@~�!?�0͓�@�����ٿ�D䴩�@�Y(S��3@��@~�!?�0͓�@T�WC�ٿ�T-��@����3@�!v5�!?�߈R0��@T�WC�ٿ�T-��@����3@�!v5�!?�߈R0��@d�ce!�ٿ����@ k�)�3@Y����!?/V9�A3�@d�ce!�ٿ����@ k�)�3@Y����!?/V9�A3�@d�ce!�ٿ����@ k�)�3@Y����!?/V9�A3�@d�ce!�ٿ����@ k�)�3@Y����!?/V9�A3�@d�ce!�ٿ����@ k�)�3@Y����!?/V9�A3�@wQ�)��ٿѫ����@u]���4@%Q�!?�Vl�b�@��.k��ٿ��Ņ��@眽ޅ�3@(��!?sP�܌J�@��.k��ٿ��Ņ��@眽ޅ�3@(��!?sP�܌J�@0t���ٿ��ԴY��@$�����3@�9.a�!?f��:k�@0t���ٿ��ԴY��@$�����3@�9.a�!?f��:k�@0t���ٿ��ԴY��@$�����3@�9.a�!?f��:k�@����<�ٿa�'���@f�3,A4@�:�5:�!?�����r�@����6�ٿ�$�^9�@|ڑ�j�3@�uU��!?��-�(�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@0[��ٿ�[Mo׽�@�Q���3@�u�`�!?Q>�c�@��8�a�ٿ�h����@l�����3@짺Ј�!?����gg�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@�F�Aq�ٿ���]���@M=p�O�3@�S�[��!?g�JTi�@����ٿt���@��Jj8�3@1&=.Ő!?b�x#��@����ٿt���@��Jj8�3@1&=.Ő!?b�x#��@^\��
�ٿ�<2`��@��?��3@S�Iq��!?.�����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@��͌�ٿ8��j��@2�l��3@<YEä�!?Dm
����@�T��1�ٿ V�����@]�Y���3@�oTK�!?Grs&�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@s>�Oڛٿ����]�@�u�x4@>6��A�!?��{@�@jc'���ٿ2c:B��@Z�Ay4@fUI�!?!���_�@jc'���ٿ2c:B��@Z�Ay4@fUI�!?!���_�@jc'���ٿ2c:B��@Z�Ay4@fUI�!?!���_�@�Q~��ٿ��j�0�@t(_��4@qhv�G�!?�NS<��@�Q~��ٿ��j�0�@t(_��4@qhv�G�!?�NS<��@�Q~��ٿ��j�0�@t(_��4@qhv�G�!?�NS<��@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�t��e�ٿ�"�}]k�@���
�3@c,升�!?�z���-�@�wQ��ٿ�٩4���@�
&�W�3@T`k�z�!?c��ֵ�@�wQ��ٿ�٩4���@�
&�W�3@T`k�z�!?c��ֵ�@�wQ��ٿ�٩4���@�
&�W�3@T`k�z�!?c��ֵ�@�o�4��ٿXh����@��:L��3@�����!?�Qf\y�@�o�4��ٿXh����@��:L��3@�����!?�Qf\y�@}5l�Y�ٿ���I*�@*�q���3@L�dJ�!?ybn���@}5l�Y�ٿ���I*�@*�q���3@L�dJ�!?ybn���@}5l�Y�ٿ���I*�@*�q���3@L�dJ�!?ybn���@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�u^��ٿ7�5'd�@[w�63�3@�?4i�!?�.�}�\�@�����ٿ���ޝ��@�,�&4@�b����!?���O�@�����ٿ���ޝ��@�,�&4@�b����!?���O�@�����ٿ���ޝ��@�,�&4@�b����!?���O�@�����ٿ���ޝ��@�,�&4@�b����!?���O�@�����ٿ���ޝ��@�,�&4@�b����!?���O�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@_�[���ٿؠbXK>�@7�a�i�3@��̟��!?�X9��j�@��̭&�ٿL����@�>'�3@kd|J�!?��b|�@��̭&�ٿL����@�>'�3@kd|J�!?��b|�@��̭&�ٿL����@�>'�3@kd|J�!?��b|�@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@se���ٿ��=8S�@�@����3@.���!?H���δ@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@<�����ٿ����-�@�]D��3@�ĕ�(�!?���%�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@)1��a�ٿ��s:�b�@HDv���3@b[?gn�!?��5�@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@a�9���ٿ��~,�@�p��]�3@b��)Z�!?�5�#��@�-|%�ٿ�W�Y��@t����3@��av�!?/�R״@�-|%�ٿ�W�Y��@t����3@��av�!?/�R״@�-|%�ٿ�W�Y��@t����3@��av�!?/�R״@�?ݧ�ٿ���a}��@�B���3@or��?�!?Cs�p�5�@�?ݧ�ٿ���a}��@�B���3@or��?�!?Cs�p�5�@T��a��ٿ���I��@�0�<��3@�BaOZ�!?�)q5�r�@�D���ٿ0����@~d0j�3@�>8�f�!? k��@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@�jt�d�ٿFfh���@f���3@��吐!?
&�3�@��E�ٿ�QzISO�@K>$��3@+���!?� �o�@���ٿ����B�@◇���3@2�* �!?w�r��@���ٿ����B�@◇���3@2�* �!?w�r��@���ٿ����B�@◇���3@2�* �!?w�r��@���ٿ����B�@◇���3@2�* �!?w�r��@!p�$��ٿ�|�:S�@���p�3@�`�쥐!?�u;�Xe�@!p�$��ٿ�|�:S�@���p�3@�`�쥐!?�u;�Xe�@!p�$��ٿ�|�:S�@���p�3@�`�쥐!?�u;�Xe�@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@�q���ٿ�����@o���3@μ����!?x�Z䖴@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��N�i�ٿ��	�@�$�d��3@{���А!?"���ˇ�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@��u�ٿ��ֵ)��@W"�_��3@��j�2�!?'4u��+�@���Ǚٿ�)� >h�@��]��3@��~�!?���>u�@���Ǚٿ�)� >h�@��]��3@��~�!?���>u�@���Ǚٿ�)� >h�@��]��3@��~�!?���>u�@���Ǚٿ�)� >h�@��]��3@��~�!?���>u�@k����ٿ6��8���@��1s�3@d	��M�!?�v�a�Ӵ@s��ٿx��_ �@�/x��3@!L.`�!?���ت��@���T�ٿ!+��!��@El=	�3@�0\F��!?�&��m~�@���T�ٿ!+��!��@El=	�3@�0\F��!?�&��m~�@���T�ٿ!+��!��@El=	�3@�0\F��!?�&��m~�@���T�ٿ!+��!��@El=	�3@�0\F��!?�&��m~�@BM�+��ٿ��Q
��@���V�3@���ˢ�!? ��y��@BM�+��ٿ��Q
��@���V�3@���ˢ�!? ��y��@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�ڮ�3�ٿᰲ���@�Z��n�3@!z�Er�!?�R��t�@�D�x1�ٿ�Q�0��@�UW��3@�=�ゐ!?#8ac�@�D�x1�ٿ�Q�0��@�UW��3@�=�ゐ!?#8ac�@�D�x1�ٿ�Q�0��@�UW��3@�=�ゐ!?#8ac�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@,7�@'�ٿy��NQ�@N��F�3@�c�*~�!?9��R�@&�K�ٿ)!c]��@��Y�3@g_��Y�!?$�����@�Ų���ٿ,����@��=���3@��'�B�!?��R�!��@�u�x�ٿ3<?����@#��M%4@��4�!?:d,ީ�@]�#��ٿ����T�@߯���3@y�*܍�!?�ȇ4z��@]�#��ٿ����T�@߯���3@y�*܍�!?�ȇ4z��@]�#��ٿ����T�@߯���3@y�*܍�!?�ȇ4z��@]�#��ٿ����T�@߯���3@y�*܍�!?�ȇ4z��@LWƣԕٿ��Y��(�@cz�+��3@��L��!?,��Ǫ��@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@�ߛ���ٿ����m�@܃ʹ$�3@r�!?4���'�@+��iӑٿx�?h���@m��8��3@�U�`{�!?���uo��@��x�ٿ���}*�@�m'L��3@����!?"��7~��@��x�ٿ���}*�@�m'L��3@����!?"��7~��@��x�ٿ���}*�@�m'L��3@����!?"��7~��@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@W�?�9�ٿ*NOi��@��Z�3@R�3g�!?[�Ђ͵@�	��ٿ@�,9+^�@	g,��3@e��{�!?2"��P%�@�	��ٿ@�,9+^�@	g,��3@e��{�!?2"��P%�@�	��ٿ@�,9+^�@	g,��3@e��{�!?2"��P%�@+�&�/�ٿ�3����@KU�v�3@r�g�
�!?�z��#��@+�&�/�ٿ�3����@KU�v�3@r�g�
�!?�z��#��@�*�n�ٿ���>��@>�B��3@��EA'�!?ӟ`  ��@F�I�Аٿ��dݵ��@����Y4@#�5/�!?�2�=-�@F�I�Аٿ��dݵ��@����Y4@#�5/�!?�2�=-�@F�I�Аٿ��dݵ��@����Y4@#�5/�!?�2�=-�@�� ��ٿ������@� J�$�3@Z~涏!?)7��*��@�� ��ٿ������@� J�$�3@Z~涏!?)7��*��@h�x�)�ٿ��#@-[�@%��k�3@8���!?6v�;���@h�x�)�ٿ��#@-[�@%��k�3@8���!?6v�;���@h�x�)�ٿ��#@-[�@%��k�3@8���!?6v�;���@h�x�)�ٿ��#@-[�@%��k�3@8���!?6v�;���@���܈�ٿ^��*�@oVY�y�3@��?��!?9���Ҵ@���܈�ٿ^��*�@oVY�y�3@��?��!?9���Ҵ@���܈�ٿ^��*�@oVY�y�3@��?��!?9���Ҵ@�dn��ٿ=��E��@&H\��3@}_$��!?2	>�Z�@�dn��ٿ=��E��@&H\��3@}_$��!?2	>�Z�@�dn��ٿ=��E��@&H\��3@}_$��!?2	>�Z�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@0q%ƌ�ٿ9f|����@�|۱�3@�6���!?C*qSS�@���E�ٿ1���@���"��3@��<!?A��U��@���E�ٿ1���@���"��3@��<!?A��U��@���E�ٿ1���@���"��3@��<!?A��U��@���E�ٿ1���@���"��3@��<!?A��U��@b '��ٿ���^�"�@�x�_��3@��I��!?
��+��@b '��ٿ���^�"�@�x�_��3@��I��!?
��+��@b '��ٿ���^�"�@�x�_��3@��I��!?
��+��@b '��ٿ���^�"�@�x�_��3@��I��!?
��+��@��!���ٿ�1���*�@E����3@���͏!?[-�;�@��!���ٿ�1���*�@E����3@���͏!?[-�;�@;%�V��ٿ5�x��@�+�W_�3@�-�*n�!?��n3G�@;%�V��ٿ5�x��@�+�W_�3@�-�*n�!?��n3G�@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@N�+q�ٿ).8d3��@�3_�9�3@6f/Ψ�!?u8�4�ɴ@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�,��ٿ�����@�ȍ��3@F�;qF�!?O%8J���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@�@��ٿQ��a
�@K�x̳�3@v�R��!?C�j���@��U���ٿש;�&��@�-TR%�3@�e6/�!?�k�O��@��U���ٿש;�&��@�-TR%�3@�e6/�!?�k�O��@��U���ٿש;�&��@�-TR%�3@�e6/�!?�k�O��@�}�γ�ٿ
X�P�@˂�D��3@Z�KL�!?��&��6�@�}�γ�ٿ
X�P�@˂�D��3@Z�KL�!?��&��6�@�}�γ�ٿ
X�P�@˂�D��3@Z�KL�!?��&��6�@�}�γ�ٿ
X�P�@˂�D��3@Z�KL�!?��&��6�@�}�γ�ٿ
X�P�@˂�D��3@Z�KL�!?��&��6�@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@�N�Z*�ٿ �ـ���@���3@�Waj6�!?oF����@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@��_�ٿ$Ɓ�U�@X%���3@��n�!?6�"�*�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@D�4���ٿ�P���a�@ߢ4�:�3@N����!?����S�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@L�ؠ��ٿb;0ŉX�@DsD���3@^��7�!?T�m��x�@Q�:�ٿ�l�~�@\h�:�4@�T	�!? ��)dK�@Q�:�ٿ�l�~�@\h�:�4@�T	�!? ��)dK�@Q�:�ٿ�l�~�@\h�:�4@�T	�!? ��)dK�@Q�:�ٿ�l�~�@\h�:�4@�T	�!? ��)dK�@Q�:�ٿ�l�~�@\h�:�4@�T	�!? ��)dK�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@Ӗ�$�ٿ=������@�I4@	���1�!?Z�!Ns*�@PWӡ�ٿg$Y�u�@̃$e
4@1��^a�!?��ǽ��@PWӡ�ٿg$Y�u�@̃$e
4@1��^a�!?��ǽ��@PWӡ�ٿg$Y�u�@̃$e
4@1��^a�!?��ǽ��@PWӡ�ٿg$Y�u�@̃$e
4@1��^a�!?��ǽ��@x ��a�ٿZ�6jn�@�0����3@`3n��!?��3�@x ��a�ٿZ�6jn�@�0����3@`3n��!?��3�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@�����ٿ�ރ��@�h���3@�0,��!?�!2�ބ�@i\C���ٿ2�Q��@�X����3@�H%�!?eB�����@i\C���ٿ2�Q��@�X����3@�H%�!?eB�����@i\C���ٿ2�Q��@�X����3@�H%�!?eB�����@i\C���ٿ2�Q��@�X����3@�H%�!?eB�����@��u���ٿg�z3�@���tr�3@��^)�!?Q�kˣ�@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@�!� �ٿ��-�{�@{28��3@��r�!?&�,@��@��W��ٿ�5��0��@��pw�3@P3/��!?����H�@��W��ٿ�5��0��@��pw�3@P3/��!?����H�@��W��ٿ�5��0��@��pw�3@P3/��!?����H�@��W��ٿ�5��0��@��pw�3@P3/��!?����H�@��LϜٿA���&��@�4�~��3@X�✐!?�H����@��LϜٿA���&��@�4�~��3@X�✐!?�H����@��LϜٿA���&��@�4�~��3@X�✐!?�H����@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@N|Xɜ�ٿ�N���@Q���3@�O?�/�!?1L�V�w�@Gu��m�ٿ���\�@h����3@ h8�!?�3f뿪�@Gu��m�ٿ���\�@h����3@ h8�!?�3f뿪�@Gu��m�ٿ���\�@h����3@ h8�!?�3f뿪�@Gu��m�ٿ���\�@h����3@ h8�!?�3f뿪�@Gu��m�ٿ���\�@h����3@ h8�!?�3f뿪�@�1U�_�ٿ�W#Q�@pi9��3@ߜ�I5�!?��d��@�1U�_�ٿ�W#Q�@pi9��3@ߜ�I5�!?��d��@�1U�_�ٿ�W#Q�@pi9��3@ߜ�I5�!?��d��@����'�ٿ�wY&!��@�wA���3@G�L��!?��8#"�@����'�ٿ�wY&!��@�wA���3@G�L��!?��8#"�@��9�ϒٿ��T�!�@7ZK��3@�ڤ�E�!?~f����@��9�ϒٿ��T�!�@7ZK��3@�ڤ�E�!?~f����@��9�ϒٿ��T�!�@7ZK��3@�ڤ�E�!?~f����@��9�ϒٿ��T�!�@7ZK��3@�ڤ�E�!?~f����@���^Ԓٿ+0��=��@���+�3@�w6���!?W��LҴ@���^Ԓٿ+0��=��@���+�3@�w6���!?W��LҴ@���^Ԓٿ+0��=��@���+�3@�w6���!?W��LҴ@���^Ԓٿ+0��=��@���+�3@�w6���!?W��LҴ@���^Ԓٿ+0��=��@���+�3@�w6���!?W��LҴ@5f��5�ٿG��N�@�<R|[�3@�|�ȥ�!?z�ӂ�״@5f��5�ٿG��N�@�<R|[�3@�|�ȥ�!?z�ӂ�״@�Z�v�ٿf����=�@����o�3@K�l���!?��P�c7�@�Xֵ�ٿYCHl}��@�&,\U4@��
~{�!?C��`V��@�Xֵ�ٿYCHl}��@�&,\U4@��
~{�!?C��`V��@��R��ٿ����W�@�+k3�4@�KVa�!?���Ƶ@��R��ٿ����W�@�+k3�4@�KVa�!?���Ƶ@��R��ٿ����W�@�+k3�4@�KVa�!?���Ƶ@��R��ٿ����W�@�+k3�4@�KVa�!?���Ƶ@��R��ٿ����W�@�+k3�4@�KVa�!?���Ƶ@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@�4�Ŗٿ���>��@
�D��3@腿k�!?��o�U�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@��`�F�ٿf�	�$��@�Xy� �3@wE!�>�!?'�Nr7i�@eᏧ,�ٿ+O�^)�@�f8��3@��T囐!?��� �@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@�`+Ԭ�ٿ���3��@w֑)Y�3@@Q��_�!?e��[�H�@��~�ٿzz�T<�@�Q�O�3@�]>��!?��IfL�@���ٿ֡+%y�@vU(��3@O�(��!?��#�?�@S����ٿIue��'�@������3@��lܛ�!?�gk�L:�@S����ٿIue��'�@������3@��lܛ�!?�gk�L:�@S����ٿIue��'�@������3@��lܛ�!?�gk�L:�@S����ٿIue��'�@������3@��lܛ�!?�gk�L:�@�B�іٿ{f��L�@�3��3@�G	\]�!?��cL96�@�B�іٿ{f��L�@�3��3@�G	\]�!?��cL96�@sӷ�H�ٿs{�'��@C��s�3@��^_�!?�Z+b�@sӷ�H�ٿs{�'��@C��s�3@��^_�!?�Z+b�@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@k�M��ٿ�1(��G�@*����3@��ջ�!?����@�
`�'�ٿ*I�{:.�@�@Һa�3@��)��!?X�nX��@�
`�'�ٿ*I�{:.�@�@Һa�3@��)��!?X�nX��@�
`�'�ٿ*I�{:.�@�@Һa�3@��)��!?X�nX��@�
`�'�ٿ*I�{:.�@�@Һa�3@��)��!?X�nX��@�
`�'�ٿ*I�{:.�@�@Һa�3@��)��!?X�nX��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@2��#��ٿPڞ����@�&����3@�=o��!?�ޠ��@ ���^�ٿ�Z,j1�@��sN�3@^Y��!?j��Qv�@��q�<�ٿ|L���;�@�V�8�3@K4|�]�!?c��(1��@��q�<�ٿ|L���;�@�V�8�3@K4|�]�!?c��(1��@���(�ٿh�����@8�ۓc4@���0��!?���Q3�@���(�ٿh�����@8�ۓc4@���0��!?���Q3�@�9�ᮓٿ�k&G�|�@����b�3@08�oY�!?����\�@�p���ٿV�V���@͆�Q�3@�}�H�!?�!t=�@�p���ٿV�V���@͆�Q�3@�}�H�!?�!t=�@�p���ٿV�V���@͆�Q�3@�}�H�!?�!t=�@�p���ٿV�V���@͆�Q�3@�}�H�!?�!t=�@�p���ٿV�V���@͆�Q�3@�}�H�!?�!t=�@t�2��ٿWd?�N��@��n���3@���:�!?/j���o�@t�2��ٿWd?�N��@��n���3@���:�!?/j���o�@t�2��ٿWd?�N��@��n���3@���:�!?/j���o�@*%	�7�ٿ�`��t�@EB1P��3@K���/�!?��C3��@��f��ٿN���.�@$U���3@`���%�!?5lwK��@��f��ٿN���.�@$U���3@`���%�!?5lwK��@"��M�ٿ�����@��K�3@���L�!?�5s�/�@"��M�ٿ�����@��K�3@���L�!?�5s�/�@<���O�ٿk�#_L�@�(���3@���b�!?�Su$@�@<���O�ٿk�#_L�@�(���3@���b�!?�Su$@�@�t�b@�ٿE20
���@������3@"E���!?��sJ! �@�t�b@�ٿE20
���@������3@"E���!?��sJ! �@�t�b@�ٿE20
���@������3@"E���!?��sJ! �@3Y�V�ٿ���|�@�ϡz�3@��-Ԑ!?Tr�;#6�@3Y�V�ٿ���|�@�ϡz�3@��-Ԑ!?Tr�;#6�@�
��a�ٿ]w�L�@���k�3@6ɐ!?�ȮoѴ@7��B�ٿ�M�\D.�@Z�$"�3@G��K�!?q�A�G�@7��B�ٿ�M�\D.�@Z�$"�3@G��K�!?q�A�G�@��+�S�ٿ�m�3W�@P��S�3@�IB.�!?��P�n�@��+�S�ٿ�m�3W�@P��S�3@�IB.�!?��P�n�@V{՘N�ٿ���W�X�@�*\�3@(�e̋�!?�n��}�@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@()I�ٿ�����@vw��)4@��O�{�!?b��JZ��@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@���[�ٿ.�C�@�C�[n�3@ZE&��!?��[�ڴ@�{�l�ٿs�7���@ｐ�\�3@<_됐!?������@�{�l�ٿs�7���@ｐ�\�3@<_됐!?������@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@9E�J/�ٿ\��(�@�]Z���3@��u�3�!?�)���@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@�~�j��ٿ �l{w��@c%�E�3@�,��}�!?�����@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@wn�"ɒٿ�Ӯg*�@�?�O�3@�,J�`�!?s�pGM�@l]�Q�ٿ�T
:��@</:���3@��k��!?����婴@l]�Q�ٿ�T
:��@</:���3@��k��!?����婴@l]�Q�ٿ�T
:��@</:���3@��k��!?����婴@l]�Q�ٿ�T
:��@</:���3@��k��!?����婴@l]�Q�ٿ�T
:��@</:���3@��k��!?����婴@9cK��ٿ�h�}g��@K4��9�3@��ӥ-�!?=�+ܤ�@9cK��ٿ�h�}g��@K4��9�3@��ӥ-�!?=�+ܤ�@9cK��ٿ�h�}g��@K4��9�3@��ӥ-�!?=�+ܤ�@Z�2��ٿ�%�a��@J����3@Հ/[	�!?��|�U�@Z�2��ٿ�%�a��@J����3@Հ/[	�!?��|�U�@Z�2��ٿ�%�a��@J����3@Հ/[	�!?��|�U�@Z�2��ٿ�%�a��@J����3@Հ/[	�!?��|�U�@,�n��ٿ�!{)E�@��Cb�3@-��%�!?��YtM�@�:�u�ٿg<%r��@x���3@�j��!?�m�Ѝڴ@�:�u�ٿg<%r��@x���3@�j��!?�m�Ѝڴ@�:�u�ٿg<%r��@x���3@�j��!?�m�Ѝڴ@/D@�ٿ�Q��V*�@��y�3@��K+%�!?RI�O���@/D@�ٿ�Q��V*�@��y�3@��K+%�!?RI�O���@/D@�ٿ�Q��V*�@��y�3@��K+%�!?RI�O���@�=�q�ٿ8���m��@�*r�@�3@�Y���!?U���@��@�=�q�ٿ8���m��@�*r�@�3@�Y���!?U���@��@�=�q�ٿ8���m��@�*r�@�3@�Y���!?U���@��@��1p&�ٿ��p����@�(-V��3@w�e{g�!?:��r�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@�	󅏚ٿ"�QA�M�@����R�3@�八N�!?z���	F�@���nٿ��'6L�@���$��3@ �aoN�!?y�0��@���nٿ��'6L�@���$��3@ �aoN�!?y�0��@on��>�ٿrj�^�@���_�3@H����!?p���G�@on��>�ٿrj�^�@���_�3@H����!?p���G�@�ҷ��ٿ���h��@2�ԋ 4@���M$�!?{�4O.��@�ҷ��ٿ���h��@2�ԋ 4@���M$�!?{�4O.��@�ҷ��ٿ���h��@2�ԋ 4@���M$�!?{�4O.��@����ٿ�#��D�@�����4@Y���i�!?��hzl�@����ٿ�#��D�@�����4@Y���i�!?��hzl�@����ٿ�#��D�@�����4@Y���i�!?��hzl�@����ٿ�#��D�@�����4@Y���i�!?��hzl�@����ٿ�#��D�@�����4@Y���i�!?��hzl�@����ٿ�#��D�@�����4@Y���i�!?��hzl�@?�ل�ٿ��t�{�@]�����3@e��j_�!?���B�@ϯ�K*�ٿ	��0R��@ns@�4@1��!?�u���5�@ϯ�K*�ٿ	��0R��@ns@�4@1��!?�u���5�@	�Mҗٿ��pA�@��ej�4@����z�!?Ұ���@	�Mҗٿ��pA�@��ej�4@����z�!?Ұ���@_�*ٿ�~����@6�h�-4@T�,|�!?�(ӝ+�@o��:S�ٿ6�E4��@��(��3@�:w4	�!?o`��j�@o��:S�ٿ6�E4��@��(��3@�:w4	�!?o`��j�@o��:S�ٿ6�E4��@��(��3@�:w4	�!?o`��j�@o��:S�ٿ6�E4��@��(��3@�:w4	�!?o`��j�@1��f�ٿu���*�@p��$s�3@�Ec �!?!e��'��@1��f�ٿu���*�@p��$s�3@�Ec �!?!e��'��@1��f�ٿu���*�@p��$s�3@�Ec �!?!e��'��@1��f�ٿu���*�@p��$s�3@�Ec �!?!e��'��@1��f�ٿu���*�@p��$s�3@�Ec �!?!e��'��@�o@�T�ٿ3popU��@7�D4c�3@
�c��!?Fn(���@�o@�T�ٿ3popU��@7�D4c�3@
�c��!?Fn(���@�o@�T�ٿ3popU��@7�D4c�3@
�c��!?Fn(���@�o@�T�ٿ3popU��@7�D4c�3@
�c��!?Fn(���@��)�ٿz�jz��@�޷3��3@\��C�!?4kiO�:�@��)�ٿz�jz��@�޷3��3@\��C�!?4kiO�:�@��)�ٿz�jz��@�޷3��3@\��C�!?4kiO�:�@���ٿy5I^��@���k&�3@ĺX�!?��0�)�@���ٿy5I^��@���k&�3@ĺX�!?��0�)�@���ٿy5I^��@���k&�3@ĺX�!?��0�)�@���ٿy5I^��@���k&�3@ĺX�!?��0�)�@�!��ٿ�>�ܲ��@��/P1�3@�9W�!?�C>t �@�!��ٿ�>�ܲ��@��/P1�3@�9W�!?�C>t �@�!��ٿ�>�ܲ��@��/P1�3@�9W�!?�C>t �@�!��ٿ�>�ܲ��@��/P1�3@�9W�!?�C>t �@�!��ٿ�>�ܲ��@��/P1�3@�9W�!?�C>t �@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@2p�ٿj2�h��@>}v��3@���^�!?4��E��@�f�ȗ�ٿ@mт��@d�j���3@�9�垐!?��>�,��@h�sJ�ٿ��s?{�@�i����3@
>�<�!?�6 ����@h�sJ�ٿ��s?{�@�i����3@
>�<�!?�6 ����@h�sJ�ٿ��s?{�@�i����3@
>�<�!?�6 ����@t���ٿ�\7"4��@z?	��3@����!?E��O�*�@t���ٿ�\7"4��@z?	��3@����!?E��O�*�@t���ٿ�\7"4��@z?	��3@����!?E��O�*�@�HU��ٿ�{|��X�@>+��3@.m���!? ׽��E�@�HU��ٿ�{|��X�@>+��3@.m���!? ׽��E�@�HU��ٿ�{|��X�@>+��3@.m���!? ׽��E�@�HU��ٿ�{|��X�@>+��3@.m���!? ׽��E�@�HU��ٿ�{|��X�@>+��3@.m���!? ׽��E�@����ٿ0�H"���@[����3@�򃞡�!?�1 �E�@����ٿ0�H"���@[����3@�򃞡�!?�1 �E�@����ٿ0�H"���@[����3@�򃞡�!?�1 �E�@����ٿ0�H"���@[����3@�򃞡�!?�1 �E�@�W���ٿ�e�O��@B?�'��3@?�7���!?�\h�@�W���ٿ�e�O��@B?�'��3@?�7���!?�\h�@H��{N�ٿ�n��P��@*����4@).�L�!?XT� w�@H��{N�ٿ�n��P��@*����4@).�L�!?XT� w�@H��{N�ٿ�n��P��@*����4@).�L�!?XT� w�@H��{N�ٿ�n��P��@*����4@).�L�!?XT� w�@���ΐٿy���?�@0D1�i4@a0pc1�!???E���@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@JC��ٿ
�\5t�@ߡ[��4@�)�Q�!?ѐ��p��@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�8�(q�ٿ 3�!r�@��~s�4@�2%߫�!?�
�DĴ@�;]&�ٿ�О3&,�@2`��3@�:p���!?��1;״@�K�O��ٿ�ķkEz�@��Qe�3@�{�?�!?T�eI
��@�K�O��ٿ�ķkEz�@��Qe�3@�{�?�!?T�eI
��@�K�O��ٿ�ķkEz�@��Qe�3@�{�?�!?T�eI
��@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@�� �U�ٿq��Hf�@�i}�4@�V!�8�!?�
8K���@��;��ٿ1②��@��Fp�4@�|�+�!?߽/�m�@��;��ٿ1②��@��Fp�4@�|�+�!?߽/�m�@��;��ٿ1②��@��Fp�4@�|�+�!?߽/�m�@b:�Y��ٿ��%�@<����3@��nA�!?j\�8�*�@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@��f�4�ٿ(*�+��@���9�3@;B��(�!?CA�-��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@'9��+�ٿM�+O��@���p�3@�'_8h�!?D���>��@���s�ٿ]uP����@��ܻ��3@�\	$g�!?�}�u8,�@���s�ٿ]uP����@��ܻ��3@�\	$g�!?�}�u8,�@���s�ٿ]uP����@��ܻ��3@�\	$g�!?�}�u8,�@G�1��ٿ?��߇�@�p�%��3@����?�!?�}�,�@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@>�/�C�ٿ��<���@�p�U�3@�eظR�!?W��~��@J�ǹ��ٿ��\�Ti�@�D�/`�3@��spm�!?0&4znJ�@J�ǹ��ٿ��\�Ti�@�D�/`�3@��spm�!?0&4znJ�@��If�ٿ�$-� �@�?'s�3@=\!v�!?����q�@���]Ŗٿ-'ږ��@?�[�3@�l0��!?m�x�`��@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@����S�ٿH{�8-�@�c��{�3@��R�!?�%�Heȵ@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@���q�ٿ[eT���@6AD��3@�l����!?�Ҵ�Zz�@QPh&��ٿ\::q��@�o1}��3@��9>�!?�0�fĵ@QPh&��ٿ\::q��@�o1}��3@��9>�!?�0�fĵ@QPh&��ٿ\::q��@�o1}��3@��9>�!?�0�fĵ@QPh&��ٿ\::q��@�o1}��3@��9>�!?�0�fĵ@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@�>d�ٿ)���jl�@�w��3@�J�r�!?��U-� �@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@F�#�ٿ"�%͉��@:�2)�3@�+"y�!?�`�4Kk�@�N=�T�ٿ��) 	9�@��z9�3@��n�!?��l�W��@e�l�ٿn�%�\�@����3@�>ˬ��!?A�@�刵@e�l�ٿn�%�\�@����3@�>ˬ��!?A�@�刵@e�l�ٿn�%�\�@����3@�>ˬ��!?A�@�刵@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@�����ٿZ� �J��@-��� �3@B�C�h�!?#�{��@��ܜ.�ٿ��j3DQ�@!�=�y�3@`�;A�!?S<fF�m�@��ܜ.�ٿ��j3DQ�@!�=�y�3@`�;A�!?S<fF�m�@��ܜ.�ٿ��j3DQ�@!�=�y�3@`�;A�!?S<fF�m�@EGa�r�ٿ��)_��@���-t�3@j��k�!?h'6<�@EGa�r�ٿ��)_��@���-t�3@j��k�!?h'6<�@EGa�r�ٿ��)_��@���-t�3@j��k�!?h'6<�@EGa�r�ٿ��)_��@���-t�3@j��k�!?h'6<�@EGa�r�ٿ��)_��@���-t�3@j��k�!?h'6<�@i�9f��ٿJό� d�@~�w��3@�rbg�!?i����@i�9f��ٿJό� d�@~�w��3@�rbg�!?i����@i�9f��ٿJό� d�@~�w��3@�rbg�!?i����@��#��ٿ�L�]��@i��3@l�DI�!?g�^V"�@��#��ٿ�L�]��@i��3@l�DI�!?g�^V"�@��#��ٿ�L�]��@i��3@l�DI�!?g�^V"�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@lW��ʓٿ��쐈�@�t���3@O�4�K�!?Ko|�B�@�)C�ޗٿ��sE|��@ɦ�'<�3@��9=7�!?f�a�Z��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�e{ڙٿ��]���@�X`���3@�+m��!?\^2��@�!�:�ٿX�*����@H(2��3@M'�H��!?b8����@�!�:�ٿX�*����@H(2��3@M'�H��!?b8����@�����ٿ�髁ں�@S�l��3@`{�j��!?ת�iǵ@�����ٿ�髁ں�@S�l��3@`{�j��!?ת�iǵ@�����ٿ�髁ں�@S�l��3@`{�j��!?ת�iǵ@�����ٿ�髁ں�@S�l��3@`{�j��!?ת�iǵ@�:z���ٿ��/��@����3@β���!?�z��
�@�:z���ٿ��/��@����3@β���!?�z��
�@�>�x�ٿ�M[?�b�@�����3@_pj��!?(P/��@q+y��ٿ���pN�@k�.!*�3@��3���!?����^�@��N<�ٿŷL<���@�-
� 4@��'��!?D��s�H�@��N<�ٿŷL<���@�-
� 4@��'��!?D��s�H�@��8��ٿPefz1��@?c[Q�3@z�;��!?x�	�ll�@o-���ٿ5�`Y���@Y�؊D�3@�Q��!?Ŗ�B:�@o-���ٿ5�`Y���@Y�؊D�3@�Q��!?Ŗ�B:�@o-���ٿ5�`Y���@Y�؊D�3@�Q��!?Ŗ�B:�@>!�g�ٿ����@�Qߥ��3@݋�8�!?�A��u��@>!�g�ٿ����@�Qߥ��3@݋�8�!?�A��u��@>!�g�ٿ����@�Qߥ��3@݋�8�!?�A��u��@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@��}��ٿ�"��Dc�@a�!��3@���|5�!?�`�%@�@f8z��ٿoiO�u�@����3@ӑE�O�!?�(���r�@����ٿ��MR���@��.6�3@^�)�#�!?~�U�5�@����ٿ��MR���@��.6�3@^�)�#�!?~�U�5�@����ٿ��MR���@��.6�3@^�)�#�!?~�U�5�@����ٿ��MR���@��.6�3@^�)�#�!?~�U�5�@����ٿ��MR���@��.6�3@^�)�#�!?~�U�5�@*�,^�ٿ��
���@�rYL�4@M���%�!?rƚ�@*�,^�ٿ��
���@�rYL�4@M���%�!?rƚ�@*�,^�ٿ��
���@�rYL�4@M���%�!?rƚ�@*�,^�ٿ��
���@�rYL�4@M���%�!?rƚ�@�?�vדٿ9v׬Z�@��Ԅ��3@Y�Q�w�!?U�˱�l�@�?�vדٿ9v׬Z�@��Ԅ��3@Y�Q�w�!?U�˱�l�@�?�vדٿ9v׬Z�@��Ԅ��3@Y�Q�w�!?U�˱�l�@�����ٿ��W�S�@Y�+���3@|4�z�!?͊��.�@�����ٿ��W�S�@Y�+���3@|4�z�!?͊��.�@�����ٿ��W�S�@Y�+���3@|4�z�!?͊��.�@�����ٿ��W�S�@Y�+���3@|4�z�!?͊��.�@/[�@�ٿ2�\8f�@�1;��3@��F��!?�:6a��@/[�@�ٿ2�\8f�@�1;��3@��F��!?�:6a��@/[�@�ٿ2�\8f�@�1;��3@��F��!?�:6a��@/[�@�ٿ2�\8f�@�1;��3@��F��!?�:6a��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@û[ ��ٿ�^N��@xD�a��3@���vP�!?=�J��@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@�[(P�ٿ���}��@�����3@��-!X�!?p���@`,��c�ٿ�~�r��@���.�3@�k��<�!?1�E�@�Q���ٿSOVy��@P��3�3@�O|O}�!?�ʁS��@�Q���ٿSOVy��@P��3�3@�O|O}�!?�ʁS��@�Q���ٿSOVy��@P��3�3@�O|O}�!?�ʁS��@�Q���ٿSOVy��@P��3�3@�O|O}�!?�ʁS��@�Q���ٿSOVy��@P��3�3@�O|O}�!?�ʁS��@ ����ٿ�e+�ɵ�@���9�3@�G�_B�!?�x?�?�@�_�z�ٿ�Mmv���@�6h�v�3@��n�!?Z�{Ӵ@�_�z�ٿ�Mmv���@�6h�v�3@��n�!?Z�{Ӵ@�_�z�ٿ�Mmv���@�6h�v�3@��n�!?Z�{Ӵ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@�Vl_U�ٿ���f�I�@��k��3@�~�!?�!6�Xܴ@��ty9�ٿN��� ��@����d4@DQ���!?\ŭ�;�@��ty9�ٿN��� ��@����d4@DQ���!?\ŭ�;�@��ty9�ٿN��� ��@����d4@DQ���!?\ŭ�;�@��ty9�ٿN��� ��@����d4@DQ���!?\ŭ�;�@��ty9�ٿN��� ��@����d4@DQ���!?\ŭ�;�@s��ّٿ�,�����@6���4@�(���!?쬏���@s��ّٿ�,�����@6���4@�(���!?쬏���@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@iê��ٿ��tx��@���c�3@:�hc�!?���R5%�@�l�	j�ٿ{*�����@�d^^�3@��| �!?�S�	���@�l�	j�ٿ{*�����@�d^^�3@��| �!?�S�	���@�l�	j�ٿ{*�����@�d^^�3@��| �!?�S�	���@�l�	j�ٿ{*�����@�d^^�3@��| �!?�S�	���@�l�	j�ٿ{*�����@�d^^�3@��| �!?�S�	���@P�2�ٿ|"8�^��@���$H�3@��g6|�!?��-��R�@c�����ٿ��'i�(�@��HW��3@ۜ�퇐!?��X�7�@c�����ٿ��'i�(�@��HW��3@ۜ�퇐!?��X�7�@�q���ٿ�q2����@2+���3@qFzh�!?t���d�@�3n疏ٿ���g6�@q3��s�3@�+Q��!?u�+�C�@�3n疏ٿ���g6�@q3��s�3@�+Q��!?u�+�C�@�3n疏ٿ���g6�@q3��s�3@�+Q��!?u�+�C�@�3n疏ٿ���g6�@q3��s�3@�+Q��!?u�+�C�@�O��ٿ.�UfDi�@����P�3@���Y�!?Q����|�@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@0�眒ٿ�{L!׮�@y��-�3@��CdB�!?��L���@�6M�8�ٿ�?�J0�@��u?��3@ʌ�p�!?�eU�@�6M�8�ٿ�?�J0�@��u?��3@ʌ�p�!?�eU�@�6M�8�ٿ�?�J0�@��u?��3@ʌ�p�!?�eU�@7�3���ٿ�.����@0s���3@λx.�!?����@7�3���ٿ�.����@0s���3@λx.�!?����@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@K�����ٿ�Ah����@-c�3@��Y9�!?p��JH´@��}��ٿ���@�@�z���3@�����!?�@o�@�lƃ�ٿ���8�@H'աi�3@�k,c�!??�`�X�@�lƃ�ٿ���8�@H'աi�3@�k,c�!??�`�X�@�_#���ٿ�۠����@U�n�6�3@42{V	�!?���[�@�_#���ٿ�۠����@U�n�6�3@42{V	�!?���[�@�_#���ٿ�۠����@U�n�6�3@42{V	�!?���[�@�_o�ٿ��9���@�WUB�3@��*,�!?ܶj!е@8�D�@�ٿ��L@ �@$�R�Y�3@$�1�!?>?nq���@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�v|�ٿ]�r�q��@g�+Sh�3@����!?'���ĵ@�n����ٿ�nϞ[e�@�2��J4@{�s1�!?��n�J�@�n����ٿ�nϞ[e�@�2��J4@{�s1�!?��n�J�@~�%��ٿ$��V��@���{14@��@>'�!?M"r�@~�%��ٿ$��V��@���{14@��@>'�!?M"r�@K���ٿ�#Zy+��@�lӂ�3@<�fo�!?��q��I�@K���ٿ�#Zy+��@�lӂ�3@<�fo�!?��q��I�@Ḅ�?�ٿ,3�-3��@��`���3@M:!�m�!?YǓ���@��4�m�ٿFk����@�"v.�3@�[�!?y��!o�@��4�m�ٿFk����@�"v.�3@�[�!?y��!o�@��4�m�ٿFk����@�"v.�3@�[�!?y��!o�@��4�m�ٿFk����@�"v.�3@�[�!?y��!o�@��4�m�ٿFk����@�"v.�3@�[�!?y��!o�@@Q�ٿ$���M�@�ܥp��3@N���4�!?4յ���@@Q�ٿ$���M�@�ܥp��3@N���4�!?4յ���@@Q�ٿ$���M�@�ܥp��3@N���4�!?4յ���@d��0�ٿ�;��K��@l�����3@�hyW	�!?��!�o�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@�w_`�ٿ��<.�@$;����3@�@��2�!?����b�@f�;�ٿ�K`+ �@��s{��3@�sb1�!?�|C0�v�@f�;�ٿ�K`+ �@��s{��3@�sb1�!?�|C0�v�@f�;�ٿ�K`+ �@��s{��3@�sb1�!?�|C0�v�@f�;�ٿ�K`+ �@��s{��3@�sb1�!?�|C0�v�@�>-�ٿ-���a�@���Ko4@�i�#�!?Kr��@�m;|�ٿ�k�Y��@���w4@�mm�L�!?�����@Q��i�ٿ#�M�m�@4*���3@���7�!?Ш�᝷�@Q��i�ٿ#�M�m�@4*���3@���7�!?Ш�᝷�@Q��i�ٿ#�M�m�@4*���3@���7�!?Ш�᝷�@Q��i�ٿ#�M�m�@4*���3@���7�!?Ш�᝷�@Q��i�ٿ#�M�m�@4*���3@���7�!?Ш�᝷�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@�}���ٿ�tT?���@{Y���3@�8�( �!?��D�q�@��խ�ٿ�%ߡ��@���_�3@��:8�!?�/㿴@.��	�ٿ�˪�$��@����L�3@���F�!?#Vƪy�@.��	�ٿ�˪�$��@����L�3@���F�!?#Vƪy�@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@��7���ٿ��֗�@��>��3@�.R9�!?����@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@-���Z�ٿBV� �@>%D��3@��3P�!?��8𢆴@�Յ�}�ٿNM�wl�@�����3@`+i+z�!?3 ��NM�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@���T�ٿ�47��@�WJ��3@�0I4|�!?�6C�x�@�Zv�\�ٿ�{:�8��@]&|�3@�Z���!?�[D�0�@�7J��ٿS���e�@�^� 4@%N�x�!?�b��쳴@�7J��ٿS���e�@�^� 4@%N�x�!?�b��쳴@�Y'�ٿ�� �aT�@?O�^�3@Wv��&�!?�n��u��@�Y'�ٿ�� �aT�@?O�^�3@Wv��&�!?�n��u��@�Y'�ٿ�� �aT�@?O�^�3@Wv��&�!?�n��u��@�Y'�ٿ�� �aT�@?O�^�3@Wv��&�!?�n��u��@���ʔٿUm��U�@H�8LJ�3@�i�'�!?��k�p�@���ʔٿUm��U�@H�8LJ�3@�i�'�!?��k�p�@���ʔٿUm��U�@H�8LJ�3@�i�'�!?��k�p�@nu�ߖٿqx�C�>�@
��t,�3@i]�T�!?��_��W�@w-8,]�ٿs.��,P�@g!���3@a@c.�!?���x�ȴ@w-8,]�ٿs.��,P�@g!���3@a@c.�!?���x�ȴ@w-8,]�ٿs.��,P�@g!���3@a@c.�!?���x�ȴ@w-8,]�ٿs.��,P�@g!���3@a@c.�!?���x�ȴ@w-8,]�ٿs.��,P�@g!���3@a@c.�!?���x�ȴ@���ՙ�ٿ���r5�@�|)�X�3@���@��!?��"C��@���ՙ�ٿ���r5�@�|)�X�3@���@��!?��"C��@u��ٿ�#�j��@��=Փ�3@��R���!?��д@u��ٿ�#�j��@��=Փ�3@��R���!?��д@��N��ٿ<0m�9�@������3@��XhE�!?�4�1?Q�@��N��ٿ<0m�9�@������3@��XhE�!?�4�1?Q�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@#�$w~�ٿv�k� ��@Cz9+�3@���<�!?b���`'�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@]L���ٿ�NwZ��@d�SI��3@�=GkS�!?���L�n�@\��j�ٿ����@�����3@�wֈ�!?��Q�
µ@\��j�ٿ����@�����3@�wֈ�!?��Q�
µ@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@kW�*��ٿ�u���@��S���3@;e�l�!?�`�Ĥ�@�5��ٿ�t�ц�@BQl�w�3@z��H��!?�>0	��@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@X�̻��ٿcWQG��@�����3@�7TА!?�ΠIô@Ѡ�7=�ٿ����a4�@�wr�5�3@��)Ȑ!?�0�L�@�:-�ȓٿu��hn�@����4@ ��w�!?�4�u@�@q$��n�ٿD�]N�@Ƚ8���3@�Uc�d�!?������@q$��n�ٿD�]N�@Ƚ8���3@�Uc�d�!?������@q$��n�ٿD�]N�@Ƚ8���3@�Uc�d�!?������@q$��n�ٿD�]N�@Ƚ8���3@�Uc�d�!?������@q$��n�ٿD�]N�@Ƚ8���3@�Uc�d�!?������@�7�P��ٿf�$�@5�@�&~��3@�|���!?]����@�7�P��ٿf�$�@5�@�&~��3@�|���!?]����@�7�P��ٿf�$�@5�@�&~��3@�|���!?]����@�qI�ٿ�	���@�M��3@['Cُ!?�PX�!�@�qI�ٿ�	���@�M��3@['Cُ!?�PX�!�@���.��ٿ��~j-��@���3@�>����!?�a��'�@���.��ٿ��~j-��@���3@�>����!?�a��'�@���.��ٿ��~j-��@���3@�>����!?�a��'�@���.��ٿ��~j-��@���3@�>����!?�a��'�@���.��ٿ��~j-��@���3@�>����!?�a��'�@y�0�o�ٿ�$�%�@'�����3@���I�!?���l@ʴ@y�0�o�ٿ�$�%�@'�����3@���I�!?���l@ʴ@y�0�o�ٿ�$�%�@'�����3@���I�!?���l@ʴ@y�0�o�ٿ�$�%�@'�����3@���I�!?���l@ʴ@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@m0\t��ٿ��E*���@���3@���X�!?L7N�O�@p|-+7�ٿ�E�S��@�2_��3@ �X��!?A�l�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@ȧ���ٿ���ʣ�@���/D�3@3�9&�!?p4"`	*�@+j��ٿ��@l�Q�@2q@˵�3@��J�!?M'��I�@+j��ٿ��@l�Q�@2q@˵�3@��J�!?M'��I�@+j��ٿ��@l�Q�@2q@˵�3@��J�!?M'��I�@+j��ٿ��@l�Q�@2q@˵�3@��J�!?M'��I�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@���r�ٿS��dJ]�@\1eW�3@X��\.�!?N���4�@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@�I���ٿ�c�V���@zPMD��3@�B�uޏ!?����@5�ѡ�ٿ��Le]�@�Ӯ12�3@�=�Ə!?�՝����@\��t�ٿ�8�p?=�@f��3@ܕL�!?����;4�@\��t�ٿ�8�p?=�@f��3@ܕL�!?����;4�@\��t�ٿ�8�p?=�@f��3@ܕL�!?����;4�@\��t�ٿ�8�p?=�@f��3@ܕL�!?����;4�@8�ܧ�ٿ0Ɲ��^�@U�E �3@3q�!?�x�!�@�,-�ٿ{]6�F�@|��_�3@�Mk�!?����)�@�,-�ٿ{]6�F�@|��_�3@�Mk�!?����)�@�,-�ٿ{]6�F�@|��_�3@�Mk�!?����)�@�D����ٿ���2\�@K+��R�3@I�c��!?��m�mܴ@�D����ٿ���2\�@K+��R�3@I�c��!?��m�mܴ@�D����ٿ���2\�@K+��R�3@I�c��!?��m�mܴ@�D����ٿ���2\�@K+��R�3@I�c��!?��m�mܴ@�کCy�ٿҺk�
�@��!���3@KHԑ�!?�� �6�@�کCy�ٿҺk�
�@��!���3@KHԑ�!?�� �6�@d�S>A�ٿB�	\��@(��7��3@d$�Ǔ�!?���@d�S>A�ٿB�	\��@(��7��3@d$�Ǔ�!?���@9o|�ҕٿg���@B�-h� 4@��Iy�!?�3��	�@���"�ٿ� 6���@ ����3@��b�!?�����޴@���"�ٿ� 6���@ ����3@��b�!?�����޴@���"�ٿ� 6���@ ����3@��b�!?�����޴@���"�ٿ� 6���@ ����3@��b�!?�����޴@���"�ٿ� 6���@ ����3@��b�!?�����޴@� �ٿ_$���@a�����3@�o�!?��ھ��@� �ٿ_$���@a�����3@�o�!?��ھ��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�_e�_�ٿ����Y�@B�g�3@�(#%d�!?�n�I;��@�O�ٿe����@����3@'ab��!?wc�F}�@�Č��ٿR(���-�@.��E�3@h5�!?������@�K��ٿ�r��M!�@]_����3@���B�!?�sB&���@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@:ܰ��ٿ����m�@�\���3@�bu�!?D�B�@�zS��ٿ��^(��@ـ���3@�c9>�!?f��8���@�O1�ٿ,���;�@�,�+��3@Q���G�!?�A>ь��@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�E3� �ٿ�aP��j�@�~�n�3@�\�7�!?� �ô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@�PJqu�ٿ-�c�*_�@+�i��3@V��+u�!?� ENô@8�C�ٿ8,.s,�@�� "��3@�����!?�g�1]�@8�C�ٿ8,.s,�@�� "��3@�����!?�g�1]�@+oT^�ٿ�TI]��@���s� 4@#�[�M�!?��L�FB�@+oT^�ٿ�TI]��@���s� 4@#�[�M�!?��L�FB�@+oT^�ٿ�TI]��@���s� 4@#�[�M�!?��L�FB�@�/ ��ٿ�!א�~�@��߭� 4@<$����!?�o�D�c�@�/ ��ٿ�!א�~�@��߭� 4@<$����!?�o�D�c�@�/ ��ٿ�!א�~�@��߭� 4@<$����!?�o�D�c�@�/ ��ٿ�!א�~�@��߭� 4@<$����!?�o�D�c�@�/ ��ٿ�!א�~�@��߭� 4@<$����!?�o�D�c�@W��s�ٿ���lخ�@,�����3@JO��!?]�)�T�@W��s�ٿ���lخ�@,�����3@JO��!?]�)�T�@�f��ؑٿǑ����@�(�2��3@���u�!?�;ڴ@��Ԁ�ٿ_6;u��@���31�3@Kt�p��!?�.�����@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@��Sʗٿ6�;v�@�,����3@���[�!?r�Ǒ�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@ �f�^�ٿ��*g��@'���3@3S��^�!?��ݳOP�@���ٿ�<yec�@z�{���3@���\�!?ӪA�!�@���ٿ�<yec�@z�{���3@���\�!?ӪA�!�@���ٿ�<yec�@z�{���3@���\�!?ӪA�!�@���ٿ�<yec�@z�{���3@���\�!?ӪA�!�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@�8n2�ٿ֖�HkR�@yƦ�)�3@v�vB�!?�fUw=�@*�a��ٿxw�9�5�@���n��3@�=LΏ!?��ʬ���@*�a��ٿxw�9�5�@���n��3@�=LΏ!?��ʬ���@*�a��ٿxw�9�5�@���n��3@�=LΏ!?��ʬ���@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@���-�ٿ}+��@<�aH�4@��O�!?J]<	H=�@�/g�@�ٿ�_+�$�@閤e�3@��4�!?%]b�I�@�/g�@�ٿ�_+�$�@閤e�3@��4�!?%]b�I�@�/g�@�ٿ�_+�$�@閤e�3@��4�!?%]b�I�@�^Ϋy�ٿ?��pt��@-�8���3@N����!?�bmޫ2�@�^Ϋy�ٿ?��pt��@-�8���3@N����!?�bmޫ2�@�^Ϋy�ٿ?��pt��@-�8���3@N����!?�bmޫ2�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@&>�5�ٿ$m��$�@���Ae�3@5��O�!?��*?.�@�J��#�ٿ�,/i.�@̻\B�4@�}?Џ�!?��ks�@�J��#�ٿ�,/i.�@̻\B�4@�}?Џ�!?��ks�@�J��#�ٿ�,/i.�@̻\B�4@�}?Џ�!?��ks�@�J��#�ٿ�,/i.�@̻\B�4@�}?Џ�!?��ks�@�J��#�ٿ�,/i.�@̻\B�4@�}?Џ�!?��ks�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@+d�?B�ٿ�����@Eև*�4@RʛL�!?G��}�@�i}R$�ٿV�B�a��@D9��4@���|!�!?�i(�m��@��:�!�ٿL�@��@��J7�4@P��ޏ!?#ƻ�ZP�@��>ݢٿr ��u�@R� j��3@�	�!?�s���>�@��>ݢٿr ��u�@R� j��3@�	�!?�s���>�@(5��ٿ��v��@�����3@�	�� �!?��]G�@(5��ٿ��v��@�����3@�	�� �!?��]G�@(5��ٿ��v��@�����3@�	�� �!?��]G�@(5��ٿ��v��@�����3@�	�� �!?��]G�@wmU�G�ٿ�ߚ�;@�@<=�\��3@��=��!?m!�ܴ@wmU�G�ٿ�ߚ�;@�@<=�\��3@��=��!?m!�ܴ@wmU�G�ٿ�ߚ�;@�@<=�\��3@��=��!?m!�ܴ@wmU�G�ٿ�ߚ�;@�@<=�\��3@��=��!?m!�ܴ@�f�,�ٿc���1M�@��=ab�3@���P�!?��\1��@|F�"�ٿ�ֆ[�D�@�����3@_��<d�!?!�>Z�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@�i©Ȗٿ8s�L�
�@#�@{0�3@�;�1�!?�]���)�@C9pKv�ٿ����9�@�ДJ��3@��9kQ�!?�P$�@&4aL�ٿ3_rA2�@{�1���3@'!0O0�!?RRH9��@&4aL�ٿ3_rA2�@{�1���3@'!0O0�!?RRH9��@���j�ٿ�i.��J�@3F�F�3@c�L�\�!?k�B�|C�@���j�ٿ�i.��J�@3F�F�3@c�L�\�!?k�B�|C�@���j�ٿ�i.��J�@3F�F�3@c�L�\�!?k�B�|C�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@xGӒٿ�v��@~���2�3@����f�!?��{B�@3�*ߊ�ٿ|� {�@ފ���3@�)}�"�!?��`�3��@3�*ߊ�ٿ|� {�@ފ���3@�)}�"�!?��`�3��@3�*ߊ�ٿ|� {�@ފ���3@�)}�"�!?��`�3��@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@�#�봑ٿ��!Hʼ�@��)�3@k[>�!?���c���@Rv��ٿ^��a.�@�?��v�3@�W�e�!?�M�d�ʴ@Rv��ٿ^��a.�@�?��v�3@�W�e�!?�M�d�ʴ@Bc�3N�ٿ�?�q�a�@`׹��3@*�eY�!?�<E�H��@Bc�3N�ٿ�?�q�a�@`׹��3@*�eY�!?�<E�H��@Bc�3N�ٿ�?�q�a�@`׹��3@*�eY�!?�<E�H��@Bc�3N�ٿ�?�q�a�@`׹��3@*�eY�!?�<E�H��@Bc�3N�ٿ�?�q�a�@`׹��3@*�eY�!?�<E�H��@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�o1̕ٿnfDI�G�@~A��4@X5�h�!?E�?Ѵ@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@�hY��ٿ�֜E�3�@0ʮ&��3@�#v2��!? �}]�H�@���K�ٿ�["���@�
�d�3@{�[ڴ�!?������@Og���ٿ��|���@eHOC��3@���7��!?��5`��@'�a��ٿA$��s�@�XP��3@���̐!?q.Qb��@'�a��ٿA$��s�@�XP��3@���̐!?q.Qb��@'�a��ٿA$��s�@�XP��3@���̐!?q.Qb��@���*b�ٿ�,�ki;�@t���l�3@JW��!?��P��@"M�;�ٿ2sɞ�@�#x��3@&ý̐!?��?��@"M�;�ٿ2sɞ�@�#x��3@&ý̐!?��?��@"M�;�ٿ2sɞ�@�#x��3@&ý̐!?��?��@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@��Y0��ٿ �����@�L7��3@=�EӐ!?Q����L�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@V���ٿiIat��@�o���3@�O�Ӝ�!?K ��q�@��_}j�ٿ~)C����@�-�E�3@�4�!?�+j?�մ@��_}j�ٿ~)C����@�-�E�3@�4�!?�+j?�մ@Gc}'Ԕٿ�*�|�"�@���4@��q�!?*Z��|�@Gc}'Ԕٿ�*�|�"�@���4@��q�!?*Z��|�@Gc}'Ԕٿ�*�|�"�@���4@��q�!?*Z��|�@�� ���ٿ�0qLW��@�����3@���m�!?nNG(J�@�� ���ٿ�0qLW��@�����3@���m�!?nNG(J�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@vZ՘ٿ��a���@""���3@�=ς�!? Jr��:�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@.�m=@�ٿ��wۢ�@�( ���3@'�v�)�!?�����@�@�-679�ٿ>9)���@T�~���3@��jȐ�!?H�z�=�@�j�y�ٿ�QA�\��@K��w�4@:#u]�!?�g�ÏE�@�j�y�ٿ�QA�\��@K��w�4@:#u]�!?�g�ÏE�@�*ɚ��ٿ !�"C�@[��J�3@I�#��!?��zzU�@�*ɚ��ٿ !�"C�@[��J�3@I�#��!?��zzU�@�*ɚ��ٿ !�"C�@[��J�3@I�#��!?��zzU�@�ގ���ٿ��Bf�@������3@��D�[�!?r���@�ގ���ٿ��Bf�@������3@��D�[�!?r���@�ގ���ٿ��Bf�@������3@��D�[�!?r���@�ގ���ٿ��Bf�@������3@��D�[�!?r���@�ގ���ٿ��Bf�@������3@��D�[�!?r���@�ގ���ٿ��Bf�@������3@��D�[�!?r���@d�(��ٿo��%�S�@Q]i0��3@b��!?�Cd؆h�@�����ٿ��G��@�);�3@�XjW�!?�9֛w�@�O����ٿ-������@�y���3@h6�|��!?v�#T��@�O����ٿ-������@�y���3@h6�|��!?v�#T��@�O����ٿ-������@�y���3@h6�|��!?v�#T��@�O����ٿ-������@�y���3@h6�|��!?v�#T��@�O����ٿ-������@�y���3@h6�|��!?v�#T��@q��v�ٿ�:�d�l�@�zbh� 4@����?�!?`I��t�@�.��ٿ����@
�ғ�3@�#���!?7i%�p�@�.��ٿ����@
�ғ�3@�#���!?7i%�p�@�.��ٿ����@
�ғ�3@�#���!?7i%�p�@�.��ٿ����@
�ғ�3@�#���!?7i%�p�@�.��ٿ����@
�ғ�3@�#���!?7i%�p�@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@�� U�ٿf�n�J�@��3@�Ff�!?��^�P��@J>i|B�ٿ��xx>��@;����3@�E���!?o�L���@J>i|B�ٿ��xx>��@;����3@�E���!?o�L���@�\��k�ٿ~�x�j�@�P0��3@��tO��!?P�S�?�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@q�;݄�ٿ�ZK��@{�dp��3@aw�I�!?7��E�@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@D.|��ٿ}�V��y�@���1��3@�� ��!?���{��@'�n�ٿx����@�G�/4@�?Ј�!?@�	bĵ@'�n�ٿx����@�G�/4@�?Ј�!?@�	bĵ@�	�삙ٿY�0
j��@d�N���3@J4��)�!?��Ԡ�ϵ@�	�삙ٿY�0
j��@d�N���3@J4��)�!?��Ԡ�ϵ@�	�삙ٿY�0
j��@d�N���3@J4��)�!?��Ԡ�ϵ@>��ݘٿ�<o7���@)tāU�3@�E�L!�!?']�#J�@O9r�[�ٿ�	ϥ���@ކ��3@�e��l�!?c�dӁ��@O9r�[�ٿ�	ϥ���@ކ��3@�e��l�!?c�dӁ��@,�Iߜٿ��r��Y�@KJ��3@E>��R�!?F��'��@,�Iߜٿ��r��Y�@KJ��3@E>��R�!?F��'��@,�Iߜٿ��r��Y�@KJ��3@E>��R�!?F��'��@��%�_�ٿ�vu}�@��<~e4@����T�!?b/��7|�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@/�b��ٿ����@�����3@��A4�!?,+��v�@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@�D7��ٿ2����@�6��3@�>a��!?���'Դ@���ٿ��̉�Ŀ@�L����3@��U�B�!?��{ႃ�@���ٿ��̉�Ŀ@�L����3@��U�B�!?��{ႃ�@{��hs�ٿl���#�@1���`�3@U?EX��!?�f8�е@{��hs�ٿl���#�@1���`�3@U?EX��!?�f8�е@{��hs�ٿl���#�@1���`�3@U?EX��!?�f8�е@�yG�ٿ��L����@��C��3@h�B���!?���,�_�@�yG�ٿ��L����@��C��3@h�B���!?���,�_�@�yG�ٿ��L����@��C��3@h�B���!?���,�_�@!���֙ٿ$���d�@A=�TA�3@���h�!?v}��H��@!���֙ٿ$���d�@A=�TA�3@���h�!?v}��H��@�v#��ٿg��6:��@�F'D4@�Y��B�!?��ΟɁ�@i�[��ٿo~y�(A�@����I 4@��0K�!?*^?M.W�@i�[��ٿo~y�(A�@����I 4@��0K�!?*^?M.W�@�pj0��ٿ�T��]�@�	�4@�%��P�!?%���g��@�pj0��ٿ�T��]�@�	�4@�%��P�!?%���g��@�pj0��ٿ�T��]�@�	�4@�%��P�!?%���g��@�D�k�ٿѓ���@���i�3@�J�y�!?��%-D!�@�D�k�ٿѓ���@���i�3@�J�y�!?��%-D!�@��e��ٿ���1��@e����4@FIL�l�!?��7{�@��e��ٿ���1��@e����4@FIL�l�!?��7{�@��e��ٿ���1��@e����4@FIL�l�!?��7{�@�V�[�ٿ�;��Q8�@9y�jz
4@�Zbv�!?�%\�Q=�@�oaL�ٿW:����@Tg�.�3@��9�!?݄�մ@�oaL�ٿW:����@Tg�.�3@��9�!?݄�մ@�oaL�ٿW:����@Tg�.�3@��9�!?݄�մ@�oaL�ٿW:����@Tg�.�3@��9�!?݄�մ@�oaL�ٿW:����@Tg�.�3@��9�!?݄�մ@�~7f�ٿ��u=�@��4�3@d��!?�`M&;�@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�0�w�ٿ�U-����@����3@��]R!�!?�����@�g���ٿ6��LV(�@?�fL�3@�,ʉ�!?��5,
�@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@��	���ٿ����W�@�|����3@�P�C�!?�.�� �@i�p�ٿFU���@@�����3@�n/�!?�D����@i�p�ٿFU���@@�����3@�n/�!?�D����@i�p�ٿFU���@@�����3@�n/�!?�D����@����Ñٿ@
c̠�@:�N4��3@�F��!?ӷ���ٴ@����Ñٿ@
c̠�@:�N4��3@�F��!?ӷ���ٴ@����Ñٿ@
c̠�@:�N4��3@�F��!?ӷ���ٴ@����Ñٿ@
c̠�@:�N4��3@�F��!?ӷ���ٴ@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@��)�h�ٿʈ��o�@�܈��3@Y�wQ��!?����+k�@����_�ٿtm� ���@���3@~f9x�!?�����״@T��wW�ٿ�*Mm؄�@CsH�]4@;-�Q�!?���Ij��@T��wW�ٿ�*Mm؄�@CsH�]4@;-�Q�!?���Ij��@T��wW�ٿ�*Mm؄�@CsH�]4@;-�Q�!?���Ij��@T��wW�ٿ�*Mm؄�@CsH�]4@;-�Q�!?���Ij��@��XŜٿD��L�@h�&M-�3@�5�$ѐ!?�8Ps�b�@��XŜٿD��L�@h�&M-�3@�5�$ѐ!?�8Ps�b�@��XŜٿD��L�@h�&M-�3@�5�$ѐ!?�8Ps�b�@��XŜٿD��L�@h�&M-�3@�5�$ѐ!?�8Ps�b�@��XŜٿD��L�@h�&M-�3@�5�$ѐ!?�8Ps�b�@�`���ٿ�Ux��@��#��3@;�И�!?p�ڇFԳ@:&��4�ٿy��l^�@Gy�{�4@��W�!?7���8�@:&��4�ٿy��l^�@Gy�{�4@��W�!?7���8�@��ʑٿ��=��@j�!���3@p[%�d�!?.#᯿��@��ʑٿ��=��@j�!���3@p[%�d�!?.#᯿��@����R�ٿ�;�V��@3;hA�3@� u`��!?�V:|R�@����R�ٿ�;�V��@3;hA�3@� u`��!?�V:|R�@����R�ٿ�;�V��@3;hA�3@� u`��!?�V:|R�@����R�ٿ�;�V��@3;hA�3@� u`��!?�V:|R�@����R�ٿ�;�V��@3;hA�3@� u`��!?�V:|R�@**��ٿS��
� �@7��|�3@ߌ�!?�i-r�V�@**��ٿS��
� �@7��|�3@ߌ�!?�i-r�V�@**��ٿS��
� �@7��|�3@ߌ�!?�i-r�V�@**��ٿS��
� �@7��|�3@ߌ�!?�i-r�V�@~�R���ٿO$}g��@��Ȯ�3@=q3��!?��E���@~�R���ٿO$}g��@��Ȯ�3@=q3��!?��E���@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@L�ɏ��ٿ
`����@��f��3@��*h�!?l.�/�@�4��ٿ �+q8>�@��SM�3@x;#V�!?���@��K.�ٿ^��2��@c�*$U�3@I�*�Y�!?\w�9'�@��K.�ٿ^��2��@c�*$U�3@I�*�Y�!?\w�9'�@��K.�ٿ^��2��@c�*$U�3@I�*�Y�!?\w�9'�@��K.�ٿ^��2��@c�*$U�3@I�*�Y�!?\w�9'�@��K.�ٿ^��2��@c�*$U�3@I�*�Y�!?\w�9'�@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@:�ew�ٿo�J��@���6N�3@�1\X�!?��\���@�M}.U�ٿr���4*�@�qx�B�3@5��fZ�!?"�2�S�@�M}.U�ٿr���4*�@�qx�B�3@5��fZ�!?"�2�S�@�M}.U�ٿr���4*�@�qx�B�3@5��fZ�!?"�2�S�@�M}.U�ٿr���4*�@�qx�B�3@5��fZ�!?"�2�S�@���ٿ}������@G5���3@�{-Xɏ!?��r�B�@���ٿ}������@G5���3@�{-Xɏ!?��r�B�@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�ti¥�ٿ3yXt���@�
B��3@o��!?L�l���@�U�$�ٿ��^�L�@�Ȁ��3@��M�!?�(AP���@�U�$�ٿ��^�L�@�Ȁ��3@��M�!?�(AP���@�U�$�ٿ��^�L�@�Ȁ��3@��M�!?�(AP���@�U�$�ٿ��^�L�@�Ȁ��3@��M�!?�(AP���@�U�$�ٿ��^�L�@�Ȁ��3@��M�!?�(AP���@S@�sy�ٿ%
cl��@n���<�3@���6�!?�ି�ϴ@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@ P�E�ٿ���~�@���P��3@$�w�!?;v)���@̓+��ٿ��ϳ���@	�#F��3@4�fӏ!?�*6j@�@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@TfR��ٿk���@��d��3@���!?��Qr9Ĵ@��[�̒ٿ��p�=b�@�I*nY�3@��I�.�!?�K�㛿�@��[�̒ٿ��p�=b�@�I*nY�3@��I�.�!?�K�㛿�@��[�̒ٿ��p�=b�@�I*nY�3@��I�.�!?�K�㛿�@��[�̒ٿ��p�=b�@�I*nY�3@��I�.�!?�K�㛿�@��[�̒ٿ��p�=b�@�I*nY�3@��I�.�!?�K�㛿�@��Y��ٿ�<���@%�j���3@��$"�!?����D�@��Y��ٿ�<���@%�j���3@��$"�!?����D�@��Y��ٿ�<���@%�j���3@��$"�!?����D�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@=�Q ��ٿ�r�>��@LPg!4@��2.�!?���ae?�@�M(o��ٿ�Dآ�@�#�4@%��A�!? A�G^5�@�M(o��ٿ�Dآ�@�#�4@%��A�!? A�G^5�@�M(o��ٿ�Dآ�@�#�4@%��A�!? A�G^5�@�M(o��ٿ�Dآ�@�#�4@%��A�!? A�G^5�@@��0A�ٿ��T���@�:��7�3@�i� я!?4��N�@@��0A�ٿ��T���@�:��7�3@�i� я!?4��N�@@��0A�ٿ��T���@�:��7�3@�i� я!?4��N�@ؠs��ٿ�O,��L�@q�פ��3@z��]�!?K��{e��@ؠs��ٿ�O,��L�@q�פ��3@z��]�!?K��{e��@ؠs��ٿ�O,��L�@q�פ��3@z��]�!?K��{e��@X`�N�ٿ��Z����@}��bi 4@��!-C�!?㦀SR��@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@�|S��ٿH�h�o�@��J���3@��jc�!?˱T��[�@� (��ٿ��Lc+��@wr��3@�")$
�!?y;�YBV�@u�tI�ٿB�t��@�F�`�3@��6��!?l�Љ´@u�tI�ٿB�t��@�F�`�3@��6��!?l�Љ´@u�tI�ٿB�t��@�F�`�3@��6��!?l�Љ´@u�tI�ٿB�t��@�F�`�3@��6��!?l�Љ´@u�tI�ٿB�t��@�F�`�3@��6��!?l�Љ´@X �t�ٿ7�ђ�K�@OS��3@t��%�!?F�5����@X �t�ٿ7�ђ�K�@OS��3@t��%�!?F�5����@���~p�ٿ�tv�W�@�u�Q��3@{�32�!?:�X2��@���~p�ٿ�tv�W�@�u�Q��3@{�32�!?:�X2��@���~p�ٿ�tv�W�@�u�Q��3@{�32�!?:�X2��@���~p�ٿ�tv�W�@�u�Q��3@{�32�!?:�X2��@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@`��z�ٿ]��{P�@)a�=�3@� �LX�!?�o��4�@���"��ٿd�Y/�:�@$�nfL�3@����p�!?!}��F8�@���"��ٿd�Y/�:�@$�nfL�3@����p�!?!}��F8�@���"��ٿd�Y/�:�@$�nfL�3@����p�!?!}��F8�@���"��ٿd�Y/�:�@$�nfL�3@����p�!?!}��F8�@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@�Jr��ٿ�3Yi�v�@�C,���3@��B5i�!?�ͅ5��@(� Rz�ٿ�sn����@_�ܡo�3@:W6� �!?0���B��@(� Rz�ٿ�sn����@_�ܡo�3@:W6� �!?0���B��@���W|�ٿ/[m��G�@�h�|�4@q3%	=�!?ȣ!Xv]�@���W|�ٿ/[m��G�@�h�|�4@q3%	=�!?ȣ!Xv]�@<�?E�ٿ_blw��@.%�4@�?��!?�s�?�|�@<�?E�ٿ_blw��@.%�4@�?��!?�s�?�|�@<�?E�ٿ_blw��@.%�4@�?��!?�s�?�|�@MKl��ٿ��}�BW�@��'�R�3@��q�!?`�����@MKl��ٿ��}�BW�@��'�R�3@��q�!?`�����@MKl��ٿ��}�BW�@��'�R�3@��q�!?`�����@e(t=�ٿ�bZ����@:��Q�3@2�>(��!?��m=Y��@e(t=�ٿ�bZ����@:��Q�3@2�>(��!?��m=Y��@t7��Z�ٿ���C�6�@RU��z4@NY}j�!?Ϣ@�յ@������ٿ�9��c�@�~�k��3@��\=�!?�sq\��@������ٿ�9��c�@�~�k��3@��\=�!?�sq\��@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@?ϡŘٿ�7pFG��@L$y��3@���T�!?�l�!���@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@!N��N�ٿ(E���L�@R���3@Tq�A�!?h��@��<⊛ٿ��M��@i��R!�3@E��{B�!?D��8^̴@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@h�$Wיٿ̎ �	7�@�ܒR,�3@�+/�!?4�T�
�@-M� �ٿ����@�2l���3@s��A�!?R��̒�@-M� �ٿ����@�2l���3@s��A�!?R��̒�@-M� �ٿ����@�2l���3@s��A�!?R��̒�@u�^Ԙٿ-F����@��mY�3@�2fwڏ!?x�x���@������ٿ*���8?�@[}�H��3@l�~"��!?�!��ܴ@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@$�x�ğٿ�D�K�@�Q%���3@3�p�!?ͪ�`�O�@���Иٿ/�R���@����3@܅)k�!?�i�x��@���Иٿ/�R���@����3@܅)k�!?�i�x��@���Иٿ/�R���@����3@܅)k�!?�i�x��@���Иٿ/�R���@����3@܅)k�!?�i�x��@B�Q��ٿn6f�r�@��T�3@(��2��!?��-���@B�Q��ٿn6f�r�@��T�3@(��2��!?��-���@06H�ٿ!^����@�ω���3@)�}�y�!?Z'��#\�@06H�ٿ!^����@�ω���3@)�}�y�!?Z'��#\�@��tJ
�ٿMИ��@{�P���3@�Ƙp�!?K�j�qǴ@��tJ
�ٿMИ��@{�P���3@�Ƙp�!?K�j�qǴ@�Еٿ��·Y�@���v�3@~,OqR�!?��Ac�P�@�Еٿ��·Y�@���v�3@~,OqR�!?��Ac�P�@�Еٿ��·Y�@���v�3@~,OqR�!?��Ac�P�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@f�=ߕٿLg�j�9�@����6�3@�W;�!?^{�v*�@*櫔ٿ%�b�+��@�_�-�3@�c�u�!?�[��5�@*櫔ٿ%�b�+��@�_�-�3@�c�u�!?�[��5�@*櫔ٿ%�b�+��@�_�-�3@�c�u�!?�[��5�@�x]�n�ٿ����y��@������3@�	Vߌ�!?�k~tJ�@�k��T�ٿ�� ��7�@O�o��3@3jdޓ�!?_L���[�@�k��T�ٿ�� ��7�@O�o��3@3jdޓ�!?_L���[�@�k��T�ٿ�� ��7�@O�o��3@3jdޓ�!?_L���[�@�k��T�ٿ�� ��7�@O�o��3@3jdޓ�!?_L���[�@8�j���ٿٖ�	�@o��E�4@�o=�r�!?���Xˑ�@8�j���ٿٖ�	�@o��E�4@�o=�r�!?���Xˑ�@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@5"DȘ�ٿ�^� e�@l�^]F�3@,�+g4�!?ڒY��@����ٿl�Ii���@3����3@�`���!?�����Q�@����ٿl�Ii���@3����3@�`���!?�����Q�@tG08�ٿ�|��I��@>*�j�4@ٌ\�ڏ!?��)���@tG08�ٿ�|��I��@>*�j�4@ٌ\�ڏ!?��)���@tG08�ٿ�|��I��@>*�j�4@ٌ\�ڏ!?��)���@tG08�ٿ�|��I��@>*�j�4@ٌ\�ڏ!?��)���@tG08�ٿ�|��I��@>*�j�4@ٌ\�ڏ!?��)���@��襌�ٿ�5@����@ST�4@�=φ�!?���UL�@�	�x͚ٿ7��(��@_u�:4@�Fƽ~�!?�U��\s�@�~���ٿ�8��'�@Y_�)d4@~��'0�!?t���閴@�~���ٿ�8��'�@Y_�)d4@~��'0�!?t���閴@�~���ٿ�8��'�@Y_�)d4@~��'0�!?t���閴@�~���ٿ�8��'�@Y_�)d4@~��'0�!?t���閴@��%A��ٿ���k��@~�'�x4@1�U���!?�R�� ��@.d�K�ٿ7��c�@Մ�I��3@�_!x�!?�:���@.d�K�ٿ7��c�@Մ�I��3@�_!x�!?�:���@�_H5Q�ٿn��j�v�@w�����3@�T�x�!?�~���&�@5 Qz��ٿ�E)O:��@��]T�3@�QL(��!? '���?�@5 Qz��ٿ�E)O:��@��]T�3@�QL(��!? '���?�@5 Qz��ٿ�E)O:��@��]T�3@�QL(��!? '���?�@�_
�ٿX�s%d�@>y",Q�3@��TO�!?t@�G�޴@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@��؋�ٿ�B��-�@�Q���3@Õ��n�!?7HQm�$�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@RŽMq�ٿ��y��u�@�����3@�m�1b�!?Q�)I{�@��)���ٿH!-�@̨|@d�3@
��h�!?�����@��)���ٿH!-�@̨|@d�3@
��h�!?�����@��)���ٿH!-�@̨|@d�3@
��h�!?�����@��)���ٿH!-�@̨|@d�3@
��h�!?�����@�U�e��ٿ�Cfsr[�@�$���3@��Q�m�!?�X@����@/q��o�ٿ�����@'jR^e�3@���!?�i�|�@/q��o�ٿ�����@'jR^e�3@���!?�i�|�@/q��o�ٿ�����@'jR^e�3@���!?�i�|�@/q��o�ٿ�����@'jR^e�3@���!?�i�|�@/q��o�ٿ�����@'jR^e�3@���!?�i�|�@�����ٿ��oHJ�@ZN���3@���Z�!? �ѷ�>�@�����ٿ��oHJ�@ZN���3@���Z�!? �ѷ�>�@�����ٿ��oHJ�@ZN���3@���Z�!? �ѷ�>�@�����ٿ��oHJ�@ZN���3@���Z�!? �ѷ�>�@h1�C��ٿq��!��@
�+_+�3@�_ᐐ!?�����Y�@yrU\�ٿUή���@���+D4@t�I�|�!?XjY�:�@yrU\�ٿUή���@���+D4@t�I�|�!?XjY�:�@��ٙٿi�q����@nI��y�3@N�bb��!?N1���@eLO��ٿ�����@�^ �(�3@ �ꑣ�!?��dİI�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@~,��ٿ�Lr.�%�@h�P��4@��{]א!?���t�@�u:��ٿ�\�(�@�A9q4@�p3��!?)��k�@�u:��ٿ�\�(�@�A9q4@�p3��!?)��k�@�u:��ٿ�\�(�@�A9q4@�p3��!?)��k�@�u:��ٿ�\�(�@�A9q4@�p3��!?)��k�@*�};͙ٿZ�#-2V�@��p��3@k�w�ʐ!?umG����@*�};͙ٿZ�#-2V�@��p��3@k�w�ʐ!?umG����@P4$�ٿ�zZ�x��@���3@�E ���!?�, ۴@:��]�ٿ��=:V��@�NL�3@���ߐ!?[�G>�Դ@���b�ٿ,�,�O�@�S/(��3@@�M��!?vбuM��@���b�ٿ,�,�O�@�S/(��3@@�M��!?vбuM��@���b�ٿ,�,�O�@�S/(��3@@�M��!?vбuM��@���b�ٿ,�,�O�@�S/(��3@@�M��!?vбuM��@���b�ٿ,�,�O�@�S/(��3@@�M��!?vбuM��@Q���&�ٿע�U*�@�϶���3@��l	�!?X�rFS�@Q���&�ٿע�U*�@�϶���3@��l	�!?X�rFS�@Q���&�ٿע�U*�@�϶���3@��l	�!?X�rFS�@�a����ٿ��¯
�@s��B�3@��K��!?|k,��@�a����ٿ��¯
�@s��B�3@��K��!?|k,��@�a����ٿ��¯
�@s��B�3@��K��!?|k,��@�M�.;�ٿ�b�4>�@�v��w�3@��<��!?��o�	q�@f�i�$�ٿAX,��o�@���u��3@Qw�*��!?�0c���@f�i�$�ٿAX,��o�@���u��3@Qw�*��!?�0c���@f�i�$�ٿAX,��o�@���u��3@Qw�*��!?�0c���@f�i�$�ٿAX,��o�@���u��3@Qw�*��!?�0c���@��U?��ٿ��{k��@?b�ϥ�3@@x��w�!?�%Gn/�@��U?��ٿ��{k��@?b�ϥ�3@@x��w�!?�%Gn/�@��U?��ٿ��{k��@?b�ϥ�3@@x��w�!?�%Gn/�@��U?��ٿ��{k��@?b�ϥ�3@@x��w�!?�%Gn/�@��q�&�ٿVy�n��@��Nq��3@�۽�!?���|��@��q�&�ٿVy�n��@��Nq��3@�۽�!?���|��@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@!d
���ٿ!��#<�@=�!�3@�ؿ�!?.��Dג�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@�t��}�ٿ�}��@�=J�3@D��À�!?�Αڛ�@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@-�t�6�ٿS���@��j�~�3@ѩ��!?e^G���@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@Q�|Y�ٿBf(����@Zܨ�Q�3@V�A�!?Y�QN�u�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�p�e��ٿ��fO�A�@��3�]�3@	q�{}�!?�ӎ�Q8�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�I�	�ٿ�i0��@,,�W�3@���h�!?�K�
h�@�����ٿ��\��@H����3@+�7�!?�iɅ�'�@�����ٿ��\��@H����3@+�7�!?�iɅ�'�@�����ٿ��\��@H����3@+�7�!?�iɅ�'�@�=儛ٿ�H9�5��@D�ςH�3@k����!?�z5��)�@���_��ٿ
:����@�Y���3@UB�Z(�!?�ej���@���_��ٿ
:����@�Y���3@UB�Z(�!?�ej���@���_��ٿ
:����@�Y���3@UB�Z(�!?�ej���@���_��ٿ
:����@�Y���3@UB�Z(�!?�ej���@���_��ٿ
:����@�Y���3@UB�Z(�!?�ej���@���h�ٿPk;�e�@wc	�T�3@��FN�!?�v�G���@C�V��ٿ��X��@�%�p�3@v_a+�!?<��*���@C�V��ٿ��X��@�%�p�3@v_a+�!?<��*���@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@�f1P��ٿ�n�A`��@�^J�F�3@B�)�5�!?�	�<:e�@
ɔ�V�ٿz�'z �@��w
4@�|b�B�!?�a���ε@Wx T̗ٿR.Q�@�*E�4@.o8Ik�!?�п8ն�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@���(��ٿJ��J�@�k���3@$��;��!?)�UT�{�@�T���ٿ�&)�"�@��$�[�3@���W�!?����S�@�T���ٿ�&)�"�@��$�[�3@���W�!?����S�@�T���ٿ�&)�"�@��$�[�3@���W�!?����S�@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�M��,�ٿ&��	�@���3@�:Y�V�!?3�����@�g�*ّٿ���wQ�@5J���3@cC�|�!?9�2K�@�g�*ّٿ���wQ�@5J���3@cC�|�!?9�2K�@�g�*ّٿ���wQ�@5J���3@cC�|�!?9�2K�@�g�*ّٿ���wQ�@5J���3@cC�|�!?9�2K�@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@���Xۘٿ�\��;�@�����3@�K��{�!?�z��@g��2��ٿ��ܟ���@�?*�l�3@�cwne�!?7��˴@d�3�ٿ����x�@�l��A�3@#X����!?N�͗��@d�3�ٿ����x�@�l��A�3@#X����!?N�͗��@�a���ٿ�t��&�@��}��3@>ΐ�!?��b��e�@M@�P��ٿ?��>G�@�}���3@�s�!?/�����@M@�P��ٿ?��>G�@�}���3@�s�!?/�����@M@�P��ٿ?��>G�@�}���3@�s�!?/�����@M@�P��ٿ?��>G�@�}���3@�s�!?/�����@����ٿ�6t�E�@�)v"�3@ߎ��!?��u50�@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@�=���ٿ�!�7W��@D�c���3@7D�	�!?/�����@��g�ٿ^�����@P�44�3@��<>��!?sCԴ@��g�ٿ^�����@P�44�3@��<>��!?sCԴ@��g�ٿ^�����@P�44�3@��<>��!?sCԴ@��g�ٿ^�����@P�44�3@��<>��!?sCԴ@��g�ٿ^�����@P�44�3@��<>��!?sCԴ@�;וٿ�3����@}����3@fE�.��!?��/�@�;וٿ�3����@}����3@fE�.��!?��/�@�L���ٿRo_����@����4@�q0\�!?��i���@�L���ٿRo_����@����4@�q0\�!?��i���@E���ٿj�
��l�@9���3@���I�!?����O�@E���ٿj�
��l�@9���3@���I�!?����O�@E���ٿj�
��l�@9���3@���I�!?����O�@E���ٿj�
��l�@9���3@���I�!?����O�@٢���ٿ,y+��@���b��3@�K�	5�!?ŝ��w��@٢���ٿ,y+��@���b��3@�K�	5�!?ŝ��w��@)�dw��ٿ�5e\��@�w�.�3@`��"*�!?�x)h��@)�dw��ٿ�5e\��@�w�.�3@`��"*�!?�x)h��@������ٿ�<�2,�@⡤���3@��?��!?�x���C�@���sO�ٿ�QX{7�@�l憹�3@�LKk:�!?-�M���@���sO�ٿ�QX{7�@�l憹�3@�LKk:�!?-�M���@���sO�ٿ�QX{7�@�l憹�3@�LKk:�!?-�M���@���sO�ٿ�QX{7�@�l憹�3@�LKk:�!?-�M���@��qp0�ٿoM�{ٹ�@��V��3@g�����!?"�e��@�=�k�ٿ�ɾ�v�@`�;	�3@����!? ��M�@�=�k�ٿ�ɾ�v�@`�;	�3@����!? ��M�@�=�k�ٿ�ɾ�v�@`�;	�3@����!? ��M�@�=�k�ٿ�ɾ�v�@`�;	�3@����!? ��M�@�5̌�ٿ�oߎ�<�@Ϭ}�3@s��>G�!?��6��~�@�5̌�ٿ�oߎ�<�@Ϭ}�3@s��>G�!?��6��~�@�5̌�ٿ�oߎ�<�@Ϭ}�3@s��>G�!?��6��~�@�y����ٿq����@Q�B ��3@+�'Q�!?{�ў�@�y����ٿq����@Q�B ��3@+�'Q�!?{�ў�@�y����ٿq����@Q�B ��3@+�'Q�!?{�ў�@�y����ٿq����@Q�B ��3@+�'Q�!?{�ў�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@x�b$�ٿ!n�)�g�@W߯���3@�_�1�!?$�N*$�@
'�z)�ٿq�Q���@}J�ǣ�3@�0ETI�!?���˺�@
'�z)�ٿq�Q���@}J�ǣ�3@�0ETI�!?���˺�@��,0ٔٿ*�ލd�@R*��3@zb&;�!?�S���l�@��,0ٔٿ*�ލd�@R*��3@zb&;�!?�S���l�@��,0ٔٿ*�ލd�@R*��3@zb&;�!?�S���l�@��,0ٔٿ*�ލd�@R*��3@zb&;�!?�S���l�@��,0ٔٿ*�ލd�@R*��3@zb&;�!?�S���l�@2��l�ٿ�!h�@2uX��4@�G�o�!?�Xk)o�@2��l�ٿ�!h�@2uX��4@�G�o�!?�Xk)o�@2��l�ٿ�!h�@2uX��4@�G�o�!?�Xk)o�@2��l�ٿ�!h�@2uX��4@�G�o�!?�Xk)o�@2��l�ٿ�!h�@2uX��4@�G�o�!?�Xk)o�@�<��ٿ��vc�@֠��P4@=	�<�!?Oz2�@�Hr���ٿ�����@AU�G�3@�\��!?Eskh�Q�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@X�3��ٿ0�]�c0�@x3�
4@ɾ�	�!?$n��p�@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@���:��ٿ���1QO�@b�n&�4@�y0D:�!?O�����@�]�s��ٿ%���#�@�CɅ4@��1�!?w,�yF�@�]�s��ٿ%���#�@�CɅ4@��1�!?w,�yF�@�]�s��ٿ%���#�@�CɅ4@��1�!?w,�yF�@";��-�ٿ�=�����@�Qk`l�3@U�ɑo�!?j2BW��@";��-�ٿ�=�����@�Qk`l�3@U�ɑo�!?j2BW��@��`��ٿ��y��@o~�)�3@u'� =�!?xÆ�?�@��`��ٿ��y��@o~�)�3@u'� =�!?xÆ�?�@��`��ٿ��y��@o~�)�3@u'� =�!?xÆ�?�@��`��ٿ��y��@o~�)�3@u'� =�!?xÆ�?�@��`��ٿ��y��@o~�)�3@u'� =�!?xÆ�?�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@K��-�ٿq��ۖ(�@���W�3@{-�B�!?hF#�]�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@�Դ���ٿ� G���@��<�3@��'��!?�O\x�H�@P�i��ٿ�+�:��@�`�L�3@xz�3m�!?�,,K��@�O��ٿ��E���@`�p���3@%1|,��!?��uB!�@�O��ٿ��E���@`�p���3@%1|,��!?��uB!�@�_l�ٿ���t�@�����3@�`"��!?X����@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@|��e2�ٿ��*\�@�nH�t4@@܄�{�!?��Rn�D�@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@4\����ٿ�
i���@X��b��3@���Ys�!?%0w�w��@��֜��ٿM��d\��@��6N��3@�zofӏ!?���ƒ�@��֜��ٿM��d\��@��6N��3@�zofӏ!?���ƒ�@��֜��ٿM��d\��@��6N��3@�zofӏ!?���ƒ�@��֜��ٿM��d\��@��6N��3@�zofӏ!?���ƒ�@��֜��ٿM��d\��@��6N��3@�zofӏ!?���ƒ�@n�5�ٿ��N���@�3���3@9�Fڏ!?��;*�K�@�D���ٿ��w�� �@${lm��3@H6���!?���H�&�@�/�s��ٿ{L�<,�@'�C���3@Of��&�!?���W���@�/�s��ٿ{L�<,�@'�C���3@Of��&�!?���W���@�/�s��ٿ{L�<,�@'�C���3@Of��&�!?���W���@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@rmd��ٿ����h|�@9�4@Y����!?�(��Re�@��ÒٿD<�4���@�O��c4@�p�Qa�!?*��(��@R��јٿ&/8�#�@�����4@B��!?1�"�YE�@��s�Q�ٿ��:�w�@�Y�>+�3@(���#�!?ߺ����@��s�Q�ٿ��:�w�@�Y�>+�3@(���#�!?ߺ����@����ٿ⊧���@�Jz<��3@髻S(�!?��C�@����ٿ⊧���@�Jz<��3@髻S(�!?��C�@����ٿ⊧���@�Jz<��3@髻S(�!?��C�@����ٿ⊧���@�Jz<��3@髻S(�!?��C�@����ٿ⊧���@�Jz<��3@髻S(�!?��C�@(��%�ٿ'�Wͳk�@��/�3@�w�؏!?���(�@(��%�ٿ'�Wͳk�@��/�3@�w�؏!?���(�@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@+�y���ٿ�/����@���lF�3@Yl)4�!?Я�N+ȴ@��7�ٿ8u*����@b3�DC�3@��uY�!?g4���@��7�ٿ8u*����@b3�DC�3@��uY�!?g4���@^�~���ٿ:�qV7�@��O��3@D[�c��!?n���@^�~���ٿ:�qV7�@��O��3@D[�c��!?n���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�*�TP�ٿ˽(<��@(M�r�3@P(|ˊ�!?��h���@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�M.���ٿF��	�@��Vن�3@�<���!?��3c1�@�C��u�ٿ �܊�]�@�G>@�3@�0��m�!?sa��Y��@�C��u�ٿ �܊�]�@�G>@�3@�0��m�!?sa��Y��@�C��u�ٿ �܊�]�@�G>@�3@�0��m�!?sa��Y��@�I)�
�ٿ%�i����@���3@cP�3@�!?��-����@�I)�
�ٿ%�i����@���3@cP�3@�!?��-����@�I)�
�ٿ%�i����@���3@cP�3@�!?��-����@r��H�ٿ"��d��@)Y蛤�3@1��p�!?�#��@r��H�ٿ"��d��@)Y蛤�3@1��p�!?�#��@r��H�ٿ"��d��@)Y蛤�3@1��p�!?�#��@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@���P��ٿJ��V�@��T�e�3@]�1�t�!?���ܴ@����ɕٿቤɊ�@l&0�4�3@�����!?�LXO�@����ɕٿቤɊ�@l&0�4�3@�����!?�LXO�@����ɕٿቤɊ�@l&0�4�3@�����!?�LXO�@W�N�řٿW^.�@�/��"�3@�]��!?�ߜ��@W�N�řٿW^.�@�/��"�3@�]��!?�ߜ��@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@�0]�ٿU&�t�@?��}�3@�1S&�!?��V�W4�@b����ٿq-� ��@*��K�3@~�:r�!?	�j�3�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@b��yĘٿ/��%�@"��H��3@�*�3w�!?��\q�@a�T�v�ٿ_�m���@t0�^7�3@)�aG��!?��v��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@/�Zf�ٿ�&����@���ڳ�3@�W�a�!?�h�r��@x�~AÕٿ�� �n��@�Yc�/�3@
dV�h�!?��Mҵ@x�~AÕٿ�� �n��@�Yc�/�3@
dV�h�!?��Mҵ@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@��� �ٿ4cB�a�@�1�0�3@mĄV�!?�*Q�l��@^1M׉�ٿXw�o�I�@�2i�3@ExV�3�!?RTyש�@�e�l�ٿ��)��@�@A����3@���ŏ!?-��<�@�e�l�ٿ��)��@�@A����3@���ŏ!?-��<�@E�)�ٿ!��!%��@�B����3@�{���!?�t�����@E�)�ٿ!��!%��@�B����3@�{���!?�t�����@E�)�ٿ!��!%��@�B����3@�{���!?�t�����@E�)�ٿ!��!%��@�B����3@�{���!?�t�����@ISޛ~�ٿ�/��@�K~-�3@��ٓ�!?SM�+���@ISޛ~�ٿ�/��@�K~-�3@��ٓ�!?SM�+���@ISޛ~�ٿ�/��@�K~-�3@��ٓ�!?SM�+���@ISޛ~�ٿ�/��@�K~-�3@��ٓ�!?SM�+���@ISޛ~�ٿ�/��@�K~-�3@��ٓ�!?SM�+���@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�˧�ٿ���[V�@������3@���L@�!?l�ј�g�@�����ٿZ��
��@�ŉ���3@%�Z�!?F�蘆�@�����ٿZ��
��@�ŉ���3@%�Z�!?F�蘆�@�����ٿZ��
��@�ŉ���3@%�Z�!?F�蘆�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@�~�Q�ٿ�|�-$��@�����3@�q�b.�!?�s�;�L�@Y�ÙV�ٿB2���@����3@b(�y�!?E-#�z�@?ϰ���ٿt�;"��@��Y�3@�ט��!?���X�@?ϰ���ٿt�;"��@��Y�3@�ט��!?���X�@?ϰ���ٿt�;"��@��Y�3@�ט��!?���X�@W2�J�ٿw����@�A���3@�?-�v�!?���td�@W2�J�ٿw����@�A���3@�?-�v�!?���td�@�"��ٿs�.���@kfm���3@��K�M�!?_�B,*�@�"��ٿs�.���@kfm���3@��K�M�!?_�B,*�@���r�ٿ���
;�@3�fpT�3@��!?�YRW�@4s��,�ٿ)//#�@��7x��3@0����!?���P��@4s��,�ٿ)//#�@��7x��3@0����!?���P��@4s��,�ٿ)//#�@��7x��3@0����!?���P��@��v�ٿ��>6�"�@X���3@)j��F�!?w�Z�Nq�@��v�ٿ��>6�"�@X���3@)j��F�!?w�Z�Nq�@��v�ٿ��>6�"�@X���3@)j��F�!?w�Z�Nq�@��v�ٿ��>6�"�@X���3@)j��F�!?w�Z�Nq�@��v�ٿ��>6�"�@X���3@)j��F�!?w�Z�Nq�@c"���ٿ�A���.�@�|�W4@�.l�V�!?Bף�.A�@c"���ٿ�A���.�@�|�W4@�.l�V�!?Bף�.A�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@B��^�ٿW�7�)#�@��Ҩf�3@бd��!?�J�3�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�SJ�V�ٿ|V�jnc�@�Xup��3@E���Q�!?��i'0�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@�D�s�ٿ+zt��@h�[(s�3@=��9�!?\>m�;$�@Vy���ٿ� �d��@\+����3@��U�!?(��-���@Vy���ٿ� �d��@\+����3@��U�!?(��-���@Vy���ٿ� �d��@\+����3@��U�!?(��-���@���7�ٿ�O�p���@�[�T��3@�!e%�!?����	�@���7�ٿ�O�p���@�[�T��3@�!e%�!?����	�@���7�ٿ�O�p���@�[�T��3@�!e%�!?����	�@���7�ٿ�O�p���@�[�T��3@�!e%�!?����	�@���7�ٿ�O�p���@�[�T��3@�!e%�!?����	�@4�)>�ٿ�b�hD��@G����3@R#b~�!?�u��6�@4�)>�ٿ�b�hD��@G����3@R#b~�!?�u��6�@4�)>�ٿ�b�hD��@G����3@R#b~�!?�u��6�@�����ٿ��IJEL�@�Z�7r�3@�T�*��!?�����L�@XY��ٿu�Q����@��� 4@���'Y�!?Y)J�Ss�@XY��ٿu�Q����@��� 4@���'Y�!?Y)J�Ss�@XY��ٿu�Q����@��� 4@���'Y�!?Y)J�Ss�@XY��ٿu�Q����@��� 4@���'Y�!?Y)J�Ss�@XY��ٿu�Q����@��� 4@���'Y�!?Y)J�Ss�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@��<�N�ٿ̽�1��@�eg���3@K�n�q�!?�Y�l9�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@N|xܘٿ�����@�ʏ�3@c�p+A�!?��?3�@�:S�\�ٿE�lm@��@+����3@�M1>�!?�����@�
քA�ٿ������@V��"N�3@���n�!?�v�䬴@�
քA�ٿ������@V��"N�3@���n�!?�v�䬴@LAIӶ�ٿP�P#�=�@�g/���3@�v�LX�!?`'�k�@LAIӶ�ٿP�P#�=�@�g/���3@�v�LX�!?`'�k�@LAIӶ�ٿP�P#�=�@�g/���3@�v�LX�!?`'�k�@LAIӶ�ٿP�P#�=�@�g/���3@�v�LX�!?`'�k�@s�+�ٿ!�%���@JR�4@靽eU�!?\��0��@s�+�ٿ!�%���@JR�4@靽eU�!?\��0��@s�+�ٿ!�%���@JR�4@靽eU�!?\��0��@s�+�ٿ!�%���@JR�4@靽eU�!?\��0��@s�+�ٿ!�%���@JR�4@靽eU�!?\��0��@L�Z��ٿ�ˆ�{��@��h�3@�B�;�!?N��;�@L�Z��ٿ�ˆ�{��@��h�3@�B�;�!?N��;�@L�Z��ٿ�ˆ�{��@��h�3@�B�;�!?N��;�@L�Z��ٿ�ˆ�{��@��h�3@�B�;�!?N��;�@L�Z��ٿ�ˆ�{��@��h�3@�B�;�!?N��;�@�5A�ٿ��/,���@=D����3@�B#�z�!?�Ё�V�@�5A�ٿ��/,���@=D����3@�B#�z�!?�Ё�V�@�5A�ٿ��/,���@=D����3@�B#�z�!?�Ё�V�@e�Ф�ٿR��ϔc�@̨ϫ�3@�4��c�!?���'C�@e�Ф�ٿR��ϔc�@̨ϫ�3@�4��c�!?���'C�@e�Ф�ٿR��ϔc�@̨ϫ�3@�4��c�!?���'C�@e�Ф�ٿR��ϔc�@̨ϫ�3@�4��c�!?���'C�@{'�͛ٿ�����@�+ #��3@���"�!?S���L��@{'�͛ٿ�����@�+ #��3@���"�!?S���L��@{'�͛ٿ�����@�+ #��3@���"�!?S���L��@{'�͛ٿ�����@�+ #��3@���"�!?S���L��@{'�͛ٿ�����@�+ #��3@���"�!?S���L��@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@� �;��ٿ����J3�@������3@ �0�O�!?ٝ�Q�@���Rњٿr2����@D�<o�4@���S�!?$�G�t��@���Rњٿr2����@D�<o�4@���S�!?$�G�t��@����-�ٿ��΋\3�@f�Hj��3@Ӟ�](�!?���h�ʴ@����-�ٿ��΋\3�@f�Hj��3@Ӟ�](�!?���h�ʴ@����-�ٿ��΋\3�@f�Hj��3@Ӟ�](�!?���h�ʴ@����-�ٿ��΋\3�@f�Hj��3@Ӟ�](�!?���h�ʴ@:�?�n�ٿ-���d�@4��4@T��Jm�!?>���E�@:�?�n�ٿ-���d�@4��4@T��Jm�!?>���E�@:�?�n�ٿ-���d�@4��4@T��Jm�!?>���E�@:�?�n�ٿ-���d�@4��4@T��Jm�!?>���E�@��#�u�ٿ��"�@q,~;*4@�E�]?�!?Up���C�@��#�u�ٿ��"�@q,~;*4@�E�]?�!?Up���C�@��#�u�ٿ��"�@q,~;*4@�E�]?�!?Up���C�@��#�u�ٿ��"�@q,~;*4@�E�]?�!?Up���C�@��#�u�ٿ��"�@q,~;*4@�E�]?�!?Up���C�@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@� ��ٿ=jyPI�@��k�4@��!?��Kx��@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@��`�Вٿ_��q��@���E��3@!;qN�!?t҅-�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@֏�M�ٿ
�a���@��:��3@v�8��!?r ���j�@��ѫW�ٿQ�ZN�p�@������3@Z��	�!?�u	���@�1��?�ٿ�e׸g=�@��	� 4@-�X:�!?Y��@�1��?�ٿ�e׸g=�@��	� 4@-�X:�!?Y��@�1��?�ٿ�e׸g=�@��	� 4@-�X:�!?Y��@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@�[����ٿ�HRm<��@wQ��3@$��G�!?1�B倵@c�q�ٿ���ё�@�}0��3@��a�!?���B�@�5_��ٿ�`�7�@�
+���3@UVw4j�!?N8�PD�@�5_��ٿ�`�7�@�
+���3@UVw4j�!?N8�PD�@�5_��ٿ�`�7�@�
+���3@UVw4j�!?N8�PD�@�k�ę�ٿ���+��@���ul�3@�ˈQg�!?^Ťr�i�@J2xL͘ٿ�%4���@��G�@�3@���!?�)��	m�@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@���8'�ٿ=��4tn�@'#BP��3@��oƂ�!?B����@�6ŷ�ٿΌ�RV�@Dہ���3@�E����!?� ����@�6ŷ�ٿΌ�RV�@Dہ���3@�E����!?� ����@�6ŷ�ٿΌ�RV�@Dہ���3@�E����!?� ����@'(dz�ٿ+�#�/��@c8$0��3@�e.u[�!?�6��7V�@'(dz�ٿ+�#�/��@c8$0��3@�e.u[�!?�6��7V�@��'��ٿ秡���@M+�-�3@F�n<�!?1�m%�@��'��ٿ秡���@M+�-�3@F�n<�!?1�m%�@6C�-�ٿ$ƞ�2��@� �3@����q�!?R����0�@6C�-�ٿ$ƞ�2��@� �3@����q�!?R����0�@6C�-�ٿ$ƞ�2��@� �3@����q�!?R����0�@6C�-�ٿ$ƞ�2��@� �3@����q�!?R����0�@F����ٿ-���o��@�M���3@m:�,�!?��j﮴@��/��ٿ���ͣ>�@�@���3@�r��̏!?$�~R
O�@��/��ٿ���ͣ>�@�@���3@�r��̏!?$�~R
O�@7��ʘٿ�����B�@�]���3@�ל�!?N����@7��ʘٿ�����B�@�]���3@�ל�!?N����@7��ʘٿ�����B�@�]���3@�ל�!?N����@7��ʘٿ�����B�@�]���3@�ל�!?N����@�P���ٿ�3�����@��<!�3@�r�Kˏ!?����'��@ɦ��/�ٿ�"���D�@t[���3@�>�!�!?y/��?�@���h�ٿ��r����@LoVPX�3@��5��!?�
���@���h�ٿ��r����@LoVPX�3@��5��!?�
���@�X�#��ٿm�`,c�@
�q�z�3@��8��!?n�zjz��@�X�#��ٿm�`,c�@
�q�z�3@��8��!?n�zjz��@�X�#��ٿm�`,c�@
�q�z�3@��8��!?n�zjz��@�X�#��ٿm�`,c�@
�q�z�3@��8��!?n�zjz��@�X�#��ٿm�`,c�@
�q�z�3@��8��!?n�zjz��@��q�ٿ�X���j�@�<��v�3@Xs�"�!?��h��@��q�ٿ�X���j�@�<��v�3@Xs�"�!?��h��@9�}���ٿ;,�s���@MF��=�3@�t=�!?��*$t��@9�}���ٿ;,�s���@MF��=�3@�t=�!?��*$t��@9�}���ٿ;,�s���@MF��=�3@�t=�!?��*$t��@��ro[�ٿ�(����@�@Wb�3@n䘋R�!?�C���@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�5�b�ٿ
���[D�@l+�X��3@��")�!?�\��״@�?T��ٿ�����@���&��3@���P�!?4�����@�?T��ٿ�����@���&��3@���P�!?4�����@�?T��ٿ�����@���&��3@���P�!?4�����@a�b�Y�ٿz���Em�@-�h�3@���@!�!?�Q���<�@a�b�Y�ٿz���Em�@-�h�3@���@!�!?�Q���<�@�ژ�S�ٿ^6�]���@������3@����,�!?�}ꕠ̴@�ژ�S�ٿ^6�]���@������3@����,�!?�}ꕠ̴@�ژ�S�ٿ^6�]���@������3@����,�!?�}ꕠ̴@W*7e:�ٿS�FrkP�@vDS�4@�Vz�Y�!?��eT�@�ӎ�O�ٿ:Uc���@:5R
�3@�����!?�C�_�r�@������ٿ�޷���@(V��V4@��,�!�!?���\+�@������ٿ�޷���@(V��V4@��,�!�!?���\+�@ ��H�ٿ86�4���@��׉4@Zք�"�!?�x���ĵ@ ��H�ٿ86�4���@��׉4@Zք�"�!?�x���ĵ@ ��H�ٿ86�4���@��׉4@Zք�"�!?�x���ĵ@�+>���ٿ�k����@C��g�3@X����!?'�3����@�+>���ٿ�k����@C��g�3@X����!?'�3����@�l̥ٖٿ(���@t��	��3@�N�l�!?�-:��-�@�l̥ٖٿ(���@t��	��3@�N�l�!?�-:��-�@S~ņ%�ٿ�T���@��V'�3@i/�O6�!?��9��]�@�O.��ٿ򎐨j�@L{D_��3@�
�|�!?O��/�4�@�O.��ٿ򎐨j�@L{D_��3@�
�|�!?O��/�4�@�O.��ٿ򎐨j�@L{D_��3@�
�|�!?O��/�4�@��4^�ٿS�ws�@��3@��3P�!?,��N�P�@��4^�ٿS�ws�@��3@��3P�!?,��N�P�@td�{�ٿNT��@b�V���3@<�#�!?�ZX*=#�@td�{�ٿNT��@b�V���3@<�#�!?�ZX*=#�@td�{�ٿNT��@b�V���3@<�#�!?�ZX*=#�@td�{�ٿNT��@b�V���3@<�#�!?�ZX*=#�@td�{�ٿNT��@b�V���3@<�#�!?�ZX*=#�@�"��Вٿ(f�B�'�@5����3@o��yB�!?F�C���@�"��Вٿ(f�B�'�@5����3@o��yB�!?F�C���@!ʁ��ٿ��s'��@���zC�3@�{l�!?��W3Hz�@^�I�O�ٿ�j9�aV�@5��F�3@��;G�!?_�㗵@^�I�O�ٿ�j9�aV�@5��F�3@��;G�!?_�㗵@6����ٿB�&@D.�@��e��3@#��C1�!?�N$��@6����ٿB�&@D.�@��e��3@#��C1�!?�N$��@6����ٿB�&@D.�@��e��3@#��C1�!?�N$��@6����ٿB�&@D.�@��e��3@#��C1�!?�N$��@���ٿ�<�X�K�@�b/��3@��s5�!?�ho�
�@���ٿ�<�X�K�@�b/��3@��s5�!?�ho�
�@���ٿ�<�X�K�@�b/��3@��s5�!?�ho�
�@��t�ٿ�� ;���@���3@���{E�!?��O|*�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@G��wW�ٿBK��΢�@ְ˧4�3@�
GG�!?[�L�4�@��[�2�ٿ3f���@E_7��3@�X�aL�!?f�9{��@��ē�ٿG��n��@Z_[�`�3@�L0v@�!?}v��@��ē�ٿG��n��@Z_[�`�3@�L0v@�!?}v��@��ē�ٿG��n��@Z_[�`�3@�L0v@�!?}v��@��ē�ٿG��n��@Z_[�`�3@�L0v@�!?}v��@��ē�ٿG��n��@Z_[�`�3@�L0v@�!?}v��@9]I���ٿT~�ډ��@=�#Y��3@�]"x�!?"�D~(y�@9]I���ٿT~�ډ��@=�#Y��3@�]"x�!?"�D~(y�@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�.�qv�ٿ�M��@F�a���3@'���!?��9����@�����ٿ�/Bxq�@fJB&0�3@���x�!?����U�@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@���ٿ�;'(���@L��ː�3@��ï{�!?;��8մ@��͸�ٿ
�:@�R�@�#2��3@���s�!?�J-���@��͸�ٿ
�:@�R�@�#2��3@���s�!?�J-���@��͸�ٿ
�:@�R�@�#2��3@���s�!?�J-���@��͸�ٿ
�:@�R�@�#2��3@���s�!?�J-���@��&1\�ٿ~�4�'q�@d P�F�3@��(�!?���U�@��&1\�ٿ~�4�'q�@d P�F�3@��(�!?���U�@��&1\�ٿ~�4�'q�@d P�F�3@��(�!?���U�@����ќٿI�Z�%�@{jm���3@��eD�!?��XKL�@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@6J]�0�ٿ����@_��N�3@k���u�!?"��GQ��@[tied�ٿ��va���@΀�!��3@�}�̆�!?&ko�>��@[tied�ٿ��va���@΀�!��3@�}�̆�!?&ko�>��@��/��ٿP+	�@2�A�=�3@����!?is�.q�@��+�ٿ���%?O�@�G+ 4@����I�!?6$�˶�@��+�ٿ���%?O�@�G+ 4@����I�!?6$�˶�@��+�ٿ���%?O�@�G+ 4@����I�!?6$�˶�@��+�ٿ���%?O�@�G+ 4@����I�!?6$�˶�@��+�ٿ���%?O�@�G+ 4@����I�!?6$�˶�@��0ȝٿt��JG�@����A4@~sn.B�!?�����Ǵ@8��]�ٿo���@�e];�3@�/�Q�!?�����d�@8��]�ٿo���@�e];�3@�/�Q�!?�����d�@�	�ٿ��o k��@v��q 4@��jpO�!?g\�@�t֝ٿڀv���@SC;d4@���я�!?����L�@�t֝ٿڀv���@SC;d4@���я�!?����L�@�fDn�ٿ2Lb��-�@�h��b4@U�/Q��!?e�f8���@�fDn�ٿ2Lb��-�@�h��b4@U�/Q��!?e�f8���@2��� �ٿ�E-���@�m���3@	vu�w�!?���RO�@2��� �ٿ�E-���@�m���3@	vu�w�!?���RO�@2��� �ٿ�E-���@�m���3@	vu�w�!?���RO�@���U~�ٿ�	����@cnt<4@�򖳐!?&| �^�@���U~�ٿ�	����@cnt<4@�򖳐!?&| �^�@���U~�ٿ�	����@cnt<4@�򖳐!?&| �^�@h�#/��ٿ��f�#�@�+�ۢ4@=�;o��!?!���@h�#/��ٿ��f�#�@�+�ۢ4@=�;o��!?!���@h�#/��ٿ��f�#�@�+�ۢ4@=�;o��!?!���@c}�.�ٿ�	�W��@�O#�4@�0��d�!?������@��H�j�ٿ�k�#8�@vK����3@Y㺠�!?G��M�@��H�j�ٿ�k�#8�@vK����3@Y㺠�!?G��M�@��H�j�ٿ�k�#8�@vK����3@Y㺠�!?G��M�@��H�j�ٿ�k�#8�@vK����3@Y㺠�!?G��M�@�&	�ٿ���a���@;]J�'�3@��D��!?&�)���@�����ٿ40^��@D��OQ�3@�zgB�!?i�� Ե@�����ٿ40^��@D��OQ�3@�zgB�!?i�� Ե@�����ٿ40^��@D��OQ�3@�zgB�!?i�� Ե@�����ٿ40^��@D��OQ�3@�zgB�!?i�� Ե@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@"l��ٿmZ���G�@�����3@�Lݩ�!?/f�7o�@�2m�{�ٿm@�D��@Wg��3@���(i�!?bL�:��@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@0��B�ٿ4�5쒫�@�`b�4�3@'�B6b�!?�S�Ǹz�@�|���ٿ�5"��@B��|4@�-47�!?fA�/G�@�|���ٿ�5"��@B��|4@�-47�!?fA�/G�@Co�/��ٿ�[��A�@�g���3@�!?w<����@�_� �ٿ7����@��BI��3@B�#�!?�ŝ��s�@�_� �ٿ7����@��BI��3@B�#�!?�ŝ��s�@�_� �ٿ7����@��BI��3@B�#�!?�ŝ��s�@�8� ��ٿ ��6���@�K�%��3@����M�!?x7���@�8� ��ٿ ��6���@�K�%��3@����M�!?x7���@��#�ٿO���J�@U
��3@z�zrm�!??4�~��@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@�`�
�ٿ]������@�QL.�3@�^([��!?o��`���@Z1�N�ٿ�D*�X,�@������3@�_��_�!?�t¥��@C��-�ٿ�������@����3@N�1�D�!?�l���j�@=8��ɛٿ�&݈��@�ट��3@|s�X�!?�0�
ߴ@=8��ɛٿ�&݈��@�ट��3@|s�X�!?�0�
ߴ@=8��ɛٿ�&݈��@�ट��3@|s�X�!?�0�
ߴ@=8��ɛٿ�&݈��@�ट��3@|s�X�!?�0�
ߴ@=8��ɛٿ�&݈��@�ट��3@|s�X�!?�0�
ߴ@&5~i�ٿ�	��� �@��W6��3@��s�!?�x!�9��@&5~i�ٿ�	��� �@��W6��3@��s�!?�x!�9��@��inr�ٿ�Ya��a�@������3@6b:_8�!?��e�z�@��inr�ٿ�Ya��a�@������3@6b:_8�!?��e�z�@��inr�ٿ�Ya��a�@������3@6b:_8�!?��e�z�@��inr�ٿ�Ya��a�@������3@6b:_8�!?��e�z�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@���J�ٿ�NN����@�޹���3@�P\�)�!?��m|�O�@�TT��ٿ�#���@�G�`4@!�.�L�!?m�*�@9�����ٿ=M��-��@;��u�3@}�;,f�!?V$(��@9�����ٿ=M��-��@;��u�3@}�;,f�!?V$(��@9�����ٿ=M��-��@;��u�3@}�;,f�!?V$(��@��)HM�ٿ1���q��@Tc���3@6E�i�!?o9��h�@�iD�Бٿ�"߂��@���8X�3@���gc�!?jii:�M�@�iD�Бٿ�"߂��@���8X�3@���gc�!?jii:�M�@�iD�Бٿ�"߂��@���8X�3@���gc�!?jii:�M�@�<5�ٿ��2bhO�@��ǫK�3@�,��!?p��J/�@1���Țٿ��N����@�-����3@B���!?0W5h0��@P�o�ٿo5�;�@�����3@e�Y���!?4Bo���@������ٿ�ML����@G��q��3@	����!?��F�7��@���=�ٿ/�&��f�@�|jk�3@�G��v�!?�N�<ʹ@���=�ٿ/�&��f�@�|jk�3@�G��v�!?�N�<ʹ@<]P��ٿ&eEa��@>Y���3@�B.�!?�>��Y�@<]P��ٿ&eEa��@>Y���3@�B.�!?�>��Y�@��ѕ�ٿ����O��@����3@[��i�!?�IF�U9�@��ѕ�ٿ����O��@����3@[��i�!?�IF�U9�@l��m�ٿ�Oo���@��Ÿ�3@@x�
�!?�_%��@l��m�ٿ�Oo���@��Ÿ�3@@x�
�!?�_%��@l��m�ٿ�Oo���@��Ÿ�3@@x�
�!?�_%��@l��m�ٿ�Oo���@��Ÿ�3@@x�
�!?�_%��@ݮ!n�ٿk�W�@T6a:�3@)ܰ,N�!?�gJ��f�@ݮ!n�ٿk�W�@T6a:�3@)ܰ,N�!?�gJ��f�@ݮ!n�ٿk�W�@T6a:�3@)ܰ,N�!?�gJ��f�@ݮ!n�ٿk�W�@T6a:�3@)ܰ,N�!?�gJ��f�@�vМ�ٿ$~�#Ai�@��Ť��3@Ij��*�!?���TK�@�vМ�ٿ$~�#Ai�@��Ť��3@Ij��*�!?���TK�@����ٿ�#>����@qQ����3@8�]./�!?��E<`@�@����ٿ�#>����@qQ����3@8�]./�!?��E<`@�@����ٿ�#>����@qQ����3@8�]./�!?��E<`@�@����ٿ�#>����@qQ����3@8�]./�!?��E<`@�@���>��ٿ >�Ϋ=�@�7��M�3@˒f�!?S�&�6�@���>��ٿ >�Ϋ=�@�7��M�3@˒f�!?S�&�6�@���>��ٿ >�Ϋ=�@�7��M�3@˒f�!?S�&�6�@T����ٿ쌿���@����3@�2�Dm�!?W<L�o"�@T����ٿ쌿���@����3@�2�Dm�!?W<L�o"�@ZP��ٿg��
��@,`Hbc�3@;�<h�!?.%���@ZP��ٿg��
��@,`Hbc�3@;�<h�!?.%���@ZP��ٿg��
��@,`Hbc�3@;�<h�!?.%���@���}��ٿ��C�W��@u�V~o�3@�d*�!?��o逌�@���}��ٿ��C�W��@u�V~o�3@�d*�!?��o逌�@7�q�&�ٿ�:)lEZ�@�=J��3@5�7�/�!?�j�9PD�@f��k��ٿ8*�X��@_5���3@RT�]�!?u�$t�@f��k��ٿ8*�X��@_5���3@RT�]�!?u�$t�@f��k��ٿ8*�X��@_5���3@RT�]�!?u�$t�@��[˕ٿ��J3��@ҿ�Ȉ�3@~A�E�!?��z��@��[˕ٿ��J3��@ҿ�Ȉ�3@~A�E�!?��z��@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@q�k�ٿr���Z�@|��>��3@hJ����!?I�2	���@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@8��L�ٿ9F�<�@�KN���3@&��C�!?�B�F�µ@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@�,��|�ٿ��?���@�Z4�A�3@Z4�!?Ր��M��@H����ٿ�!|��@
{�z�3@���X$�!?�Id��@H����ٿ�!|��@
{�z�3@���X$�!?�Id��@���ٿ��GRm"�@En5\�3@�����!?K����@���ٿ��GRm"�@En5\�3@�����!?K����@���ٿ��GRm"�@En5\�3@�����!?K����@���ٿ��GRm"�@En5\�3@�����!?K����@���ٿ��GRm"�@En5\�3@�����!?K����@���ٿ��GRm"�@En5\�3@�����!?K����@Y��֑ٿ%t�/��@�Ņ���3@�@E�!?Y���N��@+:>�ٿmC!� �@�S��3@��J7*�!?
��i|�@�����ٿ(ۆ�I��@�1��3@�qLy�!?�l���@�����ٿ(ۆ�I��@�1��3@�qLy�!?�l���@�����ٿ(ۆ�I��@�1��3@�qLy�!?�l���@�~|��ٿF�j���@�z����3@c��t|�!?�]�,�@�~|��ٿF�j���@�z����3@c��t|�!?�]�,�@�~|��ٿF�j���@�z����3@c��t|�!?�]�,�@�~|��ٿF�j���@�z����3@c��t|�!?�]�,�@������ٿ'����@Z��6�	4@2#W�y�!?���_�@U�|��ٿ���m���@ţ�E4@��.�&�!?+O:
K��@U�|��ٿ���m���@ţ�E4@��.�&�!?+O:
K��@
)�㡕ٿm�MXc�@�(`A4@;8_��!?�C)H��@
)�㡕ٿm�MXc�@�(`A4@;8_��!?�C)H��@
)�㡕ٿm�MXc�@�(`A4@;8_��!?�C)H��@�8�L�ٿ��K)Kg�@�u�u"	4@���8��!?9~��@�8�L�ٿ��K)Kg�@�u�u"	4@���8��!?9~��@ɼO�ٿ������@Ҍ��F�3@��9��!?��0+U�@ɼO�ٿ������@Ҍ��F�3@��9��!?��0+U�@ɼO�ٿ������@Ҍ��F�3@��9��!?��0+U�@������ٿ�yS�e��@��a��3@��z�^�!?ėK��q�@������ٿ�yS�e��@��a��3@��z�^�!?ėK��q�@������ٿ�yS�e��@��a��3@��z�^�!?ėK��q�@������ٿ�yS�e��@��a��3@��z�^�!?ėK��q�@A�y�ٿm	�Y�&�@����3@4G��d�!?f�_�@j�5$�ٿ������@��LP��3@=���!?�ԨC�@j�5$�ٿ������@��LP��3@=���!?�ԨC�@j�5$�ٿ������@��LP��3@=���!?�ԨC�@Pu��~�ٿ�4HX�@�^(�4@IE򟻐!?��.8�@p2w�b�ٿQ��s_�@ ��g�3@�����!?M��%���@�}Eԉ�ٿ嶦ہ$�@�[K��3@���%��!?��aȊn�@�}Eԉ�ٿ嶦ہ$�@�[K��3@���%��!?��aȊn�@�AX��ٿ-saw���@��O�4@M��ѐ!?��;��@�AX��ٿ-saw���@��O�4@M��ѐ!?��;��@
0;$>�ٿ��O%�G�@�h)�3@)Pv��!?����iT�@
0;$>�ٿ��O%�G�@�h)�3@)Pv��!?����iT�@
0;$>�ٿ��O%�G�@�h)�3@)Pv��!?����iT�@
0;$>�ٿ��O%�G�@�h)�3@)Pv��!?����iT�@
0;$>�ٿ��O%�G�@�h)�3@)Pv��!?����iT�@���x��ٿO�_����@�T
K��3@_j6��!?ZG�2�@���x��ٿO�_����@�T
K��3@_j6��!?ZG�2�@���x��ٿO�_����@�T
K��3@_j6��!?ZG�2�@��:�ҝٿ�4��Rk�@�+'�x�3@ŀ�!?Y��/��@��:�ҝٿ�4��Rk�@�+'�x�3@ŀ�!?Y��/��@��:�ҝٿ�4��Rk�@�+'�x�3@ŀ�!?Y��/��@��:�ҝٿ�4��Rk�@�+'�x�3@ŀ�!?Y��/��@��:�ҝٿ�4��Rk�@�+'�x�3@ŀ�!?Y��/��@r�{��ٿ���q�@�a�6�3@K�Z�!?���Z���@r�{��ٿ���q�@�a�6�3@K�Z�!?���Z���@r�{��ٿ���q�@�a�6�3@K�Z�!?���Z���@r�{��ٿ���q�@�a�6�3@K�Z�!?���Z���@r�{��ٿ���q�@�a�6�3@K�Z�!?���Z���@n�Z�}�ٿͼ�d��@���9�3@s���!?�e���)�@n�Z�}�ٿͼ�d��@���9�3@s���!?�e���)�@�
�F�ٿ+^���@UA��8�3@�g��!?���Tv�@�
�F�ٿ+^���@UA��8�3@�g��!?���Tv�@�
�F�ٿ+^���@UA��8�3@�g��!?���Tv�@�
�F�ٿ+^���@UA��8�3@�g��!?���Tv�@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@�M��f�ٿYB7��@�����3@���3�!?��~��@f;����ٿc^n����@�����3@*�(�!?Ȟ3h��@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@у���ٿ��>���@. | ��3@@<z5�!?�6z�G�@��躞ٿ�e���@]W'"p�3@u��%�!?y�g���@��躞ٿ�e���@]W'"p�3@u��%�!?y�g���@��躞ٿ�e���@]W'"p�3@u��%�!?y�g���@��u���ٿ�9.H��@E�
t_�3@zo��!?X�x�)�@��u���ٿ�9.H��@E�
t_�3@zo��!?X�x�)�@��u���ٿ�9.H��@E�
t_�3@zo��!?X�x�)�@��u���ٿ�9.H��@E�
t_�3@zo��!?X�x�)�@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@/lIq�ٿ�{4���@�N� v�3@X@k�f�!?m�Mb���@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��4J�ٿ�v�x0T�@K����3@��G�b�!?����@��o�Ϙٿ��(��
�@��G�/�3@±mb��!?rO��:յ@��o�Ϙٿ��(��
�@��G�/�3@±mb��!?rO��:յ@��o�Ϙٿ��(��
�@��G�/�3@±mb��!?rO��:յ@E\�I�ٿF���@|����3@	�/��!?����@E\�I�ٿF���@|����3@	�/��!?����@E\�I�ٿF���@|����3@	�/��!?����@E\�I�ٿF���@|����3@	�/��!?����@E\�I�ٿF���@|����3@	�/��!?����@E\�I�ٿF���@|����3@	�/��!?����@元l	�ٿ�L��!�@���h��3@����n�!?SP.d�@元l	�ٿ�L��!�@���h��3@����n�!?SP.d�@元l	�ٿ�L��!�@���h��3@����n�!?SP.d�@元l	�ٿ�L��!�@���h��3@����n�!?SP.d�@元l	�ٿ�L��!�@���h��3@����n�!?SP.d�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�;2Кٿ�.~�>��@GC��3@_,���!?�2�	�@�\�[J�ٿ%�=�D�@��ڟ�3@������!?��~O �@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@���HW�ٿ%�i֦b�@���q��3@��=]��!?��H��Z�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@2a�;ٝٿ�O�����@\�>�4@�gbh>�!?#
ad�@���D�ٿh�D�~�@�K5$�3@�	�,�!?b�w�@���D�ٿh�D�~�@�K5$�3@�	�,�!?b�w�@���D�ٿh�D�~�@�K5$�3@�	�,�!?b�w�@���D�ٿh�D�~�@�K5$�3@�	�,�!?b�w�@���D�ٿh�D�~�@�K5$�3@�	�,�!?b�w�@�`���ٿo��FQ��@U�9�r�3@��Y�܏!?�U��v�@�`���ٿo��FQ��@U�9�r�3@��Y�܏!?�U��v�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@���
�ٿ��^�;K�@"�
4@봾4v�!?�r�@�j�@:�2�ٿ��b��@�,�a�3@��1d�!?&x3��@:�2�ٿ��b��@�,�a�3@��1d�!?&x3��@�	C�B�ٿK�։��@-���3@`f(�K�!?�w�i$ӵ@�	C�B�ٿK�։��@-���3@`f(�K�!?�w�i$ӵ@�	C�B�ٿK�։��@-���3@`f(�K�!?�w�i$ӵ@ �ʫ�ٿ�s�~���@�Ei��3@%Ͽ�q�!?�Cs�x�@ �ʫ�ٿ�s�~���@�Ei��3@%Ͽ�q�!?�Cs�x�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@�ٿ�AF�ه�@ir���3@v��5��!?$XkP~l�@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@o���s�ٿr�ّ��@I��oJ�3@`��|T�!?� ���ص@>�ͬB�ٿ��KW=w�@���3@(8�O9�!?�Y�ϵ@g$q'��ٿ�V;�g�@|	6z�4@M·�M�!?�|K��r�@g$q'��ٿ�V;�g�@|	6z�4@M·�M�!?�|K��r�@g$q'��ٿ�V;�g�@|	6z�4@M·�M�!?�|K��r�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@�[��ٿLDp��r�@N)MJ�3@�Ċ?w�!?�nA�w�@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��Z)��ٿ?3�o�(�@*�Nh�4@�*�(��!?S\daAĴ@��T�ٿҕm
�u�@�/�x��3@+1��ߏ!?�����ô@��T�ٿҕm
�u�@�/�x��3@+1��ߏ!?�����ô@��T�ٿҕm
�u�@�/�x��3@+1��ߏ!?�����ô@��T�ٿҕm
�u�@�/�x��3@+1��ߏ!?�����ô@"�5¥�ٿ��W��@����H�3@�9qc��!?8B�靾�@"�5¥�ٿ��W��@����H�3@�9qc��!?8B�靾�@"�5¥�ٿ��W��@����H�3@�9qc��!?8B�靾�@"�5¥�ٿ��W��@����H�3@�9qc��!?8B�靾�@�*Z�'�ٿ��[���@��/�3@h�?���!?3}��Y��@Nw5_��ٿ���7���@��>\��3@�+��!?���!��@Nw5_��ٿ���7���@��>\��3@�+��!?���!��@Nw5_��ٿ���7���@��>\��3@�+��!?���!��@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@ �q�ٿ{d�D�A�@�����3@Lɛ�!?�a^fcz�@��qR��ٿv���Yƿ@4b<2�3@�aM+�!?�&%�%�@��qR��ٿv���Yƿ@4b<2�3@�aM+�!?�&%�%�@��qR��ٿv���Yƿ@4b<2�3@�aM+�!?�&%�%�@��qR��ٿv���Yƿ@4b<2�3@�aM+�!?�&%�%�@��qR��ٿv���Yƿ@4b<2�3@�aM+�!?�&%�%�@�,[��ٿ�qg�@�+7��3@���h��!?�D1���@�,[��ٿ�qg�@�+7��3@���h��!?�D1���@c�+�ٿI�>5Y$�@�X�w�3@6��,ِ!?���@�@c�+�ٿI�>5Y$�@�X�w�3@6��,ِ!?���@�@˫����ٿ������@#�����3@m)�jې!?r��⻵@'��)Əٿ���kc��@3��3@��'��!?��K���@'��)Əٿ���kc��@3��3@��'��!?��K���@'��)Əٿ���kc��@3��3@��'��!?��K���@'��)Əٿ���kc��@3��3@��'��!?��K���@'��)Əٿ���kc��@3��3@��'��!?��K���@����ٿ3��l{n�@)��w��3@����!?����n�@����ٿ3��l{n�@)��w��3@����!?����n�@����ٿ3��l{n�@)��w��3@����!?����n�@����ٿ3��l{n�@)��w��3@����!?����n�@����ٿ3��l{n�@)��w��3@����!?����n�@G��D�ٿs.^�KF�@�����3@V�z���!?��\���@9�r�K�ٿ.�>�f�@�k�J4@~Bqz�!?�p=҃�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@{l�F�ٿ�1��v��@ђ�EX4@}��&��!?�鿙\N�@c�9�ٿ��ڝ���@ �4�3@ɝ�=�!?eaT��w�@c�9�ٿ��ڝ���@ �4�3@ɝ�=�!?eaT��w�@c�9�ٿ��ڝ���@ �4�3@ɝ�=�!?eaT��w�@c�9�ٿ��ڝ���@ �4�3@ɝ�=�!?eaT��w�@pI��ٿ2���g�@d�/�@�3@���+[�!?D��{��@�![k��ٿ�E���@���f��3@���:�!?������@�![k��ٿ�E���@���f��3@���:�!?������@�~���ٿ��PXg��@bлC��3@�����!?L�e}�@Lu����ٿ �'�q\�@�o�˸�3@8��y'�!?�����@Lu����ٿ �'�q\�@�o�˸�3@8��y'�!?�����@O�Z��ٿD�AV��@�]�n��3@�e��&�!?�qc��@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@��q"�ٿ/N߯O�@�ti��3@�{=�!?uNH�۴@���o�ٿ[|�|��@������3@����׏!?�b�Gȴ@?Ʌ5�ٿ��� ���@���:�3@�Xx-�!?����z�@?Ʌ5�ٿ��� ���@���:�3@�Xx-�!?����z�@?Ʌ5�ٿ��� ���@���:�3@�Xx-�!?����z�@?Ʌ5�ٿ��� ���@���:�3@�Xx-�!?����z�@�i���ٿ�����@��F4@���T��!?�xo]��@�i���ٿ�����@��F4@���T��!?�xo]��@�i���ٿ�����@��F4@���T��!?�xo]��@H"2U�ٿn��7(��@.��>�4@�&$�!?+�'#ʴ@KD�֔ٿ��_,k�@�R�^�3@$'9y�!?��o^��@KD�֔ٿ��_,k�@�R�^�3@$'9y�!?��o^��@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@݅��ɏٿ�]Y�4��@QC���3@ai�l�!?L�'K�@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@w\�ٿ�3pQ(�@���3@ͦ!�w�!?�4�p��@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��6(�ٿ����@g��g�3@������!?��
v�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@��pR�ٿb�SX�O�@�����3@�R����!?�$ڞ�6�@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@�z�ڢ�ٿ�=�G��@#��u��3@J0Z7�!?�b�����@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@���,G�ٿ�\��v�@#�O�!�3@L>�@�!?�[��f>�@�Y�G�ٿ��=9���@�ڳF~�3@�b�3�!?Y�wvĲ�@�Y�G�ٿ��=9���@�ڳF~�3@�b�3�!?Y�wvĲ�@j'q�ۛٿ�����@�6�e?�3@�-�4�!?AJ�e��@j'q�ۛٿ�����@�6�e?�3@�-�4�!?AJ�e��@j'q�ۛٿ�����@�6�e?�3@�-�4�!?AJ�e��@j'q�ۛٿ�����@�6�e?�3@�-�4�!?AJ�e��@�Գ&��ٿ��8=�@�LmO�3@��]�n�!?H��Հ�@�Գ&��ٿ��8=�@�LmO�3@��]�n�!?H��Հ�@�Գ&��ٿ��8=�@�LmO�3@��]�n�!?H��Հ�@�Գ&��ٿ��8=�@�LmO�3@��]�n�!?H��Հ�@��7ן�ٿ{NCG��@v6ȣv�3@���6Z�!?����ڵ@��7ן�ٿ{NCG��@v6ȣv�3@���6Z�!?����ڵ@M�y�@�ٿU�ѯ�@{K�3@ҩ~�!?�Ia���@M�y�@�ٿU�ѯ�@{K�3@ҩ~�!?�Ia���@Dt�`��ٿ��@�!�@�j��3@���N`�!?a �k޵@Dt�`��ٿ��@�!�@�j��3@���N`�!?a �k޵@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@��Ԃ�ٿ��WZP�@�����3@²k+��!?if����@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@D�~w��ٿN� �@����3@oD��Z�!?{�d��W�@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�6Qƙٿ-�->�V�@�o�Y�3@��q�!?���.6޴@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@�e+�ٿ��eQb�@6�����3@^	:��!?=۳�kW�@I���ٿ̞+�g�@�
څ��3@80����!?�yd��q�@I���ٿ̞+�g�@�
څ��3@80����!?�yd��q�@I���ٿ̞+�g�@�
څ��3@80����!?�yd��q�@I���ٿ̞+�g�@�
څ��3@80����!?�yd��q�@��9l�ٿx2�7�+�@��	�B4@j� |�!?"����@��9l�ٿx2�7�+�@��	�B4@j� |�!?"����@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�eI���ٿ���s��@���q4@jZ�M��!?*`N��@�%|�Z�ٿ�	)�@��V�3@
�a"Ȑ!?lƐy��@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@u����ٿ�{f���@���l��3@��-��!?}N����@�y�(>�ٿ+�`
���@�g��3@-��@�!?��6 ��@�y�(>�ٿ+�`
���@�g��3@-��@�!?��6 ��@�H3�&�ٿZ��h��@&^k���3@\�|}�!?z��	���@�H3�&�ٿZ��h��@&^k���3@\�|}�!?z��	���@�H3�&�ٿZ��h��@&^k���3@\�|}�!?z��	���@�H3�&�ٿZ��h��@&^k���3@\�|}�!?z��	���@�H3�&�ٿZ��h��@&^k���3@\�|}�!?z��	���@	��ٿ��)1W�@���>C�3@B�{���!?j)|���@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@s�ȧɜٿ�
����@�7��}4@���!?!<�� �@	^6��ٿb�ư��@Y�lf4@� F�!?��0e���@	^6��ٿb�ư��@Y�lf4@� F�!?��0e���@;�y��ٿ2��qCd�@�k���4@��g�0�!?���N�@;�y��ٿ2��qCd�@�k���4@��g�0�!?���N�@;�y��ٿ2��qCd�@�k���4@��g�0�!?���N�@{q�͒ٿ����!��@q��^�3@E�7��!?Na���@{q�͒ٿ����!��@q��^�3@E�7��!?Na���@�@�;��ٿåTkCX�@7��v��3@�P:�!?lV�Ul�@�@�;��ٿåTkCX�@7��v��3@�P:�!?lV�Ul�@�@�;��ٿåTkCX�@7��v��3@�P:�!?lV�Ul�@�@�;��ٿåTkCX�@7��v��3@�P:�!?lV�Ul�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@�x�R��ٿ���ς��@������3@
U��B�!?��ʢ(�@���� �ٿ��d˘�@�!�V�3@�E�ޑ�!?1:ɕҪ�@���� �ٿ��d˘�@�!�V�3@�E�ޑ�!?1:ɕҪ�@���� �ٿ��d˘�@�!�V�3@�E�ޑ�!?1:ɕҪ�@���� �ٿ��d˘�@�!�V�3@�E�ޑ�!?1:ɕҪ�@�:&\�ٿt�h=��@��Y�3@�;.[��!?d��^���@�:&\�ٿt�h=��@��Y�3@�;.[��!?d��^���@6H��W�ٿ"�r���@���f��3@h��!?�*R���@6H��W�ٿ"�r���@���f��3@h��!?�*R���@�N�]��ٿ�т(-��@�����3@Y�H�!?�	e���@�����ٿ@;ZR�@]��C�3@�(�\/�!?����R�@�����ٿ@;ZR�@]��C�3@�(�\/�!?����R�@�����ٿ@;ZR�@]��C�3@�(�\/�!?����R�@�����ٿ@;ZR�@]��C�3@�(�\/�!?����R�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@5���ٿ��%��@ΛW��	4@�U`���!?�ƧiZ�@�L�ٿ֝r+-�@��X��3@�g�F��!?z\�H���@�L�ٿ֝r+-�@��X��3@�g�F��!?z\�H���@{`m�\�ٿ/Wæ�@.u��3@�-�ҏ!?[/�5"�@{`m�\�ٿ/Wæ�@.u��3@�-�ҏ!?[/�5"�@{`m�\�ٿ/Wæ�@.u��3@�-�ҏ!?[/�5"�@FU�H�ٿ���>�@��Fu��3@h���!?�Հ��r�@FU�H�ٿ���>�@��Fu��3@h���!?�Հ��r�@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@����ٿ�f;�'�@^C�E�3@Ȳ'��!?�G�$cʹ@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@��'��ٿj<\��H�@����(�3@�s��U�!?�X�c뤵@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@˿���ٿkٍB�@�����3@�� �^�!?)�-6t�@�
�RǙٿ����@��&��3@ڿxB�!?��:P���@��5C�ٿ!�����@=�$s��3@��
�!?"Z��v�@��5C�ٿ!�����@=�$s��3@��
�!?"Z��v�@��5C�ٿ!�����@=�$s��3@��
�!?"Z��v�@��5C�ٿ!�����@=�$s��3@��
�!?"Z��v�@��5C�ٿ!�����@=�$s��3@��
�!?"Z��v�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@�l���ٿ�C�2�(�@�ɉF�3@�+�@�!?d75�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@��Os�ٿdu���a�@#�v�2�3@*H�PX�!?L���՝�@'�Rؗٿ��i�&�@����4@"�Qa�!?�p��^�@'�Rؗٿ��i�&�@����4@"�Qa�!?�p��^�@'�Rؗٿ��i�&�@����4@"�Qa�!?�p��^�@'�Rؗٿ��i�&�@����4@"�Qa�!?�p��^�@'�Rؗٿ��i�&�@����4@"�Qa�!?�p��^�@O�Och�ٿ�����@gǡ5�4@ ��에!?u�7�a�@O�Och�ٿ�����@gǡ5�4@ ��에!?u�7�a�@O�Och�ٿ�����@gǡ5�4@ ��에!?u�7�a�@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@��c�ٿ8^�;�m�@l\K��3@C$F�9�!?���	��@ƶz8��ٿe�KP+�@5�Xo4@h��J�!?�-s��@S����ٿ�����@l�vx3�3@܀&�Z�!?rc���*�@S����ٿ�����@l�vx3�3@܀&�Z�!?rc���*�@S����ٿ�����@l�vx3�3@܀&�Z�!?rc���*�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@�l(V8�ٿ�t�<��@��HK�3@,훉�!?��C�M�@4S~���ٿ�Q� �q�@�"2-��3@�}�tp�!?���!)�@�M��ٿ�?\( �@�;�&��3@����%�!?%tQ�C��@_����ٿ	�"�I�@�W �3@�gO5_�!?�0�He��@_����ٿ	�"�I�@�W �3@�gO5_�!?�0�He��@_����ٿ	�"�I�@�W �3@�gO5_�!?�0�He��@_����ٿ	�"�I�@�W �3@�gO5_�!?�0�He��@_����ٿ	�"�I�@�W �3@�gO5_�!?�0�He��@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@��ZɆ�ٿO�:�v�@�e!`��3@*݀=)�!?���A!̵@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@�����ٿ�X����@Vpj�3@�L�!�!?�d��B@�@��?��ٿ��yW��@_?Φe�3@<f,P��!?�^�,>M�@W����ٿ�x}�i��@ÔM��3@��*�8�!?��*��@W����ٿ�x}�i��@ÔM��3@��*�8�!?��*��@W����ٿ�x}�i��@ÔM��3@��*�8�!?��*��@W����ٿ�x}�i��@ÔM��3@��*�8�!?��*��@�����ٿ�I�����@?`q3]4@a| [X�!?�l�j�@�����ٿ=l��/��@n�ܾX�3@�w�!?�[a�@�����ٿ=l��/��@n�ܾX�3@�w�!?�[a�@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@
�A�ٿ��׳ݭ�@�*�}�3@ظ9�*�!?>P�����@�^}���ٿ �*&���@�dD�3@�i�A�!?��9�T�@�^}���ٿ �*&���@�dD�3@�i�A�!?��9�T�@r����ٿg5\z�b�@ �z��3@C9��!?��יtȴ@r����ٿg5\z�b�@ �z��3@C9��!?��יtȴ@r����ٿg5\z�b�@ �z��3@C9��!?��יtȴ@r����ٿg5\z�b�@ �z��3@C9��!?��יtȴ@6P>t{�ٿ��%ë��@�H��3@vCS{(�!?����Zǵ@6P>t{�ٿ��%ë��@�H��3@vCS{(�!?����Zǵ@m\M��ٿ�*.Lt�@��o���3@�_I�$�!?I��ω��@m\M��ٿ�*.Lt�@��o���3@�_I�$�!?I��ω��@m\M��ٿ�*.Lt�@��o���3@�_I�$�!?I��ω��@�!�	Θٿ@l�(E��@��۸�3@�]n�!?,��t(ȴ@�!�	Θٿ@l�(E��@��۸�3@�]n�!?,��t(ȴ@�!�	Θٿ@l�(E��@��۸�3@�]n�!?,��t(ȴ@�!�	Θٿ@l�(E��@��۸�3@�]n�!?,��t(ȴ@S�/N�ٿa�y���@���u�3@�����!?�ju�n��@g���-�ٿG�� a��@Uq���3@�Ow�!?�eMg!
�@N��1�ٿℰx��@�[-�'�3@�����!?��s��@N��1�ٿℰx��@�[-�'�3@�����!?��s��@N��1�ٿℰx��@�[-�'�3@�����!?��s��@]4�b�ٿ�S���@x^�F��3@yi%D�!?�.&@̴@]4�b�ٿ�S���@x^�F��3@yi%D�!?�.&@̴@]4�b�ٿ�S���@x^�F��3@yi%D�!?�.&@̴@�B���ٿ���@�}`���3@�ۤwy�!?�l?4���@�B���ٿ���@�}`���3@�ۤwy�!?�l?4���@�f��ٿ�u{��e�@�J���3@Y���`�!?i�i!���@�f��ٿ�u{��e�@�J���3@Y���`�!?i�i!���@dj�(�ٿhk~���@������3@􏐥]�!?x!0�\ �@dj�(�ٿhk~���@������3@􏐥]�!?x!0�\ �@dj�(�ٿhk~���@������3@􏐥]�!?x!0�\ �@dj�(�ٿhk~���@������3@􏐥]�!?x!0�\ �@dj�(�ٿhk~���@������3@􏐥]�!?x!0�\ �@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@���ɖٿyk|�;�@�I+���3@�@HJ��!?b���i�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@I�>�ٿ�h�h(��@v��r��3@.��q=�!?n��l�N�@�.��Y�ٿ`��	>��@�]!���3@`nO�!?��F�lմ@�.��Y�ٿ`��	>��@�]!���3@`nO�!?��F�lմ@�.��Y�ٿ`��	>��@�]!���3@`nO�!?��F�lմ@|.H=:�ٿE�&V� �@����3@�R��!?�>�9C�@|.H=:�ٿE�&V� �@����3@�R��!?�>�9C�@|.H=:�ٿE�&V� �@����3@�R��!?�>�9C�@|.H=:�ٿE�&V� �@����3@�R��!?�>�9C�@juG�
�ٿ��{h[��@�y&��3@>�A�Ð!?D��-z�@juG�
�ٿ��{h[��@�y&��3@>�A�Ð!?D��-z�@߲�b��ٿ�E�CP��@��|�L�3@0����!?��W5o�@߲�b��ٿ�E�CP��@��|�L�3@0����!?��W5o�@߲�b��ٿ�E�CP��@��|�L�3@0����!?��W5o�@߲�b��ٿ�E�CP��@��|�L�3@0����!?��W5o�@y���y�ٿ2����@s�4@z&��!?���}�@y���y�ٿ2����@s�4@z&��!?���}�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@%7Q�i�ٿ�׷���@�P� 4@�F� `�!?�5�UM�@����c�ٿ��Lx���@���%��3@�RP�!?ܡ���8�@�w#�ٿ�`m��A�@j���3@s�����!?���|��@�w#�ٿ�`m��A�@j���3@s�����!?���|��@�w#�ٿ�`m��A�@j���3@s�����!?���|��@�w#�ٿ�`m��A�@j���3@s�����!?���|��@�w#�ٿ�`m��A�@j���3@s�����!?���|��@,��7�ٿF�;��@}�:�4@��,F��!?�yHf&m�@,��7�ٿF�;��@}�:�4@��,F��!?�yHf&m�@,��7�ٿF�;��@}�:�4@��,F��!?�yHf&m�@,��7�ٿF�;��@}�:�4@��,F��!?�yHf&m�@�Xnѹ�ٿ;�k]���@��)���3@��!?�����w�@�Xnѹ�ٿ;�k]���@��)���3@��!?�����w�@�Xnѹ�ٿ;�k]���@��)���3@��!?�����w�@���H�ٿ���̹�@�\`
�4@�d��'�!?`�ۈ�Ӵ@���H�ٿ���̹�@�\`
�4@�d��'�!?`�ۈ�Ӵ@���H�ٿ���̹�@�\`
�4@�d��'�!?`�ۈ�Ӵ@���H�ٿ���̹�@�\`
�4@�d��'�!?`�ۈ�Ӵ@���H�ٿ���̹�@�\`
�4@�d��'�!?`�ۈ�Ӵ@K��н�ٿ�eȮ���@4�\P�3@�L��|�!?dC���@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@xWLq$�ٿf���e�@�=_( 4@�>�u2�!?�VC�,�@\~r_�ٿ�$[�@�t\��3@Q!��!?i~N���@��xҏ�ٿ����a�@64@���3@a���ŏ!?�Ս�ô@��xҏ�ٿ����a�@64@���3@a���ŏ!?�Ս�ô@��xҏ�ٿ����a�@64@���3@a���ŏ!?�Ս�ô@{�>F��ٿ)P�6�@yHEm��3@��3�Ϗ!?�����˴@{�>F��ٿ)P�6�@yHEm��3@��3�Ϗ!?�����˴@�&�0�ٿ+����@v�3@t��&(�!?Y�xW#�@�&�0�ٿ+����@v�3@t��&(�!?Y�xW#�@�&�0�ٿ+����@v�3@t��&(�!?Y�xW#�@�&�0�ٿ+����@v�3@t��&(�!?Y�xW#�@���1Ȕٿm#1��t�@���X�3@<޶A�!?��.��@���1Ȕٿm#1��t�@���X�3@<޶A�!?��.��@���1Ȕٿm#1��t�@���X�3@<޶A�!?��.��@����B�ٿ�t����@[����3@���!?p���^*�@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@h��ٿ�:"�}��@ �!�3@9���n�!?�.���ʹ@��Y|�ٿ�qW��_�@�!��3@:?�	&�!?4�{�@��Y|�ٿ�qW��_�@�!��3@:?�	&�!?4�{�@��Y|�ٿ�qW��_�@�!��3@:?�	&�!?4�{�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@X	Z�^�ٿ��~�-��@x�3Y�3@&>_�*�!?Q,��,�@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@�a���ٿ��F�D��@'p���4@$Nu煐!?�aa���@47d~��ٿȵi�F��@c��j��3@窥/B�!?a�+Cδ@47d~��ٿȵi�F��@c��j��3@窥/B�!?a�+Cδ@47d~��ٿȵi�F��@c��j��3@窥/B�!?a�+Cδ@47d~��ٿȵi�F��@c��j��3@窥/B�!?a�+Cδ@47d~��ٿȵi�F��@c��j��3@窥/B�!?a�+Cδ@���{Z�ٿ�������@����T�3@r���!?���n���@���{Z�ٿ�������@����T�3@r���!?���n���@���{Z�ٿ�������@����T�3@r���!?���n���@_��Z�ٿ��2GP�@��*Y`�3@7�(�!?axp/��@_��Z�ٿ��2GP�@��*Y`�3@7�(�!?axp/��@_��Z�ٿ��2GP�@��*Y`�3@7�(�!?axp/��@�Ĳ��ٿ�i_���@���͂�3@�t�]�!?S~�\��@�Ĳ��ٿ�i_���@���͂�3@�t�]�!?S~�\��@���I�ٿiR���e�@�n�Ġ�3@�a[�%�!?�^����@�F��(�ٿ�/�;9�@#,5�g�3@�9���!?~~	���@J�(��ٿ�f\/�@�{z�>�3@d�7�}�!?�=�d�!�@J�(��ٿ�f\/�@�{z�>�3@d�7�}�!?�=�d�!�@{(�}�ٿ��ǽ%��@GLh��3@M�_�X�!?p��9��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@�G�(�ٿ9�$H���@ߕ�C��3@0<	ɏ!?@�c�o��@> q��ٿ?%��Y��@��� �3@(4.���!?�r:)5�@> q��ٿ?%��Y��@��� �3@(4.���!?�r:)5�@> q��ٿ?%��Y��@��� �3@(4.���!?�r:)5�@���ٿ������@���M�3@�UB�/�!?�iy~N�@���ٿ������@���M�3@�UB�/�!?�iy~N�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@v®�ٿ����;�@�W��3@����I�!?"�F�O�@D���ٿ�~7U���@���H��3@��J�s�!?��Bp
�@��S�ٿ`2�d�@I�� l�3@wة���!?����"�@��S�ٿ`2�d�@I�� l�3@wة���!?����"�@v�z�ٿ�N�~~Z�@�O�sj�3@���!?�0oCF�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@'���ٿ���{No�@�$�	�3@�/��!?��eaA�@��j��ٿ㋖���@=-٥��3@���!?������@Kh�ٯ�ٿ�=��@-���4@�Z��V�!?n�1L#��@�J����ٿ�Oͧ��@���4@��'E�!?�R��Gj�@�J����ٿ�Oͧ��@���4@��'E�!?�R��Gj�@�J����ٿ�Oͧ��@���4@��'E�!?�R��Gj�@�J����ٿ�Oͧ��@���4@��'E�!?�R��Gj�@�p"g�ٿ�LC��X�@ ,T�R�3@גd��!?�l���ʹ@�p"g�ٿ�LC��X�@ ,T�R�3@גd��!?�l���ʹ@�p"g�ٿ�LC��X�@ ,T�R�3@גd��!?�l���ʹ@�p"g�ٿ�LC��X�@ ,T�R�3@גd��!?�l���ʹ@�p"g�ٿ�LC��X�@ ,T�R�3@גd��!?�l���ʹ@%���I�ٿ��ZV!�@��i���3@�u� ŏ!?yb�@��@%���I�ٿ��ZV!�@��i���3@�u� ŏ!?yb�@��@%���I�ٿ��ZV!�@��i���3@�u� ŏ!?yb�@��@���}�ٿ ��_��@�M�i��3@}{��!?J�iS�@>048@�ٿ� ?����@��1�3@��`��!?�y$�D�@>048@�ٿ� ?����@��1�3@��`��!?�y$�D�@O�%��ٿ�' �|�@)76��3@�t1�	�!?��{=��@O�%��ٿ�' �|�@)76��3@�t1�	�!?��{=��@O�%��ٿ�' �|�@)76��3@�t1�	�!?��{=��@sҤ��ٿ�f�KW�@�SX���3@H���!?Z�ۡ�@sҤ��ٿ�f�KW�@�SX���3@H���!?Z�ۡ�@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@b����ٿ��'C���@�����3@��c�!?|7�/���@��<R�ٿf�7�Cv�@J>̑�3@��EZ�!?U�ｴ@��<R�ٿf�7�Cv�@J>̑�3@��EZ�!?U�ｴ@��<R�ٿf�7�Cv�@J>̑�3@��EZ�!?U�ｴ@��<R�ٿf�7�Cv�@J>̑�3@��EZ�!?U�ｴ@��<R�ٿf�7�Cv�@J>̑�3@��EZ�!?U�ｴ@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@�m`�˚ٿpI�o��@��]LC�3@�ů�x�!?��C�O�@KG�%�ٿ�r�.i��@fV� ��3@�o��!?3�G�d$�@8�K��ٿ��g��h�@I'q�:�3@nI���!?�vm�ub�@8�K��ٿ��g��h�@I'q�:�3@nI���!?�vm�ub�@��& �ٿ-��Pb��@9���s4@�0���!?crob���@��& �ٿ-��Pb��@9���s4@�0���!?crob���@b9=��ٿ�FL�"]�@A��4@ϛ��y�!?e�Ӷ]�@Ss�Z�ٿAK��@��m��3@���@�!?�*���@Ss�Z�ٿAK��@��m��3@���@�!?�*���@Ss�Z�ٿAK��@��m��3@���@�!?�*���@Ss�Z�ٿAK��@��m��3@���@�!?�*���@Ss�Z�ٿAK��@��m��3@���@�!?�*���@Ss�Z�ٿAK��@��m��3@���@�!?�*���@�"J��ٿ�Q�Z���@��|��3@�'m���!?1N۠Wȴ@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@���O�ٿq_����@~%{y�3@3��(U�!?^�~��@g��c�ٿ�Rm��@�����3@T��o��!?a�G�-�@g��c�ٿ�Rm��@�����3@T��o��!?a�G�-�@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@=h�[H�ٿ�NLP�@�O�$K�3@�S-^@�!?[],��@��+�ٿ�ޚ�oo�@��@��3@��X��!?@��l��@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@�Sm��ٿ�X�(�Q�@�7��3@ ���M�!?�g+PK�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@d?��;�ٿa���y��@��c��3@Q�k�!?��:�L�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@���Nȕٿ�<��j��@�c��%�3@���C�!?�lS�4=�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@����ʔٿSu���R�@��S���3@^��T�!??m�vy|�@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@���衚ٿ<����@����3@�;l�N�!?VIrA�δ@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@�-5;�ٿ�.�nj��@|+����3@oS��-�!?KNQnH�@��9cM�ٿ�("���@ImR��3@f�a�7�!?*|�@��9cM�ٿ�("���@ImR��3@f�a�7�!?*|�@#vp�&�ٿ$;Jh�@�%��3@Fo�I�!?����@#vp�&�ٿ$;Jh�@�%��3@Fo�I�!?����@/s/&͕ٿ;�A<��@ż�h��3@���b�!?��444��@g�+H�ٿ��.v;�@S� N�3@mZ�e;�!?���M姵@g�+H�ٿ��.v;�@S� N�3@mZ�e;�!?���M姵@g�+H�ٿ��.v;�@S� N�3@mZ�e;�!?���M姵@�2���ٿ"���&��@��a�U�3@�g�=]�!?��b�D[�@�2���ٿ"���&��@��a�U�3@�g�=]�!?��b�D[�@�2���ٿ"���&��@��a�U�3@�g�=]�!?��b�D[�@��a!�ٿ�&����@s_���3@�'���!?l����ҵ@��a!�ٿ�&����@s_���3@�'���!?l����ҵ@��a!�ٿ�&����@s_���3@�'���!?l����ҵ@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@]�����ٿs��-��@��p&P�3@ci�)�!?AY[��@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@��Q}��ٿ�A��T��@^O���3@@�<�!?}��0�k�@W�3���ٿ�qו��@�v��\�3@�� �R�!?
� ��@W�3���ٿ�qו��@�v��\�3@�� �R�!?
� ��@W�3���ٿ�qו��@�v��\�3@�� �R�!?
� ��@W�3���ٿ�qו��@�v��\�3@�� �R�!?
� ��@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@�t_b�ٿ�= ��@D���o�3@���X�!?[�;3���@��Z�;�ٿ��{xo�@Q%��3@��O '�!?ѳ� ���@��Z�;�ٿ��{xo�@Q%��3@��O '�!?ѳ� ���@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@T��19�ٿٻ;��6�@��{��3@3.cޏ!?�x���w�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@^�%�y�ٿ�:N���@$G�>K�3@�a�!?�!1袡�@�����ٿ-ແ|�@s���3@��ӄT�!?���~�@
���ٿ�s�3��@򣁆��3@��O�!?I�y/`s�@
���ٿ�s�3��@򣁆��3@��O�!?I�y/`s�@>A���ٿ���o���@	*�4�3@SxUu�!?�K7�o��@>A���ٿ���o���@	*�4�3@SxUu�!?�K7�o��@>A���ٿ���o���@	*�4�3@SxUu�!?�K7�o��@>A���ٿ���o���@	*�4�3@SxUu�!?�K7�o��@>A���ٿ���o���@	*�4�3@SxUu�!?�K7�o��@��'s�ٿm��A���@���4@֣Q�Q�!?X�_ӏ�@��X9�ٿaNs.z,�@�Fg���3@w��a`�!?�'but�@v�U���ٿ�8�Mp�@�1I�3@��r�S�!?��S\Ϊ�@v�U���ٿ�8�Mp�@�1I�3@��r�S�!?��S\Ϊ�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Zb>��ٿ�Q�=���@�����3@Mnk��!?z�A"�@Y��w�ٿ��\�@4�5���3@T���A�!?�A�8�L�@Y��w�ٿ��\�@4�5���3@T���A�!?�A�8�L�@�xvjM�ٿ�2vò��@m�.��4@�K�3�!?�����@�xvjM�ٿ�2vò��@m�.��4@�K�3�!?�����@�xvjM�ٿ�2vò��@m�.��4@�K�3�!?�����@�xvjM�ٿ�2vò��@m�.��4@�K�3�!?�����@�xvjM�ٿ�2vò��@m�.��4@�K�3�!?�����@��-͓ٿ��]����@����04@?8O�j�!?��B��@��-͓ٿ��]����@����04@?8O�j�!?��B��@��-͓ٿ��]����@����04@?8O�j�!?��B��@�r�  �ٿ3� <��@����3@����0�!?�{Kݣ�@�r�  �ٿ3� <��@����3@����0�!?�{Kݣ�@�r�  �ٿ3� <��@����3@����0�!?�{Kݣ�@�r�  �ٿ3� <��@����3@����0�!?�{Kݣ�@�r�  �ٿ3� <��@����3@����0�!?�{Kݣ�@4�SYɚٿ��&<|�@��*I?�3@�`X:�!?��z'q��@4�SYɚٿ��&<|�@��*I?�3@�`X:�!?��z'q��@4�SYɚٿ��&<|�@��*I?�3@�`X:�!?��z'q��@4�SYɚٿ��&<|�@��*I?�3@�`X:�!?��z'q��@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@���
�ٿ>*Y�}�@�����3@���Sc�!?7c;M寴@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@nH�0��ٿ���J�@p*c��3@؅��P�!?bA�~ٴ@�4⊸�ٿ@+B�.��@�)c��4@v^}m>�!?@4v�P�@�4⊸�ٿ@+B�.��@�)c��4@v^}m>�!?@4v�P�@�4⊸�ٿ@+B�.��@�)c��4@v^}m>�!?@4v�P�@�N8z�ٿtr�(���@iC�C�3@���ȏ!?����6�@�N8z�ٿtr�(���@iC�C�3@���ȏ!?����6�@�N8z�ٿtr�(���@iC�C�3@���ȏ!?����6�@�N8z�ٿtr�(���@iC�C�3@���ȏ!?����6�@YA�$�ٿ�7�����@!C�O�3@ܖ�@�!?��3F��@YA�$�ٿ�7�����@!C�O�3@ܖ�@�!?��3F��@YA�$�ٿ�7�����@!C�O�3@ܖ�@�!?��3F��@���̔ٿ�ifċ�@ml�ټ�3@�G����!?)�?a�p�@���̔ٿ�ifċ�@ml�ټ�3@�G����!?)�?a�p�@���̔ٿ�ifċ�@ml�ټ�3@�G����!?)�?a�p�@���̔ٿ�ifċ�@ml�ټ�3@�G����!?)�?a�p�@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@=t����ٿ�N6o�G�@�<�Q��3@4S5V�!?8�a�ߴ@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@�;�ےٿN7���@Ά&۱�3@(d�W�!?f <�V״@6b,�ٿ�������@ƨ��F�3@���7�!?��ϴ挴@6b,�ٿ�������@ƨ��F�3@���7�!?��ϴ挴@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@䢎�J�ٿ�[9�@�h����3@�
 s�!?Q�*�@x�tN��ٿHϱO�@U����3@��Q�!?�L��@x�tN��ٿHϱO�@U����3@��Q�!?�L��@.��3c�ٿd�뫈�@X���3@�����!?�\����@.��3c�ٿd�뫈�@X���3@�����!?�\����@.��3c�ٿd�뫈�@X���3@�����!?�\����@.��3c�ٿd�뫈�@X���3@�����!?�\����@.��3c�ٿd�뫈�@X���3@�����!?�\����@.��3c�ٿd�뫈�@X���3@�����!?�\����@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@�`T���ٿ���:�2�@�!$�c�3@w�]�!?�)�w�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@q֪kD�ٿ�f��xM�@��8�3@�֚zv�!?�j�D~M�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@7C5?�ٿ}��Z^��@�FD�3@=�E�!?:��E)�@CUk��ٿG�?���@�m����3@� �E5�!?���Nkڴ@CUk��ٿG�?���@�m����3@� �E5�!?���Nkڴ@CUk��ٿG�?���@�m����3@� �E5�!?���Nkڴ@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@��ԅ��ٿ�5/�f��@�\?��3@w�P�!?�4*��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@8��Չ�ٿ+lN���@2��M��3@��=vW�!?�?�7��@~� ��ٿ,���s�@��YM�4@K��$n�!?O�9�k�@�\���ٿ��,+��@qU6��4@C�롔�!?��y޺��@��^��ٿ�n*��@�}.��4@n�͐!?�p|�Ҵ@��^��ٿ�n*��@�}.��4@n�͐!?�p|�Ҵ@��^��ٿ�n*��@�}.��4@n�͐!?�p|�Ҵ@��^��ٿ�n*��@�}.��4@n�͐!?�p|�Ҵ@��^��ٿ�n*��@�}.��4@n�͐!?�p|�Ҵ@D�+�ٿ�&T�\�@���X�3@��(���!?G�uEŴ@�3�0�ٿ5�-{3�@aÇt��3@`'�l�!?���|�@�3�0�ٿ5�-{3�@aÇt��3@`'�l�!?���|�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@^ 9�R�ٿ�6?����@C�Ȭ��3@��},�!?�}��8�@;.��p�ٿÁz퍔�@Ll�O�3@Ŕ��4�!? ��sڴ@;.��p�ٿÁz퍔�@Ll�O�3@Ŕ��4�!? ��sڴ@;.��p�ٿÁz퍔�@Ll�O�3@Ŕ��4�!? ��sڴ@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@LYc��ٿ� �䫽�@<���3@0
tPY�!?��Dɉx�@A#-I�ٿ�:����@.A:��3@n��*�!?�z���۴@e�x�^�ٿ��n鏍�@�o�44@@��&�!?�Ŵ��˴@e�x�^�ٿ��n鏍�@�o�44@@��&�!?�Ŵ��˴@e�x�^�ٿ��n鏍�@�o�44@@��&�!?�Ŵ��˴@��"�4�ٿ*���]�@�d;��3@Rb't7�!?�č����@��"�4�ٿ*���]�@�d;��3@Rb't7�!?�č����@��"�4�ٿ*���]�@�d;��3@Rb't7�!?�č����@W���ߖٿ0��D�@ê�1�3@�����!?'�=��Y�@W���ߖٿ0��D�@ê�1�3@�����!?'�=��Y�@W���ߖٿ0��D�@ê�1�3@�����!?'�=��Y�@W���ߖٿ0��D�@ê�1�3@�����!?'�=��Y�@W���ߖٿ0��D�@ê�1�3@�����!?'�=��Y�@<�X2��ٿp˶:��@u9>_��3@�����!?�;q�@<�X2��ٿp˶:��@u9>_��3@�����!?�;q�@�c�ٿ��?m�N�@���m��3@g�9d�!?r��y=*�@�c�ٿ��?m�N�@���m��3@g�9d�!?r��y=*�@�c�ٿ��?m�N�@���m��3@g�9d�!?r��y=*�@�v��^�ٿ�����'�@�����3@��iV�!?�a`.��@�v��^�ٿ�����'�@�����3@��iV�!?�a`.��@�v��^�ٿ�����'�@�����3@��iV�!?�a`.��@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@<XȀ�ٿ0�P���@|����3@j�@���!?x���ش@{�w}�ٿkRR�B�@5јy��3@+E~�u�!?��?�7ȴ@{�w}�ٿkRR�B�@5јy��3@+E~�u�!?��?�7ȴ@{�w}�ٿkRR�B�@5јy��3@+E~�u�!?��?�7ȴ@{�w}�ٿkRR�B�@5јy��3@+E~�u�!?��?�7ȴ@����ٿ��ٳcӿ@r��d�3@��1ڄ�!?���M�@����ٿ��ٳcӿ@r��d�3@��1ڄ�!?���M�@��\0��ٿ�V0�믿@�m%��3@�&#�!?^{�&��@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@c+VD�ٿ�^h/�4�@����3@B��sD�!?�-N~/~�@���
�ٿ�����~�@����3@�l�L�!? $�*ա�@P�c �ٿ�gr\�\�@���M��3@�RRp�!?�wP�V��@P�c �ٿ�gr\�\�@���M��3@�RRp�!?�wP�V��@P�c �ٿ�gr\�\�@���M��3@�RRp�!?�wP�V��@P�c �ٿ�gr\�\�@���M��3@�RRp�!?�wP�V��@�x����ٿ�E�5�@�w>��3@��rRL�!?1�DI��@r9/�ٿV�zU�@�z.F�3@���o��!?!��*Gϴ@r9/�ٿV�zU�@�z.F�3@���o��!?!��*Gϴ@r9/�ٿV�zU�@�z.F�3@���o��!?!��*Gϴ@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@�P��ٿ~)ڳ��@���?�3@s���a�!?���Ȝ��@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@wX~Õٿ�s�'A��@/�Bb�3@�*Gr��!?��d����@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@ygg�ٿ�^�(���@};���3@n �qD�!?�H�r#�@���pZ�ٿ�d�3^�@_uͼ�3@M�g�!?��׫�@���pZ�ٿ�d�3^�@_uͼ�3@M�g�!?��׫�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@��e���ٿ �0��@�>((��3@�6WQ��!?k���l}�@������ٿ���@@��.��3@2�K�!?l%�_�:�@������ٿ���@@��.��3@2�K�!?l%�_�:�@������ٿ���@@��.��3@2�K�!?l%�_�:�@���GB�ٿ��_�4��@�ڂU!�3@�w�Rs�!?���o8��@���GB�ٿ��_�4��@�ڂU!�3@�w�Rs�!?���o8��@���GB�ٿ��_�4��@�ڂU!�3@�w�Rs�!?���o8��@n�k��ٿ�ڌ6���@�!���3@�.̹�!?�m�8\.�@n�k��ٿ�ڌ6���@�!���3@�.̹�!?�m�8\.�@n�k��ٿ�ڌ6���@�!���3@�.̹�!?�m�8\.�@n�k��ٿ�ڌ6���@�!���3@�.̹�!?�m�8\.�@n�k��ٿ�ڌ6���@�!���3@�.̹�!?�m�8\.�@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@h!=�<�ٿ��WAG�@9t��l�3@�8�|��!?d�@#��@�8��Ƙٿ��|�tj�@�.8��3@�Y�5t�!?ƃ���@�����ٿ�V���@�Ыˆ�3@�)R���!?�]ދ}��@_�d܍ٿ	���S�@����3@���Sk�!?6}pI^�@(��xW�ٿ�|'�$�@1�����3@v���F�!?�ϟ�*n�@(��xW�ٿ�|'�$�@1�����3@v���F�!?�ϟ�*n�@(��xW�ٿ�|'�$�@1�����3@v���F�!?�ϟ�*n�@(��xW�ٿ�|'�$�@1�����3@v���F�!?�ϟ�*n�@?F���ٿ�xt�C�@�VuX��3@?ӭ$��!?)��N���@?F���ٿ�xt�C�@�VuX��3@?ӭ$��!?)��N���@6�+���ٿskf�Mo�@G:c��3@YNTd�!?�'�Apе@*h�Ӳ�ٿ��q���@"!�%�3@$��o�!?p	/�4��@*h�Ӳ�ٿ��q���@"!�%�3@$��o�!?p	/�4��@*h�Ӳ�ٿ��q���@"!�%�3@$��o�!?p	/�4��@*h�Ӳ�ٿ��q���@"!�%�3@$��o�!?p	/�4��@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@���\��ٿbŮ�f��@x�x��3@h>�K�!?	���dC�@�����ٿ��~��@�d9�3@�d��E�!?����Z�@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@n�vk�ٿ��S��]�@y�<C�3@L��I�!?Tz ���@�� ΒٿU�w��M�@�MA��3@p�YL��!?�O�&��@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@Ζ�W�ٿ�9�4M��@-Ԥ��3@���gl�!?N�����@�o���ٿ0C��,i�@�f����3@O7�ɛ�!?v&n��@�o���ٿ0C��,i�@�f����3@O7�ɛ�!?v&n��@��O��ٿ�D7�\�@MF#��3@�y�b{�!?Wc��^c�@��O��ٿ�D7�\�@MF#��3@�y�b{�!?Wc��^c�@;Dm�M�ٿ`) @�g�@�+6 4@>�
A0�!?��X��8�@���y�ٿX5�0w�@6��A�3@�+�N*�!?���1[�@���y�ٿX5�0w�@6��A�3@�+�N*�!?���1[�@���y�ٿX5�0w�@6��A�3@�+�N*�!?���1[�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@�p�ٿ��/���@�tZ4�3@���qG�!?�Ԑ_L�@ۄ��ڒٿ9��+qf�@��B�o�3@HmNP<�!?7�'Q�@ۄ��ڒٿ9��+qf�@��B�o�3@HmNP<�!?7�'Q�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@��R�ٿ������@�۩Z�3@I�䦎�!?�A�'0�@!:�ʿ�ٿ�ʯn�@�_��p�3@��HIK�!?��a@�@!:�ʿ�ٿ�ʯn�@�_��p�3@��HIK�!?��a@�@!:�ʿ�ٿ�ʯn�@�_��p�3@��HIK�!?��a@�@�>��V�ٿ�b1����@��֌�3@q�8�M�!?�����i�@R��m6�ٿ�~����@Á���3@ �_=�!?O����#�@#�}E��ٿ���'"Z�@\��?�3@O��"�!?r�n�Z��@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@V�+�~�ٿ����&��@�]��P�3@�����!?�312Z�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@��ϜٿR̘<4�@_I���3@�:Ӊ;�!?����+�@n�� T�ٿ|=78�@Dr�ݑ�3@~�n�1�!?�� l�@��X�Ėٿ&�4�L
�@X���3@�R���!?���h�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@J�/k�ٿX�:��@b:-7(�3@b_1+�!?�a�EG�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@o�J�d�ٿPei�^�@ǩ��B�3@����!?���ԙ�@[���d�ٿ�A�L�@e-;�#�3@�����!?��{�@<�@[���d�ٿ�A�L�@e-;�#�3@�����!?��{�@<�@L����ٿ~*��>��@�� ���3@�W#&�!?��m���@L����ٿ~*��>��@�� ���3@�W#&�!?��m���@L����ٿ~*��>��@�� ���3@�W#&�!?��m���@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@|�@�ٿ?Wx8�@�TR�3@���:I�!?� �O��@�3KyT�ٿ0��l�P�@�h	}�3@@%t>�!?	n���@��H��ٿ�	��@/�'���3@�y���!?���3Դ@��H��ٿ�	��@/�'���3@�y���!?���3Դ@9�$�=�ٿ4���`��@EyƯ�3@�$8t,�!?t`/l"
�@9�$�=�ٿ4���`��@EyƯ�3@�$8t,�!?t`/l"
�@9�$�=�ٿ4���`��@EyƯ�3@�$8t,�!?t`/l"
�@��+Ęٿ���I�@aE�<��3@��YV�!?]vS�´@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@
&���ٿ-ǯ���@���3@�޿&F�!?�_edش@@�YH�ٿ��i�@N��Ǻ�3@����!?�3W���@)TȀ	�ٿ��$pe��@�	�?�3@�؞Ϗ!?��cb��@莖��ٿ�)���~�@�����3@��U�!?�O�?T�@�Yd�ٿG���V��@�ԟq��3@��W�!?u/��C�@�Yd�ٿG���V��@�ԟq��3@��W�!?u/��C�@���iI�ٿ�֝e��@�$��3@�QX��!?sw�۴��@��+U�ٿ�#ټ��@e�o��3@���9�!?���Q��@�D5~�ٿ�	ߧ}\�@�2��3@����E�!?���%���@5���A�ٿ�0����@��N�4@�^Agz�!?4��p+��@5���A�ٿ�0����@��N�4@�^Agz�!?4��p+��@5���A�ٿ�0����@��N�4@�^Agz�!?4��p+��@5���A�ٿ�0����@��N�4@�^Agz�!?4��p+��@z6�ڙٿ�� �?&�@�a~$�4@�����!?7uu�aD�@z6�ڙٿ�� �?&�@�a~$�4@�����!?7uu�aD�@U7�ȕٿ:՟�S)�@��W�3@���͏!?%��L-+�@&�@�ٿ�_n�.�@�;���3@��/3�!?��f$&8�@&�@�ٿ�_n�.�@�;���3@��/3�!?��f$&8�@&�@�ٿ�_n�.�@�;���3@��/3�!?��f$&8�@&�@�ٿ�_n�.�@�;���3@��/3�!?��f$&8�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=�Ӷ3�ٿ�+y���@��}�L4@����k�!?Jnu+B�@=���u�ٿ�sz����@�nʚ�4@�	/M��!?��118۴@=���u�ٿ�sz����@�nʚ�4@�	/M��!?��118۴@�w�wQ�ٿ��*���@��z�T�3@���!?N,��_5�@�w�wQ�ٿ��*���@��z�T�3@���!?N,��_5�@�w�wQ�ٿ��*���@��z�T�3@���!?N,��_5�@ AX�:�ٿ����I�@#�ܣT�3@����Ð!?'u�~ɴ@w�B�ٿ�zU(��@C�UAE�3@͕Y��!? �]Mq1�@w�B�ٿ�zU(��@C�UAE�3@͕Y��!? �]Mq1�@w�B�ٿ�zU(��@C�UAE�3@͕Y��!? �]Mq1�@M=�s �ٿs�uW���@���L�3@��򆼐!?�_�d��@M=�s �ٿs�uW���@���L�3@��򆼐!?�_�d��@M=�s �ٿs�uW���@���L�3@��򆼐!?�_�d��@M=�s �ٿs�uW���@���L�3@��򆼐!?�_�d��@;ўx`�ٿ�n��1�@4�0�3@�k�l�!?��n�Y`�@����ݗٿ���[�@�e�@��3@����!?'������@����ݗٿ���[�@�e�@��3@����!?'������@����ݗٿ���[�@�e�@��3@����!?'������@����ݗٿ���[�@�e�@��3@����!?'������@����ݗٿ���[�@�e�@��3@����!?'������@����ݗٿ���[�@�e�@��3@����!?'������@@3$�F�ٿ���0�@�煮�3@�L(��!?D��␵@�ih�ٿ-r���X�@x���4@d]Ou�!?�����'�@�ې|7�ٿ�@���@� 3I��3@	�h�!?zʜ�´@�ې|7�ٿ�@���@� 3I��3@	�h�!?zʜ�´@�ې|7�ٿ�@���@� 3I��3@	�h�!?zʜ�´@�ې|7�ٿ�@���@� 3I��3@	�h�!?zʜ�´@�ې|7�ٿ�@���@� 3I��3@	�h�!?zʜ�´@u��z��ٿ/u�K�@���/4@Ǉ �!?Q��8��@бi���ٿ���%�n�@e�tQ��3@8|!�܏!?����ݴ@	̖��ٿ�ֿ��{�@`�4@&�!?E����@�����ٿ�ju, ��@�	��i�3@�隦��!?���<Hx�@�����ٿ�ju, ��@�	��i�3@�隦��!?���<Hx�@�����ٿ�ju, ��@�	��i�3@�隦��!?���<Hx�@�f�k�ٿ;�КY�@�.��>�3@�f�Q��!?��m-Ma�@�f�k�ٿ;�КY�@�.��>�3@�f�Q��!?��m-Ma�@�f�k�ٿ;�КY�@�.��>�3@�f�Q��!?��m-Ma�@�f�k�ٿ;�КY�@�.��>�3@�f�Q��!?��m-Ma�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@��B_�ٿ�_6�@�Ϙ�p�3@Tp�e�!?D�r��E�@!=�9�ٿs�a�,�@I�6��3@��?�!?��F+��@!=�9�ٿs�a�,�@I�6��3@��?�!?��F+��@!=�9�ٿs�a�,�@I�6��3@��?�!?��F+��@!=�9�ٿs�a�,�@I�6��3@��?�!?��F+��@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@����4�ٿ�4����@vt����3@w/W��!?Ս_!�T�@q@���ٿ�1� �@�<�6i�3@/��a�!?\*��x�@q@���ٿ�1� �@�<�6i�3@/��a�!?\*��x�@q@���ٿ�1� �@�<�6i�3@/��a�!?\*��x�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@7�V��ٿ$P4���@z��V-4@��gy��!?)f�Hd�@��3�ٿ11J�&�@#|�v4@m�U�t�!?�ֲ����@�N,�ٿp����@d
�ܯ�3@P�~���!?�&N�U�@�N,�ٿp����@d
�ܯ�3@P�~���!?�&N�U�@�N,�ٿp����@d
�ܯ�3@P�~���!?�&N�U�@�'�ٿo�����@����3�3@W ]b�!?�M0Հ�@�'�ٿo�����@����3�3@W ]b�!?�M0Հ�@t�9�ٿF.`���@X�����3@����!?o��z��@�2�EG�ٿj��6k�@^�x��3@E���V�!?4�Rٳ�@{\sR�ٿO�zR��@-��z�3@Q8��!?�l˒U�@{\sR�ٿO�zR��@-��z�3@Q8��!?�l˒U�@{\sR�ٿO�zR��@-��z�3@Q8��!?�l˒U�@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@��}f�ٿ+�R�H�@��lL�3@yZw�!?�q�x��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@!3}��ٿp8~���@2)�?��3@�b�b�!?⤒'��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@P�KD�ٿ�
��I��@R:�ӎ�3@7��D{�!?�:}7��@^)��"�ٿ�lI����@��{4Z�3@{�W���!?�5���@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@����ٿ�V�t~�@�R�
�3@��ᑐ!?�R�^u�@�|�?�ٿ�V��@��ۜ�3@�Lo�i�!?H�qɏK�@�|�?�ٿ�V��@��ۜ�3@�Lo�i�!?H�qɏK�@�|�?�ٿ�V��@��ۜ�3@�Lo�i�!?H�qɏK�@U����ٿ��Q��?�@����3@��T�,�!?ևh[��@U����ٿ��Q��?�@����3@��T�,�!?ևh[��@d
�h��ٿ��	Ei�@����S�3@P�����!?�q� ��@d
�h��ٿ��	Ei�@����S�3@P�����!?�q� ��@�;�g��ٿ/i��s�@�G6S��3@��y#G�!?�u�K��@Ѭ��~�ٿ�G�FY�@�����3@�c���!?jU-mZ�@Ѭ��~�ٿ�G�FY�@�����3@�c���!?jU-mZ�@Ѭ��~�ٿ�G�FY�@�����3@�c���!?jU-mZ�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@SK�L��ٿ�*��c�@H͚���3@)UրM�!?Jp⺱�@ݍ�K�ٿ<\'���@S��\��3@���z�!?E5��@ݍ�K�ٿ<\'���@S��\��3@���z�!?E5��@ݍ�K�ٿ<\'���@S��\��3@���z�!?E5��@ݍ�K�ٿ<\'���@S��\��3@���z�!?E5��@ݍ�K�ٿ<\'���@S��\��3@���z�!?E5��@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@���J�ٿ��4���@ �����3@w�_�!?��o���@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@l��o@�ٿ��T}���@�Djr�3@�9���!?�&�`'�@���sϗٿ.�\�\�@�&j#��3@��M�,�!?�`�@���sϗٿ.�\�\�@�&j#��3@��M�,�!?�`�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@X��%ݔٿ)�Mp]��@������3@���T�!?K�bN�@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@`G����ٿ�xr�^�@9z��4@�%� W�!?s�2Q��@�R���ٿ���ꋖ�@����3@�g�P�!?�50��@�R���ٿ���ꋖ�@����3@�g�P�!?�50��@Ȝ�%�ٿ�{�E`�@�3u��3@=��[U�!?H�!��A�@Ȝ�%�ٿ�{�E`�@�3u��3@=��[U�!?H�!��A�@Ȝ�%�ٿ�{�E`�@�3u��3@=��[U�!?H�!��A�@Ȝ�%�ٿ�{�E`�@�3u��3@=��[U�!?H�!��A�@�����ٿ5ͳn���@r�Ek_�3@zCkD�!?����@i��E�ٿ`���x�@�O�x�3@�-M�s�!?Na�%�Ĵ@j�'��ٿ��}��@]>��4@��(��!?����x�@j�'��ٿ��}��@]>��4@��(��!?����x�@j�'��ٿ��}��@]>��4@��(��!?����x�@j�'��ٿ��}��@]>��4@��(��!?����x�@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@T�p�N�ٿAФP%d�@���B�3@L|?�x�!?lJ�o��@А��ٿ���h�
�@1��3@�X
�"�!?=�s�i��@А��ٿ���h�
�@1��3@�X
�"�!?=�s�i��@А��ٿ���h�
�@1��3@�X
�"�!?=�s�i��@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@5a� �ٿ�3�.���@�����3@;Xd�Q�!?,��ȴ@��HV�ٿ�A]B��@�����3@c_��!?�쒤�@��HV�ٿ�A]B��@�����3@c_��!?�쒤�@��HV�ٿ�A]B��@�����3@c_��!?�쒤�@��HV�ٿ�A]B��@�����3@c_��!?�쒤�@��HV�ٿ�A]B��@�����3@c_��!?�쒤�@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@���țٿy��(x�@�VG ��3@�ء���!?-�����@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@��t\*�ٿYp�]��@�H��/�3@����S�!?�������@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���!�ٿ�e��Q�@AU��r�3@R_��;�!?
�V_}K�@���m#�ٿ\��d,#�@AW���3@h�N��!?A�w=�*�@1&)g�ٿ���b1��@E�. 4@-��!?�i&Z��@�I�l8�ٿ���?b�@�9���3@��lf�!?�C�*�3�@�I�l8�ٿ���?b�@�9���3@��lf�!?�C�*�3�@�I�l8�ٿ���?b�@�9���3@��lf�!?�C�*�3�@��ڗٿ���T�@�W�?�3@���m�!?	�8�a�@��ڗٿ���T�@�W�?�3@���m�!?	�8�a�@��ڗٿ���T�@�W�?�3@���m�!?	�8�a�@��ڗٿ���T�@�W�?�3@���m�!?	�8�a�@�1|��ٿr��ƙ�@��N��4@;Q r�!?c9M2��@�1|��ٿr��ƙ�@��N��4@;Q r�!?c9M2��@��Z�ٿ�5&T���@E4��4@2��h�!?o��8�ŵ@�B�G��ٿ�Rq��@o�Ǯ!4@�9ZUz�!?���8x�@�B�G��ٿ�Rq��@o�Ǯ!4@�9ZUz�!?���8x�@�B�G��ٿ�Rq��@o�Ǯ!4@�9ZUz�!?���8x�@�B�G��ٿ�Rq��@o�Ǯ!4@�9ZUz�!?���8x�@S[�+�ٿ�(���@lc���4@�hM��!?cbd#��@<� 1��ٿ��b=�@���c�4@�;;���!?+�_�3�@<� 1��ٿ��b=�@���c�4@�;;���!?+�_�3�@<� 1��ٿ��b=�@���c�4@�;;���!?+�_�3�@<� 1��ٿ��b=�@���c�4@�;;���!?+�_�3�@K�Z��ٿ��a,���@.�K~4@�
֐!?4�۴@p�F�u�ٿb
5:h��@2���� 4@b�ߠ��!?,�|���@p�F�u�ٿb
5:h��@2���� 4@b�ߠ��!?,�|���@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@Sw��r�ٿX ,� �@"�(>4@�&朐!?�l�5Ѵ@H����ٿ�Ǳ����@�����3@/��ɖ�!?`4��u�@H����ٿ�Ǳ����@�����3@/��ɖ�!?`4��u�@H����ٿ�Ǳ����@�����3@/��ɖ�!?`4��u�@H����ٿ�Ǳ����@�����3@/��ɖ�!?`4��u�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@g��\�ٿI�s�V��@�(Y��3@�q��7�!?W3���f�@�N �8�ٿ�%]E�G�@_<�~�3@"��#�!?���
z��@�N �8�ٿ�%]E�G�@_<�~�3@"��#�!?���
z��@�N �8�ٿ�%]E�G�@_<�~�3@"��#�!?���
z��@�N �8�ٿ�%]E�G�@_<�~�3@"��#�!?���
z��@�N �8�ٿ�%]E�G�@_<�~�3@"��#�!?���
z��@XϢi��ٿ�����@16����3@��E�!?���,j�@R>���ٿ�|�_�n�@4�?J��3@m�k�L�!?KkN��9�@�
1��ٿ�����@زO���3@� A	�!?~��a�ε@�
1��ٿ�����@زO���3@� A	�!?~��a�ε@�
1��ٿ�����@زO���3@� A	�!?~��a�ε@ٔG� �ٿE��n��@�Kx�N�3@l��a&�!?d
�]�@ٔG� �ٿE��n��@�Kx�N�3@l��a&�!?d
�]�@X���ٿ�0�=�"�@l(R�3@:v���!?�M��,k�@X���ٿ�0�=�"�@l(R�3@:v���!?�M��,k�@X���ٿ�0�=�"�@l(R�3@:v���!?�M��,k�@hpmw��ٿ�M;5)�@���� 4@�I��!?R0rd;&�@hpmw��ٿ�M;5)�@���� 4@�I��!?R0rd;&�@�Qݔٿz4ױ�@Af��3@q!Pk8�!?j��X镵@M�\J�ٿ�xA{�!�@��ߦO 4@b��*�!?�����@M�\J�ٿ�xA{�!�@��ߦO 4@b��*�!?�����@X>e��ٿi���Yq�@#��؏�3@.����!?��wyg��@X>e��ٿi���Yq�@#��؏�3@.����!?��wyg��@X>e��ٿi���Yq�@#��؏�3@.����!?��wyg��@=����ٿ�f$9�P�@�A�[��3@��E#��!?-3Ӽ�g�@=����ٿ�f$9�P�@�A�[��3@��E#��!?-3Ӽ�g�@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@ ԫ/��ٿ��e�@��2���3@8�H�}�!?tq[��@Rg���ٿ�px��P�@���a��3@bJ�l|�!?����@�R
��ٿ�\1��@�f4���3@��Nq�!?���`ʺ�@���a��ٿ�&H(z=�@Ġ���3@ġ_n�!?�FhgА�@���a��ٿ�&H(z=�@Ġ���3@ġ_n�!?�FhgА�@�*�R�ٿl�����@Q���3@Q[�k�!?�dh�z�@�*�R�ٿl�����@Q���3@Q[�k�!?�dh�z�@�*�R�ٿl�����@Q���3@Q[�k�!?�dh�z�@�����ٿA�h���@ú��6�3@�Y71�!?��.xƒ�@�&3�N�ٿ�'J�,�@���X��3@�QxL�!?�T�Y�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�h��ٿ�qΗ~J�@�P��4@��"�!?�o�ݾ�@�B����ٿ�mKk��@|!��4@��C �!?���t�7�@�B����ٿ�mKk��@|!��4@��C �!?���t�7�@�B����ٿ�mKk��@|!��4@��C �!?���t�7�@�B����ٿ�mKk��@|!��4@��C �!?���t�7�@�B����ٿ�mKk��@|!��4@��C �!?���t�7�@;F���ٿ�ӅR�$�@C�V��	4@�� �!?M)r푴@}��m�ٿ�K�Y���@�LB�3@V4ZO�!?��ĸ�@}��m�ٿ�K�Y���@�LB�3@V4ZO�!?��ĸ�@}��m�ٿ�K�Y���@�LB�3@V4ZO�!?��ĸ�@}��m�ٿ�K�Y���@�LB�3@V4ZO�!?��ĸ�@}��m�ٿ�K�Y���@�LB�3@V4ZO�!?��ĸ�@deV�x�ٿ�fѸ�@}��p�3@��4�!?�4����@deV�x�ٿ�fѸ�@}��p�3@��4�!?�4����@deV�x�ٿ�fѸ�@}��p�3@��4�!?�4����@deV�x�ٿ�fѸ�@}��p�3@��4�!?�4����@�6�h��ٿ�[x#�B�@��SZ��3@J���&�!?"[]��@�6�h��ٿ�[x#�B�@��SZ��3@J���&�!?"[]��@e��j��ٿf��w��@������3@���:�!?C}X%�@e��j��ٿf��w��@������3@���:�!?C}X%�@e��j��ٿf��w��@������3@���:�!?C}X%�@e��j��ٿf��w��@������3@���:�!?C}X%�@���ȖٿN�iW��@oۉ��3@6����!?�b��C�@���ȖٿN�iW��@oۉ��3@6����!?�b��C�@��vV�ٿ,��ef�@�h�MB�3@#����!?x�R�z�@��vV�ٿ,��ef�@�h�MB�3@#����!?x�R�z�@��vV�ٿ,��ef�@�h�MB�3@#����!?x�R�z�@�F����ٿЄ���S�@��.c��3@c��jW�!?��6�JL�@�F����ٿЄ���S�@��.c��3@c��jW�!?��6�JL�@�F����ٿЄ���S�@��.c��3@c��jW�!?��6�JL�@�$�lf�ٿ�?[�m��@G��=��3@,Q�+�!?��ц��@J�E0��ٿ���(���@�o��v�3@thD��!?z�(��@J�E0��ٿ���(���@�o��v�3@thD��!?z�(��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@�bKq�ٿ�4GN��@�u
z�3@��4�!?�F3*>��@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��I}�ٿ�]�����@��ɄH�3@�&V�s�!?ɛo�R�@��n�ٿ��f ��@#+��3@��ƉY�!?��h�+{�@��n�ٿ��f ��@#+��3@��ƉY�!?��h�+{�@��n�ٿ��f ��@#+��3@��ƉY�!?��h�+{�@��n�ٿ��f ��@#+��3@��ƉY�!?��h�+{�@�F�S��ٿ.W��:p�@]{7��3@.��G��!?w�s	�y�@�F�S��ٿ.W��:p�@]{7��3@.��G��!?w�s	�y�@�F�S��ٿ.W��:p�@]{7��3@.��G��!?w�s	�y�@�����ٿ�n�?q/�@�S'�3@a�1j�!?drW�K��@��Ġ�ٿ��yJ�Y�@��k��3@�F���!?-����d�@��Ġ�ٿ��yJ�Y�@��k��3@�F���!?-����d�@��Ġ�ٿ��yJ�Y�@��k��3@�F���!?-����d�@��Ġ�ٿ��yJ�Y�@��k��3@�F���!?-����d�@��Ġ�ٿ��yJ�Y�@��k��3@�F���!?-����d�@���ٿ�9����@¹�h�3@8#�4�!?+�b���@���ٿ�9����@¹�h�3@8#�4�!?+�b���@���ٿ�9����@¹�h�3@8#�4�!?+�b���@���ٿ�9����@¹�h�3@8#�4�!?+�b���@���ٿ�9����@¹�h�3@8#�4�!?+�b���@|�T6&�ٿMh)�.��@�R<4�3@6���/�!?m�>�@|�T6&�ٿMh)�.��@�R<4�3@6���/�!?m�>�@|�T6&�ٿMh)�.��@�R<4�3@6���/�!?m�>�@|�T6&�ٿMh)�.��@�R<4�3@6���/�!?m�>�@|�T6&�ٿMh)�.��@�R<4�3@6���/�!?m�>�@�l���ٿ������@�8����3@��	k�!?%�V��@�/��3�ٿ1˖��0�@Eɿ��3@i���!?� �ŵ@�/��3�ٿ1˖��0�@Eɿ��3@i���!?� �ŵ@�/��3�ٿ1˖��0�@Eɿ��3@i���!?� �ŵ@7� [��ٿ�����)�@ηC��3@\GY �!?-cƣ��@7� [��ٿ�����)�@ηC��3@\GY �!?-cƣ��@7� [��ٿ�����)�@ηC��3@\GY �!?-cƣ��@7� [��ٿ�����)�@ηC��3@\GY �!?-cƣ��@:���H�ٿ�{���@L�vXt�3@z�dS.�!?���Q�@:���H�ٿ�{���@L�vXt�3@z�dS.�!?���Q�@:���H�ٿ�{���@L�vXt�3@z�dS.�!?���Q�@:���H�ٿ�{���@L�vXt�3@z�dS.�!?���Q�@:���H�ٿ�{���@L�vXt�3@z�dS.�!?���Q�@���ٿCK�b���@��z�*�3@<KD�V�!?�l�y�@d]-�8�ٿѹs�=�@Će5�3@�B;	�!?��|�W�@d]-�8�ٿѹs�=�@Će5�3@�B;	�!?��|�W�@d]-�8�ٿѹs�=�@Će5�3@�B;	�!?��|�W�@d]-�8�ٿѹs�=�@Će5�3@�B;	�!?��|�W�@���g�ٿ�ե���@W�'��3@��:�!?� �@���g�ٿ�ե���@W�'��3@��:�!?� �@���g�ٿ�ե���@W�'��3@��:�!?� �@���g�ٿ�ե���@W�'��3@��:�!?� �@��B(��ٿ���,��@ɘ�@@�3@~{�<�!?o+=��ϴ@"(�ߚ�ٿ ���a�@PK����3@.�Ш1�!?��pH��@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@���K՛ٿ@:�zҟ�@�5��E�3@�C}o�!?ͳ°�n�@4J2l�ٿ˨ά��@�����4@-�%m�!?ʐѭ��@4J2l�ٿ˨ά��@�����4@-�%m�!?ʐѭ��@��2\�ٿ�3Q�Jy�@�^*��3@�Oи��!?2�#�@��2\�ٿ�3Q�Jy�@�^*��3@�Oи��!?2�#�@���Zk�ٿ4�n����@��L���3@/��x��!?{�����@���Zk�ٿ4�n����@��L���3@/��x��!?{�����@���Zk�ٿ4�n����@��L���3@/��x��!?{�����@?����ٿ���Gi�@���l�3@�q����!?�)�]���@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@��^`��ٿ��<���@i�(��3@�����!?�,�K,�@�9	��ٿfz��f�@�
k�s�3@�c���!?X����@�9	��ٿfz��f�@�
k�s�3@�c���!?X����@Ő0ä�ٿU���B��@S�>��3@ѻ�Ķ�!?�.�@Ő0ä�ٿU���B��@S�>��3@ѻ�Ķ�!?�.�@Ő0ä�ٿU���B��@S�>��3@ѻ�Ķ�!?�.�@Ő0ä�ٿU���B��@S�>��3@ѻ�Ķ�!?�.�@Ő0ä�ٿU���B��@S�>��3@ѻ�Ķ�!?�.�@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@(�֑B�ٿ�I-=A�@�,T�4@��y�!?�x�a���@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@/3!�.�ٿe4W`+�@{Es�^�3@�n�^Q�!?RT�eߴ@���p�ٿ"�Ԟ��@���J�3@�g#H�!??�|k1��@���p�ٿ"�Ԟ��@���J�3@�g#H�!??�|k1��@���p�ٿ"�Ԟ��@���J�3@�g#H�!??�|k1��@���p�ٿ"�Ԟ��@���J�3@�g#H�!??�|k1��@���p�ٿ"�Ԟ��@���J�3@�g#H�!??�|k1��@"Qwɘٿ���]���@��K���3@�-5�!?�]uf�@"Qwɘٿ���]���@��K���3@�-5�!?�]uf�@���S�ٿ�O�	�	�@��n��3@$+M�@�!?�3H k��@���S�ٿ�O�	�	�@��n��3@$+M�@�!?�3H k��@���S�ٿ�O�	�	�@��n��3@$+M�@�!?�3H k��@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@LT�n��ٿzFt���@fSr.d�3@���bi�!?�:���2�@��ZƑٿ����@�@��զ?�3@@#d�n�!?Trh=��@��ZƑٿ����@�@��զ?�3@@#d�n�!?Trh=��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@P��nזٿ�M)˒�@�Vt�4@�:骐�!?���.*��@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@):��~�ٿ�Ӧ�*�@�@#l�4@4�"�z�!?�����@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@���%�ٿJ��U,�@"tH�4@��
�1�!?��p���@�����ٿ�;�SMn�@4jB�M
4@:uF��!? �k����@���<��ٿR�����@�I���3@+�!f�!?4)�@P�@���<��ٿR�����@�I���3@+�!f�!?4)�@P�@��Ҿ��ٿ�/]5���@'�p�J�3@��S50�!?�w�E��@��Ҿ��ٿ�/]5���@'�p�J�3@��S50�!?�w�E��@F�ߊ��ٿ-W��d��@�#�E��3@��	c�!?���D��@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@cn�=t�ٿ�2�H�@���3@�ǧʃ�!?�E�>3�@^�lyגٿ` �k�@��#kZ�3@���Z�!?_�k�ĵ@^�lyגٿ` �k�@��#kZ�3@���Z�!?_�k�ĵ@��̐ٿw�V���@{���N 4@'��c�!?��{ �N�@��̐ٿw�V���@{���N 4@'��c�!?��{ �N�@�Aݴ#�ٿ�����@����3@W��J��!?1r��0�@�Aݴ#�ٿ�����@����3@W��J��!?1r��0�@�Aݴ#�ٿ�����@����3@W��J��!?1r��0�@���f�ٿ����+��@�$G�3@J�-�~�!?��6|�@���f�ٿ����+��@�$G�3@J�-�~�!?��6|�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@�M��ٿ�B6���@�����3@��f��!?p.'�&�@���3�ٿ������@�𢸔�3@�OeY�!?xS����@��ٿ�ޏ���@��u�N�3@I��\��!?�[_��C�@��ٿ�ޏ���@��u�N�3@I��\��!?�[_��C�@��ٿ�ޏ���@��u�N�3@I��\��!?�[_��C�@��ٿ�ޏ���@��u�N�3@I��\��!?�[_��C�@��ٿ�ޏ���@��u�N�3@I��\��!?�[_��C�@���ٿ��А�@�W��\�3@�A����!?��ܫ�@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�B����ٿ��k6|�@[�V��3@�Δʅ�!?�.˕o��@�o��ٿ���l���@�+r� 4@��`Z��!?Ģ۶��@�o��ٿ���l���@�+r� 4@��`Z��!?Ģ۶��@�o��ٿ���l���@�+r� 4@��`Z��!?Ģ۶��@�o��ٿ���l���@�+r� 4@��`Z��!?Ģ۶��@�o��ٿ���l���@�+r� 4@��`Z��!?Ģ۶��@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@�>g��ٿ�o�9�W�@����3@������!?E��$�@��C�ٿ��Y��@�����3@��yŬ�!?�٩MR�@h��w��ٿD�ݢvh�@(���|�3@�
;�ڐ!?f�J�(J�@h��w��ٿD�ݢvh�@(���|�3@�
;�ڐ!?f�J�(J�@c^7h�ٿ�F����@�s�y�3@KGVs��!?.%�o��@c^7h�ٿ�F����@�s�y�3@KGVs��!?.%�o��@c^7h�ٿ�F����@�s�y�3@KGVs��!?.%�o��@c^7h�ٿ�F����@�s�y�3@KGVs��!?.%�o��@c^7h�ٿ�F����@�s�y�3@KGVs��!?.%�o��@n`�G��ٿl�T�W]�@�|.z��3@A%��!?��E�=��@n`�G��ٿl�T�W]�@�|.z��3@A%��!?��E�=��@n`�G��ٿl�T�W]�@�|.z��3@A%��!?��E�=��@T/��K�ٿL8!��@��D<�3@���wڐ!?q����@T/��K�ٿL8!��@��D<�3@���wڐ!?q����@T/��K�ٿL8!��@��D<�3@���wڐ!?q����@T/��K�ٿL8!��@��D<�3@���wڐ!?q����@T/��K�ٿL8!��@��D<�3@���wڐ!?q����@����p�ٿ�yk���@$�t�V4@��n��!?T�AYٵ@����p�ٿ�yk���@$�t�V4@��n��!?T�AYٵ@����p�ٿ�yk���@$�t�V4@��n��!?T�AYٵ@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@4Ȓ2��ٿ�)��M�@C9�N�3@r�U���!?�#����@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�7��ٿ �y �@ �3���3@Ou3z�!?���Y�@�r���ٿ�[��L.�@�lxB^�3@+��9\�!??�ݧ�L�@�r���ٿ�[��L.�@�lxB^�3@+��9\�!??�ݧ�L�@�r���ٿ�[��L.�@�lxB^�3@+��9\�!??�ݧ�L�@I�Q��ٿ�!�{h��@�R��3@1�@�r�!?�`��@I�Q��ٿ�!�{h��@�R��3@1�@�r�!?�`��@I�Q��ٿ�!�{h��@�R��3@1�@�r�!?�`��@I�Q��ٿ�!�{h��@�R��3@1�@�r�!?�`��@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@R{���ٿH8�>��@S]S�3@j��6��!?�3�u�:�@��r��ٿn.�����@�]����3@h�c��!?w��Ե@�ÔR��ٿ@����@�U�#�3@�bs��!?*f��	�@�ÔR��ٿ@����@�U�#�3@�bs��!?*f��	�@�ÔR��ٿ@����@�U�#�3@�bs��!?*f��	�@~�Sf(�ٿ$*l@�i�@��m[�3@cN��U�!?W�*£�@~�Sf(�ٿ$*l@�i�@��m[�3@cN��U�!?W�*£�@~�Sf(�ٿ$*l@�i�@��m[�3@cN��U�!?W�*£�@�#GO�ٿD�g�#�@@4��=�3@�$04d�!?��4��M�@�#GO�ٿD�g�#�@@4��=�3@�$04d�!?��4��M�@�#GO�ٿD�g�#�@@4��=�3@�$04d�!?��4��M�@�#GO�ٿD�g�#�@@4��=�3@�$04d�!?��4��M�@�#GO�ٿD�g�#�@@4��=�3@�$04d�!?��4��M�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@��`�=�ٿ���t&�@�.#���3@*K��w�!?��c˄�@rЃ���ٿ�1�����@&��@��3@j��1�!?0�/ �@rЃ���ٿ�1�����@&��@��3@j��1�!?0�/ �@rЃ���ٿ�1�����@&��@��3@j��1�!?0�/ �@rЃ���ٿ�1�����@&��@��3@j��1�!?0�/ �@W�w�ٿ�["���@t98Q��3@v���֐!?�(-	l�@W�w�ٿ�["���@t98Q��3@v���֐!?�(-	l�@Ǟ�חٿ��C8�@:�h�N�3@��+�ѐ!?��u�P�@�/>("�ٿ8iK���@�e=S��3@k?ǐ!?<��,�@�/>("�ٿ8iK���@�e=S��3@k?ǐ!?<��,�@�/>("�ٿ8iK���@�e=S��3@k?ǐ!?<��,�@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@[{�㖖ٿ&�9�R��@��g��3@�6s�i�!?ñ�eܴ@�V�O�ٿ����@]��w�3@���E��!?u�M�H'�@�V�O�ٿ����@]��w�3@���E��!?u�M�H'�@�V�O�ٿ����@]��w�3@���E��!?u�M�H'�@�V�O�ٿ����@]��w�3@���E��!?u�M�H'�@�V�O�ٿ����@]��w�3@���E��!?u�M�H'�@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@�V�8Q�ٿ��^m'g�@x ��3@�r>��!?IY����@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@���ٿ@�z#��@6��+P�3@U�+|�!?���<�´@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@���2��ٿ��C ��@�O  4@�EP���!?��4A�@���2��ٿ��C ��@�O  4@�EP���!?��4A�@���2��ٿ��C ��@�O  4@�EP���!?��4A�@���2��ٿ��C ��@�O  4@�EP���!?��4A�@���2��ٿ��C ��@�O  4@�EP���!?��4A�@�����ٿU�����@I����3@��_�!?����4A�@�����ٿU�����@I����3@��_�!?����4A�@�����ٿU�����@I����3@��_�!?����4A�@�����ٿU�����@I����3@��_�!?����4A�@�����ٿU�����@I����3@��_�!?����4A�@��˖�ٿ�/�����@�o�1��3@$����!?�Nb�4A�@��˖�ٿ�/�����@�o�1��3@$����!?�Nb�4A�@�i�ߖ�ٿܕ|����@nVp���3@�c* �!?3�,�4A�@�i�ߖ�ٿܕ|����@nVp���3@�c* �!?3�,�4A�@�i�ߖ�ٿܕ|����@nVp���3@�c* �!?3�,�4A�@�i�ߖ�ٿܕ|����@nVp���3@�c* �!?3�,�4A�@���ܞ�ٿ��n����@`��G��3@��� �!?�r��4A�@L y���ٿ�������@�����3@�va|�!?Y��4A�@qeC㠙ٿ~�����@;�.L  4@ᆏ�q�!?2M��4A�@�+���ٿ-������@_�]��3@��^��!?$�|�4A�@��ǟ�ٿ�zH����@�J���3@��3祐!?L���4A�@��$���ٿ�h�����@L
{���3@�/
m��!?}5��4A�@��$���ٿ�h�����@L
{���3@�/
m��!?}5��4A�@��$���ٿ�h�����@L
{���3@�/
m��!?}5��4A�@.����ٿc������@��n  4@�����!?Nb��4A�@.����ٿc������@��n  4@�����!?Nb��4A�@3�	���ٿ�������@T�,  4@��[�Ð!?�0^�4A�@3�	���ٿ�������@T�,  4@��[�Ð!?�0^�4A�@��hq��ٿ4�j����@��ѐ 4@�)hT��!?k\�4A�@E�0��ٿR������@}�� 4@G�J���!?�޳�4A�@E�0��ٿR������@}�� 4@G�J���!?�޳�4A�@`����ٿh�n����@ܙ�w 4@����!?�̸4A�@`����ٿh�n����@ܙ�w 4@����!?�̸4A�@UU��ٿ�־����@Dc�� 4@���Yޏ!?A�Y�4A�@���f��ٿ�<{����@6!{  4@��I8��!?>%��4A�@���f��ٿ�<{����@6!{  4@��I8��!?>%��4A�@r�=��ٿ&����@�E�g  4@m_�I�!?�%�4A�@������ٿ������@ƥs*��3@1_H�!?=�}4A�@������ٿ������@ƥs*��3@1_H�!?=�}4A�@������ٿ������@ƥs*��3@1_H�!?=�}4A�@������ٿ������@ƥs*��3@1_H�!?=�}4A�@������ٿ������@ƥs*��3@1_H�!?=�}4A�@HII���ٿ�����@�����3@aނ�!?-W�4A�@HII���ٿ�����@�����3@aނ�!?-W�4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@.Ϣ�ٿ�:�����@dd�:��3@�-(���!?�B��4A�@�蘴��ٿN����@]�=���3@�B�!?�LC�4A�@�蘴��ٿN����@]�=���3@�B�!?�LC�4A�@�蘴��ٿN����@]�=���3@�B�!?�LC�4A�@X����ٿ��
����@�����3@����!?��
�4A�@X����ٿ��
����@�����3@����!?��
�4A�@X����ٿ��
����@�����3@����!?��
�4A�@X����ٿ��
����@�����3@����!?��
�4A�@l�^ѫ�ٿ<g����@ *���3@����'�!?��׸4A�@l�^ѫ�ٿ<g����@ *���3@����'�!?��׸4A�@�Y�q��ٿwv�����@��H��3@�:K�!?���4A�@0+򋣙ٿ������@����3@�Y	�$�!?(N�4A�@�B���ٿ}G����@|��"��3@ ��)�!?f��4A�@}�+���ٿKA�����@X-���3@�R(�!?��R�4A�@��yW��ٿ�0����@s?;���3@5Q���!?g<�4A�@��yW��ٿ�0����@s?;���3@5Q���!?g<�4A�@�)�;��ٿ�b ����@.����3@��N�!?��(�4A�@�)�;��ٿ�b ����@.����3@��N�!?��(�4A�@�)�;��ٿ�b ����@.����3@��N�!?��(�4A�@�)�;��ٿ�b ����@.����3@��N�!?��(�4A�@�M\��ٿ�������@�uW���3@̟"|��!?�bљ4A�@5ý���ٿ�/f����@�>q_��3@qɺ��!?*���4A�@�b ��ٿ�3E����@�3�k��3@�0LLP�!?&'	�4A�@į���ٿ� e����@i���3@�)�Ä�!?Q�f�4A�@唶��ٿ�S?����@�^��3@';�
͐!?�8��4A�@��0d��ٿ�N7����@FQ����3@U'�^�!?���v4A�@��0d��ٿ�N7����@FQ����3@U'�^�!?���v4A�@��0d��ٿ�N7����@FQ����3@U'�^�!?���v4A�@�]ml��ٿ�������@����3@����Ð!?��%{4A�@-����ٿי�����@��L��3@��i��!?�umy4A�@-����ٿי�����@��L��3@��i��!?�umy4A�@-����ٿי�����@��L��3@��i��!?�umy4A�@-����ٿי�����@��L��3@��i��!?�umy4A�@-����ٿי�����@��L��3@��i��!?�umy4A�@G6���ٿ��]����@F�-4��3@0��%
�!?�~�p4A�@G6���ٿ��]����@F�-4��3@0��%
�!?�~�p4A�@4T���ٿ�H����@��Y��3@��:a�!?B�[n4A�@4T���ٿ�H����@��Y��3@��:a�!?B�[n4A�@b�%���ٿC�=����@R����3@mi:�.�!?�(uv4A�@z�ڱ��ٿ�o�����@di��3@95�wu�!?�)w4A�@�oh|��ٿu������@>�����3@�i��5�!?R�u4A�@�$K���ٿS������@>x���3@ ��/�!?xtz4A�@������ٿJ5{����@��oe��3@J#�?<�!?��r4A�@������ٿJ5{����@��oe��3@J#�?<�!?��r4A�@bJR>��ٿܛs����@�ذ���3@Wi�U��!?J��z4A�@��R"��ٿ�ď����@����3@<�R�!?*�x4A�@��R"��ٿ�ď����@����3@<�R�!?*�x4A�@�,`Ʒ�ٿ ^ ����@%���3@��l02�!?��n4A�@�,`Ʒ�ٿ ^ ����@%���3@��l02�!?��n4A�@6X�׹�ٿ/������@{�6���3@߸�k�!?��d4A�@u��O��ٿW������@���~��3@�-O�g�!?�le4A�@��&��ٿ����@�q���3@�����!?��ip4A�@��&��ٿ����@�q���3@�����!?��ip4A�@��&��ٿ����@�q���3@�����!?��ip4A�@_��M��ٿf۶����@�t�#��3@΁���!?�X�i4A�@�@ l��ٿ�X�����@%�79��3@\/�)U�!?�3�l4A�@���Ʊ�ٿ�	�����@��~��3@�)T",�!?���f4A�@�7#��ٿ �����@�z���3@�5���!?ed4A�@Ob P��ٿ��A����@�\���3@X�9?��!?�i4A�@Ob P��ٿ��A����@�\���3@X�9?��!?�i4A�@�ô���ٿ������@|ez���3@H�!|Z�!?��_4A�@׍���ٿ��8����@�	I��3@��@���!?��e4A�@'��&��ٿ9������@���o��3@W4(���!?b�ai4A�@�F�G��ٿ������@�����3@�Nu8�!?��Fb4A�@2v��ٿ�I�����@��i��3@U2AE�!?q�ok4A�@�Yd���ٿIB2����@Fp2���3@j�2%<�!?x�Vg4A�@r~i��ٿڴ���@�sz��3@yb�d�!?VOY4A�@������ٿw�����@%t ���3@,۔�v�!?�DK4A�@��;ٿ&�����@� �`��3@](8DJ�!?\"�M4A�@�����ٿ�iY����@6j��3@��]�!?)��U4A�@OC�м�ٿ������@@Yr���3@��~t[�!?+�3Y4A�@~�S��ٿ�b����@�/���3@��|�s�!?d� d4A�@��۴�ٿ�9�����@6K����3@F4����!?C��s4A�@�]3��ٿ]a�����@
�S���3@ɧ=�d�!?n�?m4A�@��D���ٿ�������@�m�Y��3@�2(Vo�!?ф�j4A�@l��~Ùٿ]ݳ���@s��1��3@��#;q�!?]�^4A�@�ęٿ~#V����@�3K���3@����D�!?Q�a4A�@�ęٿ~#V����@�3K���3@����D�!?Q�a4A�@]ijəٿ�M�����@�����3@!�g�!?���Z4A�@���7Ùٿ�`����@C�����3@�)��!?-h`4A�@���N��ٿv������@�3��3@���!?�Z4A�@�v����ٿ|�H����@h�z��3@ZYSB��!?
�CN4A�@�v����ٿ|�H����@h�z��3@ZYSB��!?
�CN4A�@�v����ٿ|�H����@h�z��3@ZYSB��!?
�CN4A�@K�Ic��ٿU�δ���@�n*��3@r#�Y�!?�60U4A�@�*����ٿ�������@���|��3@y�,N�!?��X4A�@�*����ٿ�������@���|��3@y�,N�!?��X4A�@�*����ٿ�������@���|��3@y�,N�!?��X4A�@�mڕ��ٿ�� ����@�#���3@(Iɼ��!?�]4A�@����ٿm^�����@i�����3@¿��z�!?�>�t4A�@d�����ٿM-H����@�ޕ���3@��<3s�!?�Rq4A�@d�����ٿM-H����@�ޕ���3@��<3s�!?�Rq4A�@S� %��ٿl^�����@������3@1/Y<�!?N��|4A�@S� %��ٿl^�����@������3@1/Y<�!?N��|4A�@S� %��ٿl^�����@������3@1/Y<�!?N��|4A�@]Z'��ٿ� �����@�,���3@�+�!?�1�4A�@�Q4ƥ�ٿ�x�����@y����3@ Bb��!?0K>�4A�@���䧙ٿ�_����@'�e���3@����!?H��4A�@��៙ٿ�����@Y>�c��3@�'�A�!?"/~�4A�@�[[랙ٿxS�����@+-�{��3@OjBSI�!?�׋�4A�@,#�@��ٿ������@*�Q���3@a�)Q]�!?A>�z4A�@T
�e��ٿsl����@Wf���3@�N%�!?���4A�@T
�e��ٿsl����@Wf���3@�N%�!?���4A�@�J�X��ٿP�����@Y}P���3@s�g��!?��}4A�@�J�X��ٿP�����@Y}P���3@s�g��!?��}4A�@�7-��ٿ �e����@2�~7��3@iWM74�!?I�k�4A�@
�g��ٿ-�L����@�r����3@�\%C?�!?
E�4A�@[����ٿ��"����@O����3@���|i�!?i8�x4A�@]q�ݲ�ٿ|�Ⱦ���@�0����3@7�L]E�!?;�v4A�@]q�ݲ�ٿ|�Ⱦ���@�0����3@7�L]E�!?;�v4A�@[.D���ٿg�����@�N���3@s��"�!?a�b4A�@ �_f��ٿ�ρ����@���3@�1)��!?���`4A�@M�����ٿ�E9����@i�����3@��'�!?	�"b4A�@�G Ǚٿ�&����@*�i^��3@�X���!?r�N4A�@��ʙٿg������@{`#��3@�K��;�!?�yUR4A�@H��ʙٿ�����@7�����3@�V�h8�!?���R4A�@bgAVǙٿ� �����@�= ���3@(�k9K�!?Q�O4A�@bgAVǙٿ� �����@�= ���3@(�k9K�!?Q�O4A�@�a2řٿ�6r����@�����3@�-�n�!?O�5S4A�@�h��ٿ\�˳���@����3@��OA�!?�CKQ4A�@@�mf��ٿ$?����@��B���3@��)b�!?A��P4A�@6�&�ʙٿU�٬���@c����3@��L�!?��F4A�@��[D��ٿ!<Z����@�g��3@�cӕ��!?��\4A�@#A[���ٿ��}����@, ��3@5�D���!?I��^4A�@���)��ٿ�~�����@,�R���3@�����!?�Jq4A�@��0
��ٿ8����@��(��3@Y���!?-��~4A�@D����ٿ��a����@g�����3@�3��!?�Ţ4A�@�`I/��ٿa�����@�����3@A͘�Z�!?��*u4A�@���գ�ٿ;�����@^�H���3@� R�!?�=m4A�@���գ�ٿ;�����@^�H���3@� R�!?�=m4A�@�t�ٿ3�����@�׉��3@h���I�!?)�wX4A�@�t�ٿ3�����@�׉��3@h���I�!?)�wX4A�@�t�ٿ3�����@�׉��3@h���I�!?)�wX4A�@=#@(��ٿR�]����@�:����3@�Q� W�!?��^4A�@ ��Խ�ٿ(Bp����@�gM��3@���M�!?��Q4A�@ ��Խ�ٿ(Bp����@�gM��3@���M�!?��Q4A�@�� ��ٿ�9�����@�N���3@8$��\�!?�?�M4A�@~�\��ٿg������@��,��3@M�#�!?H��X4A�@����ٿ�ˌ����@z<���3@V��4�!?�œQ4A�@����ٿ�ˌ����@z<���3@V��4�!?�œQ4A�@����ٿ�ˌ����@z<���3@V��4�!?�œQ4A�@����ٿ�ˌ����@z<���3@V��4�!?�œQ4A�@����ٿ�ˌ����@z<���3@V��4�!?�œQ4A�@S��S��ٿj"�����@<ܚ���3@�hZ�3�!?f*�J4A�@b����ٿ��d����@��5���3@/�A2R�!?:^_F4A�@a�g_ęٿr�@����@.C����3@���G)�!?JP?4A�@ޗ�Ùٿ򤴹���@��3p��3@�`R9�!?	͚E4A�@�H���ٿ�B�����@`u(���3@��b�!?��Z4A�@�H���ٿ�B�����@`u(���3@��b�!?��Z4A�@��B��ٿ'<ߺ���@Cg�<��3@�}IA�!?}�_e4A�@vo{k��ٿ�����@�s����3@+���	�!?&�:L4A�@� ����ٿH������@x����3@(�<؏!?�+�Y4A�@�i�ܬ�ٿj�����@��L��3@19�m��!?/�M4A�@o_)z��ٿٲ�����@�k��3@��vaŏ!?��:4A�@Z�6ʮ�ٿ�zs����@P���3@k��'܏!?	^$4A�@pa3\��ٿ{?Y����@���w��3@ڃ{	�!?q�G4A�@pa3\��ٿ{?Y����@���w��3@ڃ{	�!?q�G4A�@�+�޵�ٿ�8�����@�)���3@���,�!?l�2�3A�@zrƷ�ٿ�����@�k�Z��3@\��t:�!?>��3A�@zrƷ�ٿ�����@�k�Z��3@\��t:�!?>��3A�@躡{��ٿ�������@n�X��3@^��HJ�!?��)4A�@O�h���ٿ�����@A����3@G?a�!?�$+14A�@��1��ٿ��$����@���3@����!?�B	4A�@��1��ٿ��$����@���3@����!?�B	4A�@��1��ٿ��$����@���3@����!?�B	4A�@��1��ٿ��$����@���3@����!?�B	4A�@x����ٿ��Ʀ���@Ϗ0��3@>����!?�V4A�@rɕ[��ٿ������@CO���3@
�D�!?�A4A�@rɕ[��ٿ������@CO���3@
�D�!?�A4A�@�T����ٿ� $����@@1s���3@VɯQ�!?qF&4A�@�T����ٿ� $����@@1s���3@VɯQ�!?qF&4A�@��#���ٿ�ߏ����@p�Wg��3@z��*N�!?��F,4A�@��#���ٿ�ߏ����@p�Wg��3@z��*N�!?��F,4A�@�@���ٿfNv����@\�;���3@�=�c��!?���24A�@�N��ٿ\L�����@"h���3@����q�!?j]-4A�@��빙ٿ>Aɣ���@��s��3@����!?VkoL4A�@�+d��ٿ�Tv����@[ya���3@���]��!?���`4A�@!e���ٿ�K٨���@����3@�*�O�!?Z��r4A�@kT���ٿ|�Ș���@[a>���3@�&3�]�!?B7�V4A�@V4{���ٿ�������@���3@)L�iB�!?Z\4A�@܏��șٿ������@md��3@$�L\@�!?F�؊4A�@܏��șٿ������@md��3@$�L\@�!?F�؊4A�@��񩻙ٿ�Ŕ���@���T��3@;�zI�!?O��A4A�@ݽ����ٿn�!����@�$H���3@������!?�Dp4A�@�Q���ٿ1�}���@n���3@�z_i�!?��24A�@ɬ�C��ٿϬyw���@�/:j��3@=��>�!?�4A�@X�����ٿ�2�����@r���3@oG� ��!?�|��3A�@f-ڜ�ٿ�X�����@o����3@_��!?��3 4A�@1����ٿ�e�����@�x��3@\��!?��M4A�@4�s��ٿ+������@e>����3@Y>X�/�!?84�74A�@4�s��ٿ+������@e>����3@Y>X�/�!?84�74A�@4�s��ٿ+������@e>����3@Y>X�/�!?84�74A�@m򞣙ٿ��-����@],M���3@O=&@�!?�i<4A�@�Yƾ��ٿv�/����@U�7���3@d�^?�!?��F!4A�@�Yƾ��ٿv�/����@U�7���3@d�^?�!?��F!4A�@wb��ٿhW����@��p��3@�ʁh�!?���O4A�@wb��ٿhW����@��p��3@�ʁh�!?���O4A�@k@q��ٿʊޣ���@00�a��3@Bhݔ4�!?��-4A�@��ߚ�ٿ�"�����@Sy���3@ܦ��b�!?�-��3A�@��ߚ�ٿ�"�����@Sy���3@ܦ��b�!?�-��3A�@��Ș��ٿ��Ɠ���@���J��3@b�~j�!?Fj�3A�@3����ٿ�������@8z���3@" Ls�!?�֋�3A�@3����ٿ�������@8z���3@" Ls�!?�֋�3A�@�p|�ٿ�띕���@�1Z��3@��&��!?����3A�@�kH�}�ٿ[rD����@̦�+��3@u�D�+�!?���3A�@�kH�}�ٿ[rD����@̦�+��3@u�D�+�!?���3A�@X�T�m�ٿ �V����@�笟��3@��4V�!?���4A�@89uo�ٿ��d����@�cfe��3@Y/v�S�!?-a��3A�@��⭚�ٿ�������@Y�D^��3@�^��!?j��b4A�@0ި뒙ٿ ������@���
��3@/��:�!?"-��4A�@��r䘙ٿ�k=����@&����3@<
�E�!?��)�4A�@)&!��ٿ������@���\  4@l-�""�!?`��4A�@B�]̙ٿ�Q ��@ٹ~� 4@�F�	5�!?�֢t5A�@�`�'ϙٿ��� ��@��w� 4@u�\�4�!?�X�5A�@i\��ٿ���
 ��@A? 4@�-�_�!?~��5A�@i\��ٿ���
 ��@A? 4@�-�_�!?~��5A�@	s���ٿ��+ ��@|4`� 4@��҉�!?-�0�5A�@�-��ٿ�5 ��@��� 4@�p��2�!?�N@6A�@P���ٿ �8 ��@���� 4@}���;�!?��O�5A�@"�c/�ٿ�)�����@�pB� 4@1�[���!?�Ƴ�5A�@|܂��ٿ7\m ��@EX� 4@�� Db�!? o��5A�@�o��1�ٿ�*� ��@ 4@��me�!?L��R6A�@�o��1�ٿ�*� ��@ 4@��me�!?L��R6A�@�o��1�ٿ�*� ��@ 4@��me�!?L��R6A�@Ŋx��ٿ�Jp����@�cak��3@�b��u�!?����4A�@�<��ٿ�g)����@�f�D��3@�;n=�!?"�=5A�@���陵ٿ�������@�m���3@�F@^�!?���4A�@���N�ٿ���:���@����3@f� A�!?����2A�@)W`�ٿ�()���@C�P��3@)Kh��!?����2A�@�}�s�ٿū�	���@5����3@�D���!?ǿ��2A�@�}�s�ٿū�	���@5����3@�D���!?ǿ��2A�@�}�s�ٿū�	���@5����3@�D���!?ǿ��2A�@�}�s�ٿū�	���@5����3@�D���!?ǿ��2A�@�}�s�ٿū�	���@5����3@�D���!?ǿ��2A�@��8�H�ٿ.�j����@��=��3@�{��z�!?9�I�1A�@��8�H�ٿ.�j����@��=��3@�{��z�!?9�I�1A�@��3_Q�ٿ��z����@�s����3@�0��a�!?���I2A�@<h�g�ٿm�
���@]	����3@�vp�!?r$��2A�@���N�ٿ!����@�B��3@���O�!?��F�1A�@��)V(�ٿV�E����@t�a���3@��1�!?	(�o1A�@0�c��ٿ�"�����@z����3@�$<O$�!?=8@#/A�@0�c��ٿ�"�����@z����3@�$<O$�!?=8@#/A�@��,`ژٿ����@
��Y��3@GM�Yd�!?'F=0A�@w�cl�ٿ��D���@y�����3@���1�!?�Dq�-A�@j�R���ٿ/]�����@#{\��3@qo�kW�!?m��,A�@ ��ٿDe-4���@x<B���3@�ڑFK�!?���	3A�@F_}�y�ٿ#�� ��@���� 4@�H�~�!?��.�7A�@�v�t��ٿ������@�1-���3@q�&��!?E��3A�@NI����ٿj��>���@������3@M�&"1�!?��oI3A�@)X��ٿ+�����@Z�K��3@���0�!?0r[3A�@)X��ٿ+�����@Z�K��3@���0�!?0r[3A�@̶y��ٿ�$�`���@��"S��3@�ϛ?$�!?��.A�@���V�ٿ
lh}���@��0���3@��ڻB�!?�A�1A�@�U�4�ٿ]������@��tI��3@��f�!?e�k�0A�@��+3�ٿ�������@:����3@'�� ��!?�1��/A�@��+3�ٿ�������@:����3@'�� ��!?�1��/A�@��+3�ٿ�������@:����3@'�� ��!?�1��/A�@��+3�ٿ�������@:����3@'�� ��!?�1��/A�@���B�ٿ�_�����@�' ���3@�+w���!?O#/A�@Jz$Z3�ٿG�f� ��@He;� 4@O0���!?9B��6A�@$�;��ٿA����@'r�S# 4@n\��!?V�݋:A�@$�;��ٿA����@'r�S# 4@n\��!?V�݋:A�@7s�͙ٿ�źf ��@n�� 4@����#�!?���5A�@(T�3��ٿ�.T��@��R8 4@�T��b�!?���C<A�@U���ؙٿ}(��@c �C 4@x�5T�!?(a{8A�@U���ؙٿ}(��@c �C 4@x�5T�!?(a{8A�@�rXbi�ٿ��k��@��/Q 4@�
�wx�!?o�6A�@Q�p=E�ٿSJ�����@���:��3@{('ø�!?t��2A�@ŅH�[�ٿ�A>
��@�E?� 4@�(�a��!?� 	�6A�@ŅH�[�ٿ�A>
��@�E?� 4@�(�a��!?� 	�6A�@ŅH�[�ٿ�A>
��@�E?� 4@�(�a��!?� 	�6A�@9n���ٿ-�ob ��@��D� 4@�|az�!?�ܶ5A�@9n���ٿ-�ob ��@��D� 4@�|az�!?�ܶ5A�@��ɺ!�ٿ�b� ��@�w< 4@���U�!?���7A�@��ɺ!�ٿ�b� ��@�w< 4@���U�!?���7A�@��ɺ!�ٿ�b� ��@�w< 4@���U�!?���7A�@)�Hיٿd�
8���@/�{��3@�U��L�!? ,�3A�@i&_���ٿ1�U���@�k���3@���e�!?ɿ�X2A�@�i��ٿ��xg ��@��� 4@Gӻ��!?�}�:8A�@�כٿ��O���@eZ�P 4@:To�!?�3�?A�@��~��ٿ�'4���@�?
X 4@�S����!?��ECBA�@���؝ٿ[.h���@�n��n 4@�/W �!?���FA�@ԯ�r�ٿU�<��@��.K= 4@����!?�n�?AA�@ԯ�r�ٿU�<��@��.K= 4@����!?�n�?AA�@���׸�ٿTҞ'��@cD��R 4@���Q�!?|k#�AA�@�W�+�ٿ.�4���@�d��M 4@�oY8�!?���.BA�@�W�+�ٿ.�4���@�d��M 4@�oY8�!?���.BA�@�W�+�ٿ.�4���@�d��M 4@�oY8�!?���.BA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�\t4�ٿ�*�{��@7%yu 4@���3s�!?�F�_IA�@�O\���ٿ��ԧ��@f� 4@}n�M�!?b+��QA�@�O\���ٿ��ԧ��@f� 4@}n�M�!?b+��QA�@�O\���ٿ��ԧ��@f� 4@}n�M�!?b+��QA�@�O\���ٿ��ԧ��@f� 4@}n�M�!?b+��QA�@�O\���ٿ��ԧ��@f� 4@}n�M�!?b+��QA�@`�GQ*�ٿD�����@���� 4@�=�@�!?Ro��LA�@|5���ٿW�q����@�p?R��3@�+cu]�!?���*"A�@|5���ٿW�q����@�p?R��3@�+cu]�!?���*"A�@�g��A�ٿ����@?�+��3@��9���!?���A�@�g��A�ٿ����@?�+��3@��9���!?���A�@�g��A�ٿ����@?�+��3@��9���!?���A�@]�}/q�ٿ�Rq���@}N���3@�j�h:�!?��!>A�@#*�p�ٿli�K��@�Mv�* 4@�RW{�!?����,A�@#*�p�ٿli�K��@�Mv�* 4@�RW{�!?����,A�@}�F���ٿp�=���@��gV 4@󵻉�!?.�?v=A�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��AU�ٿVTk��@��� 4@;�Ѐ��!?�CA�@��qؖ�ٿyK����@��j+� 4@�7ZB�!?��ߨBA�@��qؖ�ٿyK����@��j+� 4@�7ZB�!?��ߨBA�@�h�鵙ٿA�����@�y|�y 4@��F;�!?a��?A�@�h�鵙ٿA�����@�y|�y 4@��F;�!?a��?A�@�h�鵙ٿA�����@�y|�y 4@��F;�!?a��?A�@�`n�ٿ�A��
��@&�B�� 4@ޥ�3@�!?����GA�@�`n�ٿ�A��
��@&�B�� 4@ޥ�3@�!?����GA�@K�^���ٿ�t7D��@�Sd0� 4@����*�!?��q>A�@K�^���ٿ�t7D��@�Sd0� 4@����*�!?��q>A�@K�^���ٿ�t7D��@�Sd0� 4@����*�!?��q>A�@K�^���ٿ�t7D��@�Sd0� 4@����*�!?��q>A�@ޛ-Z��ٿ�b����@�����4@��b��!?��QA�@ޛ-Z��ٿ�b����@�����4@��b��!?��QA�@ޛ-Z��ٿ�b����@�����4@��b��!?��QA�@ޛ-Z��ٿ�b����@�����4@��b��!?��QA�@Y"�%��ٿq2G���@`w�1V4@[�h���!?8;D�nA�@_�=�ٿ���_��@��#�]4@�m!`�!?��ҾaA�@_�=�ٿ���_��@��#�]4@�m!`�!?��ҾaA�@��Pk�ٿY��-��@�O�6 4@�ku!?h�5A�@�=5�2�ٿ'e����@a.1�j�3@2=.ꕐ!?�Z�m-A�@�=5�2�ٿ'e����@a.1�j�3@2=.ꕐ!?�Z�m-A�@ΒH0�ٿ#����@4i�� 4@�̘�!?�ܳOA�@ΒH0�ٿ#����@4i�� 4@�̘�!?�ܳOA�@ΒH0�ٿ#����@4i�� 4@�̘�!?�ܳOA�@ΒH0�ٿ#����@4i�� 4@�̘�!?�ܳOA�@�?��S�ٿx-����@�G^P� 4@�u�!?��Q;A�@�?��S�ٿx-����@�G^P� 4@�u�!?��Q;A�@�?��S�ٿx-����@�G^P� 4@�u�!?��Q;A�@�?��S�ٿx-����@�G^P� 4@�u�!?��Q;A�@�Ԃ!(�ٿ�&$��@��4@����K�!?F��NA�@����ٿ()���@�O(G� 4@m���z�!?���@A�@����ٿ()���@�O(G� 4@m���z�!?���@A�@����ٿ()���@�O(G� 4@m���z�!?���@A�@����ٿ()���@�O(G� 4@m���z�!?���@A�@����ٿ()���@�O(G� 4@m���z�!?���@A�@R�qxw�ٿߙP^��@%qsK� 4@���fh�!?adC:A�@ͣW�ٿ��Kl��@�-o��4@H���<�!?���NA�@ͣW�ٿ��Kl��@�-o��4@H���<�!?���NA�@ͣW�ٿ��Kl��@�-o��4@H���<�!?���NA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@"��}��ٿSP��
��@eF}�� 4@^�/�Z�!?Ե`5BA�@LÚ�ٿ���d��@��ٺ�4@s_��!?qޘ�HA�@LÚ�ٿ���d��@��ٺ�4@s_��!?qޘ�HA�@LÚ�ٿ���d��@��ٺ�4@s_��!?qޘ�HA�@�HZ ��ٿj�V.��@i��Q!4@DQ��!?�khA�@�HZ ��ٿj�V.��@i��Q!4@DQ��!?�khA�@e��!�ٿ<ݟ���@�*�ا4@7���!?����^A�@e��!�ٿ<ݟ���@�*�ا4@7���!?����^A�@e��!�ٿ<ݟ���@�*�ا4@7���!?����^A�@ �{5��ٿ�Y��"��@3�+4@IyJ�Տ!?�qA�@�0mM��ٿ�_"���@��)�J 4@.�_�Ȑ!?�`�+A�@�0mM��ٿ�_"���@��)�J 4@.�_�Ȑ!?�`�+A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@�Z(�R�ٿ1�	��@!���� 4@b�6�g�!?�r��@A�@��A���ٿ��M���@K����4@{c�d&�!?9\M~fA�@��A���ٿ��M���@K����4@{c�d&�!?9\M~fA�@湳缑ٿ�����@�� �4@��\�y�!?�K��NA�@湳缑ٿ�����@�� �4@��\�y�!?�K��NA�@湳缑ٿ�����@�� �4@��\�y�!?�K��NA�@湳缑ٿ�����@�� �4@��\�y�!?�K��NA�@-C�`ǒٿ�E6���@o���� 4@'ͪq�!?�3]�0A�@-C�`ǒٿ�E6���@o���� 4@'ͪq�!?�3]�0A�@-C�`ǒٿ�E6���@o���� 4@'ͪq�!?�3]�0A�@-C�`ǒٿ�E6���@o���� 4@'ͪq�!?�3]�0A�@-C�`ǒٿ�E6���@o���� 4@'ͪq�!?�3]�0A�@�z:{L�ٿ�*%��@�؟a]�3@���O�!?�cA�@��|E��ٿᱳ7��@'����3@�̼�L�!?�MA�@��|E��ٿᱳ7��@'����3@�̼�L�!?�MA�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@�)��ٿ��[���@kq��3@�+~{�!?-���@�@9�FҔٿ�5����@?�ٗ�3@v�L{��!?��DA�@?���[�ٿ�>$��@�I�n�3@�8�w�!?���A�@?���[�ٿ�>$��@�I�n�3@�8�w�!?���A�@B$���ٿ�����@s��*4@3?RMX�!?Y��HA�@B$���ٿ�����@s��*4@3?RMX�!?Y��HA�@B$���ٿ�����@s��*4@3?RMX�!?Y��HA�@B$���ٿ�����@s��*4@3?RMX�!?Y��HA�@B$���ٿ�����@s��*4@3?RMX�!?Y��HA�@&����ٿD��2��@��p�p�3@Q$����!?�o���@�@2�K��ٿq|�{&��@z�E�4@�H�+�!?�@*�oA�@2�K��ٿq|�{&��@z�E�4@�H�+�!?�@*�oA�@��o�ٿ��N_��@2��n��3@\� 2�!?��aA�@��o�ٿ��N_��@2��n��3@\� 2�!?��aA�@��o�ٿ��N_��@2��n��3@\� 2�!?��aA�@Lد�r�ٿ������@)��D�3@�1��5�!?�xS�/A�@iaU��ٿC�t���@|�v�  4@���i�!?�
J�IA�@cû���ٿ�g+��@l��U��3@1ؓ��!?���A�@cû���ٿ�g+��@l��U��3@1ؓ��!?���A�@cû���ٿ�g+��@l��U��3@1ؓ��!?���A�@����ٿbp`��@,߇]�4@�Z���!?܃��]A�@����ٿbp`��@,߇]�4@�Z���!?܃��]A�@����ٿbp`��@,߇]�4@�Z���!?܃��]A�@����ٿbp`��@,߇]�4@�Z���!?܃��]A�@A���2�ٿ\w��!��@ٯ-��4@��+P�!?|9��oA�@��\���ٿ*�0��@Lw׎�4@D: ,��!?��P`�A�@��\���ٿ*�0��@Lw׎�4@D: ,��!?��P`�A�@��\���ٿ*�0��@Lw׎�4@D: ,��!?��P`�A�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@8��6�ٿ��a��@�c�4@Q���!?>GČPA�@������ٿ%1����@pV-�+�3@�S���!?�|Ձ�@�@������ٿ%1����@pV-�+�3@�S���!?�|Ձ�@�@������ٿ%1����@pV-�+�3@�S���!?�|Ձ�@�@��l�ٿRW�3���@����3@C�">��!?���"�@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@_)���ٿD�1����@`%���3@)|7%@�!?��e@�@�s�`�ٿd��S��@����3@����5�!?�}9A�@�s�`�ٿd��S��@����3@����5�!?�}9A�@�s�`�ٿd��S��@����3@����5�!?�}9A�@�s�`�ٿd��S��@����3@����5�!?�}9A�@�s�`�ٿd��S��@����3@����5�!?�}9A�@�s�`�ٿd��S��@����3@����5�!?�}9A�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@ɗ�t�ٿ�:���@�өҀ�3@m�T���!?$�?ݭ@�@m���ٿs
��@l.I�3@�'�=�!?t�v�A�@m���ٿs
��@l.I�3@�'�=�!?t�v�A�@m���ٿs
��@l.I�3@�'�=�!?t�v�A�@m���ٿs
��@l.I�3@�'�=�!?t�v�A�@m���ٿs
��@l.I�3@�'�=�!?t�v�A�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@mF���ٿ��a���@BT���3@O�ߐ!?�WB6�@�@5j셚ٿ-��Ӈ�@��[�3@�y/�u�!?R�u��@�@5j셚ٿ-��Ӈ�@��[�3@�y/�u�!?R�u��@�@5j셚ٿ-��Ӈ�@��[�3@�y/�u�!?R�u��@�@5j셚ٿ-��Ӈ�@��[�3@�y/�u�!?R�u��@�@*Y|C�ٿ�5����@9�I��3@��l��!?�3�@�@�i��̖ٿ���<���@�
����3@�L�'>�!?'�?�P@�@�i��̖ٿ���<���@�
����3@�L�'>�!?'�?�P@�@�f%śٿ�ŋ����@�}wH�3@�7U u�!?Y7�X�@�@^��?Ýٿ��^	���@K�X���3@���-�!?�gTBC@�@^��?Ýٿ��^	���@K�X���3@���-�!?�gTBC@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@0��)��ٿ�0Qֹ��@�����3@A��%X�!?�o
�@�@t��Pj�ٿ�>Q����@�5	́4@�>V�!?�Ā��@�@R�w�@�ٿ�9ь!��@ʵ�IX�3@J��s�!?�YX^�?�@R�w�@�ٿ�9ь!��@ʵ�IX�3@J��s�!?�YX^�?�@M'J�;�ٿ.%���@X#�8��3@!�ōѐ!?����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@���_��ٿ.k�Aʇ�@S�����3@u�A�E�!?}����@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@T���ٿ������@�P&�3@��Ys9�!?.�ؖ@�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�$\�ٿ��G$��@T֞�4@R󄪐!?��i�A�@�C��ъٿ�����@ĝ\&/4@��w{k�!?$��kA�@ᘯ�!�ٿ�Z�`��@m��l�4@'�3�D�!?:uҤB�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@���ٿ�ܛ��@st\�3@�x�)�!?�4���@�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@K�H�ٿ���0��@�vk�4@n��w�!?���C{A�@��^�6�ٿ����@����&�3@�]���!?$/��@�@��^�6�ٿ����@����&�3@�]���!?$/��@�@��^�6�ٿ����@����&�3@�]���!?$/��@�@��^�6�ٿ����@����&�3@�]���!?$/��@�@��^�6�ٿ����@����&�3@�]���!?$/��@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@H]_-�ٿ��_+��@UT����3@���p�!?M]���@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@����ٿ}�-%���@~��)��3@^�;�[�!?i	&�@�@R�(Y0�ٿ=s�2���@����4@��^�!?)�U�@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�]��ܗٿ��󱵇�@��nH�3@J�1�G�!?��K �@�@�?jL�ٿ8qr�-��@�.�V;�3@q��[�!?��tg�?�@�X��s�ٿ�1ǲ/��@�����3@�fY�C�!?7����?�@�(��Ӕٿ`S��-��@�ji��3@QatM�!?.�s�?�@�(��Ӕٿ`S��-��@�ji��3@QatM�!?.�s�?�@�(��Ӕٿ`S��-��@�ji��3@QatM�!?.�s�?�@�(��Ӕٿ`S��-��@�ji��3@QatM�!?.�s�?�@e<�/��ٿ"䆁��@݇24@�]x#l�!?�i���@�@<#W���ٿ6�X��@�d΋�4@F�.ρ�!?��}~@�@<#W���ٿ6�X��@�d΋�4@F�.ρ�!?��}~@�@<#W���ٿ6�X��@�d΋�4@F�.ρ�!?��}~@�@<#W���ٿ6�X��@�d΋�4@F�.ρ�!?��}~@�@�Q���ٿ��梇�@���J�3@	GA��!?�#��@�@�F ���ٿ�\�_f��@J>����3@׎��O�!?�nI�A�@�Ë�֕ٿ�<�ҙ��@�Y���4@`jrי�!?=Rh,IB�@�Ë�֕ٿ�<�ҙ��@�Y���4@`jrי�!?=Rh,IB�@2_���ٿ!����@�Z@4@A����!?hef�B�@2_���ٿ!����@�Z@4@A����!?hef�B�@2_���ٿ!����@�Z@4@A����!?hef�B�@2_���ٿ!����@�Z@4@A����!?hef�B�@�C| �ٿt����@	0O]H4@T��CȐ!?�3vkB�@�C| �ٿt����@	0O]H4@T��CȐ!?�3vkB�@p0. �ٿ1+��x��@C���7�3@�S��V�!?�-�s�A�@p0. �ٿ1+��x��@C���7�3@�S��V�!?�-�s�A�@p0. �ٿ1+��x��@C���7�3@�S��V�!?�-�s�A�@p0. �ٿ1+��x��@C���7�3@�S��V�!?�-�s�A�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��&�O�ٿ���i��@�F�~�3@�McL�!?���@�@��3�Нٿz b4��@��
��3@��0{�!?sk͈A�@.���ٿ���p��@�I����3@yJ���!?�tC@�@�O���ٿ)�0���@z��'`�3@?�"Z�!?����?�@�O���ٿ)�0���@z��'`�3@?�"Z�!?����?�@�O���ٿ)�0���@z��'`�3@?�"Z�!?����?�@��ߛٿ��ۨ��@�
{d�4@�Bi�!?�(��?�@M	Ŵf�ٿ�b]�#��@奂ϖ�3@cpT8�!?�yIYjA�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@�hK�]�ٿ�Ӷ"���@L���r�3@�>x�3�!?-���o@�@^��ٿ�����@�g�� 4@���吐!?9V��A�@^��ٿ�����@�g�� 4@���吐!?9V��A�@^��ٿ�����@�g�� 4@���吐!?9V��A�@^��ٿ�����@�g�� 4@���吐!?9V��A�@^��ٿ�����@�g�� 4@���吐!?9V��A�@y{��ٿ�j��և�@i_x\��3@+�{G�!?�b���@�@y{��ٿ�j��և�@i_x\��3@+�{G�!?�b���@�@y{��ٿ�j��և�@i_x\��3@+�{G�!?�b���@�@y{��ٿ�j��և�@i_x\��3@+�{G�!?�b���@�@X���R�ٿ�0ud݈�@]�-e�3@�HG*r�!?��C02B�@X���R�ٿ�0ud݈�@]�-e�3@�HG*r�!?��C02B�@�\ʷ,�ٿ=�����@`�6���3@�����!?FjvYj@�@�����ٿ)��<���@���T��3@#I^".�!?��X�@�@�����ٿ)��<���@���T��3@#I^".�!?��X�@�@�����ٿ)��<���@���T��3@#I^".�!?��X�@�@�����ٿ)��<���@���T��3@#I^".�!?��X�@�@�AMH�ٿ\�癆��@�;Dܰ4@K_Sjq�!?s��7�@�@���V�ٿ�~����@r���4@o�*=+�!?��c�8?�@Z+2�~�ٿ�,�W��@C<�"�4@F+�"�!?vW��R@�@Z+2�~�ٿ�,�W��@C<�"�4@F+�"�!?vW��R@�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@>:iŜ�ٿ��I_��@�J~���3@�Fݪ�!?��3/dD�@������ٿJ(�:���@��2��3@�@'��!?;3[�D�@������ٿJ(�:���@��2��3@�@'��!?;3[�D�@������ٿJ(�:���@��2��3@�@'��!?;3[�D�@�3�f�ٿ=���T��@�+��	4@c��K~�!?"���QC�@�3�f�ٿ=���T��@�+��	4@c��K~�!?"���QC�@�3�f�ٿ=���T��@�+��	4@c��K~�!?"���QC�@����T�ٿ�O��c��@o��'z�3@�V��v�!?��
l�E�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@�s��ٿ>G0��@s�p4�3@��m�B�!?����D�@��ܣ�ٿ��\���@��u��3@X��.�!?����G�@��ܣ�ٿ��\���@��u��3@X��.�!?����G�@��ܣ�ٿ��\���@��u��3@X��.�!?����G�@��ܣ�ٿ��\���@��u��3@X��.�!?����G�@�� [��ٿ���_��@h�X��3@�,mL�!?wq�hK�@�� [��ٿ���_��@h�X��3@�,mL�!?wq�hK�@�i�]�ٿ�&�~��@�=��3@�؞���!?���J�@W2�ٿ��3�V��@�E���3@,J朳�!?�D�@۫Q�p�ٿY	��@��d(4@��?���!?b�x�<�@۫Q�p�ٿY	��@��d(4@��?���!?b�x�<�@۫Q�p�ٿY	��@��d(4@��?���!?b�x�<�@۫Q�p�ٿY	��@��d(4@��?���!?b�x�<�@������ٿ�����@aP+ 4@-}�:�!?�E�!D�@������ٿ�����@aP+ 4@-}�:�!?�E�!D�@������ٿ�����@aP+ 4@-}�:�!?�E�!D�@�(���ٿ��_���@���	4@�d�e��!?$��
�J�@�(���ٿ��_���@���	4@�d�e��!?$��
�J�@����g�ٿ|�N_ȑ�@��=c�3@ޥ\
�!?���QO�@��|Y�ٿ_�da��@�^A�v�3@�p��!?_�ѱN�@��|Y�ٿ_�da��@�^A�v�3@�p��!?_�ѱN�@��|Y�ٿ_�da��@�^A�v�3@�p��!?_�ѱN�@l��ʒٿ@2�R��@X����3@9���F�!?;i	!T�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@|�pH�ٿ�9ղޗ�@��K�4@�����!?ģ�==X�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@���
��ٿvq���@�'VL	
4@tm�FO�!?#���V�@-��7�ٿz�{;���@��Ø#4@��J� �!?�>�P�L�@-��7�ٿz�{;���@��Ø#4@��J� �!?�>�P�L�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@Ҥn[
�ٿ�[,��@a�i�3@~��!?��`,7�@�����ٿ��UQ���@W�cu�3@�s�V'�!?[�aG�@�����ٿ��UQ���@W�cu�3@�s�V'�!?[�aG�@�����ٿ��UQ���@W�cu�3@�s�V'�!?[�aG�@�����ٿ��UQ���@W�cu�3@�s�V'�!?[�aG�@�����ٿ��UQ���@W�cu�3@�s�V'�!?[�aG�@7UJJ�ٿ���۹i�@�}ب!�3@s�i��!?�X�c�@7UJJ�ٿ���۹i�@�}ب!�3@s�i��!?�X�c�@7UJJ�ٿ���۹i�@�}ب!�3@s�i��!?�X�c�@ؘ��Y�ٿ{�4��r�@�t�[�4@���um�!?���$�"�@ؘ��Y�ٿ{�4��r�@�t�[�4@���um�!?���$�"�@ؘ��Y�ٿ{�4��r�@�t�[�4@���um�!?���$�"�@ؘ��Y�ٿ{�4��r�@�t�[�4@���um�!?���$�"�@^��p�ٿ&�PT�@��-,�4@�]j�'�!?Yji5���@��*�ٿ���6�@�����	4@b��E4�!?Q�ͥ˶@��*�ٿ���6�@�����	4@b��E4�!?Q�ͥ˶@��*�ٿ���6�@�����	4@b��E4�!?Q�ͥ˶@��*�ٿ���6�@�����	4@b��E4�!?Q�ͥ˶@��*�ٿ���6�@�����	4@b��E4�!?Q�ͥ˶@2�$mߒٿd
R �@�ڔ�,�3@�~o�я!?ز7�|�@2�$mߒٿd
R �@�ڔ�,�3@�~o�я!?ز7�|�@/���R�ٿ0lu:���@$��ƒ�3@��� �!?���r�y�@/���R�ٿ0lu:���@$��ƒ�3@��� �!?���r�y�@/���R�ٿ0lu:���@$��ƒ�3@��� �!?���r�y�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@���Ao�ٿ��̥��@�*OG�3@��HWn�!?d��LWV�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@�uD}�ٿW�5)���@Yd���3@	��~`�!?`I��P�@V_��ٿ7a��kQ�@���z�3@ߧk%�!?>�$���@V_��ٿ7a��kQ�@���z�3@ߧk%�!?>�$���@V_��ٿ7a��kQ�@���z�3@ߧk%�!?>�$���@V_��ٿ7a��kQ�@���z�3@ߧk%�!?>�$���@V_��ٿ7a��kQ�@���z�3@ߧk%�!?>�$���@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@�8UBa�ٿ�����@�/ڽ��3@ia�ȏ!?�����'�@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@d|hI��ٿ۬��Ϊ�@��#n)�3@��x��!?�4�K��@�~_���ٿ:��z�@qVg��3@	��ڐ!?}�C���@�~_���ٿ:��z�@qVg��3@	��ڐ!?}�C���@�~_���ٿ:��z�@qVg��3@	��ڐ!?}�C���@�~_���ٿ:��z�@qVg��3@	��ڐ!?}�C���@�~_���ٿ:��z�@qVg��3@	��ڐ!?}�C���@�d�q��ٿ��(.��@-�6�U�3@�Z@=�!?0MA��K�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@���f�ٿ�7`�L�@}��S4@ ��H$�!?�N�8z�@K����ٿ�bDp�\�@�k"=�3@咅h��!?ѫ�٘�@K����ٿ�bDp�\�@�k"=�3@咅h��!?ѫ�٘�@K����ٿ�bDp�\�@�k"=�3@咅h��!?ѫ�٘�@C�m�"�ٿ=�	����@_��4@�t�p�!?�b�T�u�@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@��¥�ٿӽ��q��@��U�3@ŞM�N�!?5Q���@�C/5�ٿ<�:�z�@VA����3@��P�z�!?"n��=J�@9��l^�ٿ,D�j��@�L����3@�FFc܏!?h] ��@9��l^�ٿ,D�j��@�L����3@�FFc܏!?h] ��@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@sFgޑٿ�a�
g��@�U�c��3@F&nd`�!?9���@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@X�+�ٿ
�)��@*�x�<�3@MN:�b�!?Hh��P��@��7rQ�ٿXƀ���@�cs_�3@`��L�!?vӧ+=�@N�{_ٿcϛ���@�zk�3@��=�H�!?��:��@N�{_ٿcϛ���@�zk�3@��=�H�!?��:��@N�{_ٿcϛ���@�zk�3@��=�H�!?��:��@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@�X�ٿ���`P7�@"ɱq0�3@4��X��!?�y�Z�@+�Aҙٿr0�����@�2�O��3@��t]��!?�{�+�δ@+�Aҙٿr0�����@�2�O��3@��t]��!?�{�+�δ@+�Aҙٿr0�����@�2�O��3@��t]��!?�{�+�δ@+�Aҙٿr0�����@�2�O��3@��t]��!?�{�+�δ@+�Aҙٿr0�����@�2�O��3@��t]��!?�{�+�δ@G����ٿ�T�dIS�@��Fe�3@�eD�i�!?7��Dق�@G����ٿ�T�dIS�@��Fe�3@�eD�i�!?7��Dق�@G����ٿ�T�dIS�@��Fe�3@�eD�i�!?7��Dق�@�Ԥ���ٿ����\v�@�T\P��3@憓�d�!?�v^�C�@�Ԥ���ٿ����\v�@�T\P��3@憓�d�!?�v^�C�@�Ԥ���ٿ����\v�@�T\P��3@憓�d�!?�v^�C�@���q�ٿ�r�!
��@	�5��3@ e��'�!?�z�H0l�@H��s�ٿ]�J#�V�@�G"G*
4@�4\y5�!?H@����@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�u���ٿ�i,#���@�Bf5��3@�Sz�!?>�s�Դ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@�e���ٿ�>�ͤ��@}�D�3@�]H�!?&!P��ȴ@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@}�h6�ٿ�:k�@r�ӹ��3@��t�!?D|�$v2�@q�+�ٿ�P^k �@�53}��3@�#%$A�!?�=ˎ�@q�+�ٿ�P^k �@�53}��3@�#%$A�!?�=ˎ�@q�+�ٿ�P^k �@�53}��3@�#%$A�!?�=ˎ�@q�+�ٿ�P^k �@�53}��3@�#%$A�!?�=ˎ�@q�+�ٿ�P^k �@�53}��3@�#%$A�!?�=ˎ�@P=���ٿ�ȐG�@�Hf9h 4@��K���!?�x{�r�@P=���ٿ�ȐG�@�Hf9h 4@��K���!?�x{�r�@�'F�ٿ)UQty�@���3@�,�4܏!?"�[���@�'F�ٿ)UQty�@���3@�,�4܏!?"�[���@�'F�ٿ)UQty�@���3@�,�4܏!?"�[���@�'F�ٿ)UQty�@���3@�,�4܏!?"�[���@=�o��ٿ���Q��@=R���3@��4��!?��XBp�@���C�ٿeY���D�@3Dd��3@s9��R�!?G,R:2��@�jʠٿmp�;�M�@j�͊��3@
x�F"�!?��2�A{�@�jʠٿmp�;�M�@j�͊��3@
x�F"�!?��2�A{�@+�HjP�ٿ�e��Z�@��L8��3@�y4�ސ!?A���@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@*�Dm_�ٿ9T<�%�@Co����3@_Ä�D�!?~�B�A�@
,���ٿ����.�@l���3@��!?�ܧ]iN�@
,���ٿ����.�@l���3@��!?�ܧ]iN�@
,���ٿ����.�@l���3@��!?�ܧ]iN�@jb�"�ٿ�@#t�@9�Ca�3@���ΐ!?ZIqE��@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@����G�ٿJVRS��@ ��3@��::Ґ!?9�����@h5mɯ�ٿ�9��X�@�.���3@��Iٸ�!?��q����@h5mɯ�ٿ�9��X�@�.���3@��Iٸ�!?��q����@=�c�ٿj1~�s��@Ω�,�3@��Sď!?�](ߴ@=�c�ٿj1~�s��@Ω�,�3@��Sď!?�](ߴ@-Ȭ,�ٿ��ں �@���Bi�3@W���!?`�+�z9�@-Ȭ,�ٿ��ں �@���Bi�3@W���!?`�+�z9�@-Ȭ,�ٿ��ں �@���Bi�3@W���!?`�+�z9�@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@C��yb�ٿ�֕���@#W�k@�3@	�.��!?�XX�ȵ@��Q�ٿ.�����@�2����3@�z���!?'������@��Q�ٿ.�����@�2����3@�z���!?'������@��Q�ٿ.�����@�2����3@�z���!?'������@��Q�ٿ.�����@�2����3@�z���!?'������@��Q�ٿ.�����@�2����3@�z���!?'������@��Q�ٿ.�����@�2����3@�z���!?'������@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@���ݏ�ٿ,e�
��@�0����3@B�+���!?�#�sѴ@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@�s��ٿj6��w��@�����3@��P��!?���Ԯ��@6��p.�ٿY�D��n�@����4@(�]0�!?I�����@���u�ٿGv�8��@ɚ��s�3@|u�c�!?��\��@���u�ٿGv�8��@ɚ��s�3@|u�c�!?��\��@���u�ٿGv�8��@ɚ��s�3@|u�c�!?��\��@�^�q̔ٿX�{��@{e����3@?�C�U�!?X�#3m�@aK��N�ٿ���0��@��O��3@���{��!?h�&�5��@aK��N�ٿ���0��@��O��3@���{��!?h�&�5��@MHO�ٿ�������@�ED*�3@�Ua�Z�!?Py�ϴ@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@���씑ٿ6S*�V�@�//)e�3@�4n_m�!?���n҈�@��j��ٿL��("�@��4߽�3@T���Ґ!?41��<�@*��ޙ�ٿa��s��@Į`�M�3@{_����!?�0�^aֵ@*��ޙ�ٿa��s��@Į`�M�3@{_����!?�0�^aֵ@*��ޙ�ٿa��s��@Į`�M�3@{_����!?�0�^aֵ@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@B��ٿ�c�u�<�@-:���3@ۯ��!?4^��b�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@ȥ����ٿ,%��q	�@,���3@S��!�!?�.�\�@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@����ٿ���X�@dl_���3@v���[�!?�>ė��@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@Z,A��ٿ�D�w���@�g�t��3@��M�h�!?6|��ȵ@N�%��ٿ��VP�@��0��3@���~_�!?����=4�@h��g�ٿ57����@ޠ�9��3@0�H�!?�!���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�V�C�ٿ�$��={�@��~�Z�3@La���!?=�V���@�P�]ؓٿ�	FǇv�@CY��Y�3@\��я!?1���O��@�P�]ؓٿ�	FǇv�@CY��Y�3@\��я!?1���O��@�P�]ؓٿ�	FǇv�@CY��Y�3@\��я!?1���O��@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@F�:"��ٿ��$�P��@X�q�3@	쩶}�!?>�����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@�X��ٿ� o�x�@�����3@�?�_�!?��d����@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@� s�{�ٿ��Ov^%�@�4�)��3@ �p�!?O��=�A�@mz����ٿ�T��@\�	'E�3@��3o�!?@�P��	�@mz����ٿ�T��@\�	'E�3@��3o�!?@�P��	�@mz����ٿ�T��@\�	'E�3@��3o�!?@�P��	�@mz����ٿ�T��@\�	'E�3@��3o�!?@�P��	�@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@.�b�ٿb���'��@�]�I��3@
`��}�!?Ѧ9����@V&�ϗٿ��b��	�@g����3@��j׳�!?�"�͑�@{��^לٿ�pKے��@]!!��3@豨;��!?��ZGCa�@{��^לٿ�pKے��@]!!��3@豨;��!?��ZGCa�@{��^לٿ�pKے��@]!!��3@豨;��!?��ZGCa�@{��^לٿ�pKے��@]!!��3@豨;��!?��ZGCa�@!� 
�ٿD-����@}h�z74@����s�!?7R	�Mh�@!� 
�ٿD-����@}h�z74@����s�!?7R	�Mh�@!� 
�ٿD-����@}h�z74@����s�!?7R	�Mh�@!� 
�ٿD-����@}h�z74@����s�!?7R	�Mh�@e0�Q��ٿT�ŧ21�@���4@��D܏!?T��~R�@e0�Q��ٿT�ŧ21�@���4@��D܏!?T��~R�@e0�Q��ٿT�ŧ21�@���4@��D܏!?T��~R�@e0�Q��ٿT�ŧ21�@���4@��D܏!?T��~R�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@���(�ٿ� \����@�{�s8�3@z�5�!?J��+h�@�,�y�ٿ��}L�@f�� 4@���ŏ!?�u$�<x�@�,�y�ٿ��}L�@f�� 4@���ŏ!?�u$�<x�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�^k�=�ٿ��l���@����g4@Ģ �Q�!?���1:�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@�9B���ٿZ�G��]�@,��3@7�{�h�!?H/��>'�@8�ЙÖٿ�DY��g�@=oV
�3@ݢB�!?w��D1�@8�ЙÖٿ�DY��g�@=oV
�3@ݢB�!?w��D1�@8�ЙÖٿ�DY��g�@=oV
�3@ݢB�!?w��D1�@8�ЙÖٿ�DY��g�@=oV
�3@ݢB�!?w��D1�@8�ЙÖٿ�DY��g�@=oV
�3@ݢB�!?w��D1�@r�����ٿ�6�a��@��@Y�3@��<�!?YP�ݼ�@r�����ٿ�6�a��@��@Y�3@��<�!?YP�ݼ�@r�����ٿ�6�a��@��@Y�3@��<�!?YP�ݼ�@r�����ٿ�6�a��@��@Y�3@��<�!?YP�ݼ�@r�����ٿ�6�a��@��@Y�3@��<�!?YP�ݼ�@<���ʙٿ�b)?��@�d/�|�3@s_��!?�P	�7�@<���ʙٿ�b)?��@�d/�|�3@s_��!?�P	�7�@<���ʙٿ�b)?��@�d/�|�3@s_��!?�P	�7�@<���ʙٿ�b)?��@�d/�|�3@s_��!?�P	�7�@<���ʙٿ�b)?��@�d/�|�3@s_��!?�P	�7�@�ņ�ݛٿ�4�@s�@��>�A�3@ `z1��!?�=ϐ6��@�ņ�ݛٿ�4�@s�@��>�A�3@ `z1��!?�=ϐ6��@�ņ�ݛٿ�4�@s�@��>�A�3@ `z1��!?�=ϐ6��@�ņ�ݛٿ�4�@s�@��>�A�3@ `z1��!?�=ϐ6��@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@����ћٿ)�;��=�@76���3@N��SY�!?�j�D f�@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@���k��ٿ�l�6��@|%�	3�3@i#��F�!?}�C.��@7�8��ٿA5	�'�@w�xF<�3@��4���!?�.V�NI�@7�8��ٿA5	�'�@w�xF<�3@��4���!?�.V�NI�@7�8��ٿA5	�'�@w�xF<�3@��4���!?�.V�NI�@)�N�ޚٿuYe%�@�Q�3@�C�b��!?�ЍW$�@)�N�ޚٿuYe%�@�Q�3@�C�b��!?�ЍW$�@]�2���ٿ�}P�*��@��D��3@X%�⨐!?�((��Ӵ@/�;ʨ�ٿl������@����3@�WȐ!?�2�J��@"۪uD�ٿ�@	�O��@�Q)���3@}��څ�!?�Z�_�ĵ@"۪uD�ٿ�@	�O��@�Q)���3@}��څ�!?�Z�_�ĵ@"۪uD�ٿ�@	�O��@�Q)���3@}��څ�!?�Z�_�ĵ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@�����ٿ'8ް��@X����3@��(�O�!?�if�+ٴ@A��n+�ٿ7���@�[]*�3@�N_���!?O��!�@]ˊ�ٿ ����@V�N�	�3@��c�!?#����@]ˊ�ٿ ����@V�N�	�3@��c�!?#����@]ˊ�ٿ ����@V�N�	�3@��c�!?#����@]ˊ�ٿ ����@V�N�	�3@��c�!?#����@]ˊ�ٿ ����@V�N�	�3@��c�!?#����@.�.���ٿjV죌��@�b"�3@�
��!?��@��@.�.���ٿjV죌��@�b"�3@�
��!?��@��@.�.���ٿjV죌��@�b"�3@�
��!?��@��@��Œ�ٿ�8;+[�@X#!��3@��;��!?�������@��Œ�ٿ�8;+[�@X#!��3@��;��!?�������@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@��3��ٿ�nzc��@F	��3@�?szP�!?��Pu��@]���ٿ�2DQ��@{hOb�3@��:�`�!?+X���@]���ٿ�2DQ��@{hOb�3@��:�`�!?+X���@cCf���ٿ	��%r�@�/54��3@cI>ݏ!?�T�*'��@cCf���ٿ	��%r�@�/54��3@cI>ݏ!?�T�*'��@cCf���ٿ	��%r�@�/54��3@cI>ݏ!?�T�*'��@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@^( `�ٿ��K��"�@HM�)v�3@�0QC�!?�?�{v@�@K�-ɼ�ٿ��h*�*�@��S��	4@�h�Ɛ!?�U��U�@K�-ɼ�ٿ��h*�*�@��S��	4@�h�Ɛ!?�U��U�@f6�\�ٿ�jhP��@/�8\	4@�{����!?@BH��@R�-�b�ٿ��.��@��|4@��]K��!?���>�@R�-�b�ٿ��.��@��|4@��]K��!?���>�@R�-�b�ٿ��.��@��|4@��]K��!?���>�@:bR�ٿE�7>/��@mTv4@t���y�!?=��D)�@���V�ٿ��:~�@Ϋ�
i�3@��Z�!?m)]F�W�@�A,���ٿR?����@��b���3@rL����!?�s-V���@�A,���ٿR?����@��b���3@rL����!?�s-V���@�A,���ٿR?����@��b���3@rL����!?�s-V���@�A,���ٿR?����@��b���3@rL����!?�s-V���@�A,���ٿR?����@��b���3@rL����!?�s-V���@4�C	&�ٿ6��7��@��$���3@e
_7n�!?�Ihm+�@��N�ٿ�Nt���@4�|���3@{�ѐ��!?V=��z�@��N�ٿ�Nt���@4�|���3@{�ѐ��!?V=��z�@��N�ٿ�Nt���@4�|���3@{�ѐ��!?V=��z�@��N�ٿ�Nt���@4�|���3@{�ѐ��!?V=��z�@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@8ҍ�ٿ:4���@FV�E��3@K��a��!?y%�E�Ŵ@0.���ٿɯ�Z4�@��0�K�3@����!?����Z�@0.���ٿɯ�Z4�@��0�K�3@����!?����Z�@I�"l��ٿ_���@y)�ϫ�3@���Jx�!?��!$�@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@����8�ٿ��|��@\����3@X*�kT�!?`-�eӵ@�J���ٿ@�h޻��@U��b��3@���j�!??��'��@�J���ٿ@�h޻��@U��b��3@���j�!??��'��@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@<��_�ٿ|����@0×݌�3@��9�!?<-H�׿�@+"�[�ٿ�k5��*�@� /a�3@���5�!?���8qC�@+"�[�ٿ�k5��*�@� /a�3@���5�!?���8qC�@+"�[�ٿ�k5��*�@� /a�3@���5�!?���8qC�@+"�[�ٿ�k5��*�@� /a�3@���5�!?���8qC�@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@QY�Z�ٿ�1�l��@Jy-P��3@۱�*�!?�Ғ��@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@��l�ʗٿ'���a��@�*�]��3@���!?2ǲ��´@�����ٿb	�U���@* :A\�3@�'}�!?.�R�k��@�����ٿb	�U���@* :A\�3@�'}�!?.�R�k��@�����ٿb	�U���@* :A\�3@�'}�!?.�R�k��@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@�s�D��ٿ1L���@&u�B;�3@�w�2��!?$r6����@���
�ٿ[|��Y�@8B�N�3@G�L�!?4��k��@���
�ٿ[|��Y�@8B�N�3@G�L�!?4��k��@���
�ٿ[|��Y�@8B�N�3@G�L�!?4��k��@���
�ٿ[|��Y�@8B�N�3@G�L�!?4��k��@]�x���ٿ������@�7���3@s�.gy�!? BH
��@]�x���ٿ������@�7���3@s�.gy�!? BH
��@]�x���ٿ������@�7���3@s�.gy�!? BH
��@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@t�1k��ٿȠp�@��3��3@}T��X�!?1zW�@��o��ٿ�?~�n �@���P��3@�c�!?��dϊ�@��o��ٿ�?~�n �@���P��3@�c�!?��dϊ�@��o��ٿ�?~�n �@���P��3@�c�!?��dϊ�@����ߏٿ!+PHa�@<��d�3@<k%3�!?��� �@yt2���ٿ犐��W�@ud����3@b��K�!?�%�.臵@yt2���ٿ犐��W�@ud����3@b��K�!?�%�.臵@yt2���ٿ犐��W�@ud����3@b��K�!?�%�.臵@��%�U�ٿ@TV��@�,5��3@�|ͬ6�!?�kR6޴@��%�U�ٿ@TV��@�,5��3@�|ͬ6�!?�kR6޴@��%�U�ٿ@TV��@�,5��3@�|ͬ6�!?�kR6޴@=�-���ٿ��戃�@۸��r�3@���+�!?|��j��@=�-���ٿ��戃�@۸��r�3@���+�!?|��j��@=�-���ٿ��戃�@۸��r�3@���+�!?|��j��@=�-���ٿ��戃�@۸��r�3@���+�!?|��j��@=�-���ٿ��戃�@۸��r�3@���+�!?|��j��@�2�A�ٿ�7�p���@<�A��3@���\�!?ӷ~��޴@�2�A�ٿ�7�p���@<�A��3@���\�!?ӷ~��޴@�2�A�ٿ�7�p���@<�A��3@���\�!?ӷ~��޴@¯�n��ٿw������@"�?���3@'�|��!?�=;��@¯�n��ٿw������@"�?���3@'�|��!?�=;��@�
�M��ٿp�`�	�@�kq���3@��^��!?��q���@�
�M��ٿp�`�	�@�kq���3@��^��!?��q���@�
�M��ٿp�`�	�@�kq���3@��^��!?��q���@�
�M��ٿp�`�	�@�kq���3@��^��!?��q���@�
�M��ٿp�`�	�@�kq���3@��^��!?��q���@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@a{����ٿG2��@��@M�c�3@ʴ��!?l��A1޴@�X�n�ٿ�B�e/��@�u�>�3@��5B#�!?u5h�
��@��j<ɓٿȬ����@�/���3@����!?\��t˴@��j<ɓٿȬ����@�/���3@����!?\��t˴@��j<ɓٿȬ����@�/���3@����!?\��t˴@��j<ɓٿȬ����@�/���3@����!?\��t˴@tE ��ٿ$E��M��@�fX�f�3@���e�!?�;w;�@tE ��ٿ$E��M��@�fX�f�3@���e�!?�;w;�@��~���ٿꍁ$���@c��v�3@���lV�!?������@>R�)�ٿ��"5��@�a �-�3@���94�!?ol�.ʹ@>R�)�ٿ��"5��@�a �-�3@���94�!?ol�.ʹ@>R�)�ٿ��"5��@�a �-�3@���94�!?ol�.ʹ@�� �8�ٿ��˫%�@M|����3@��Ůя!?~?��U?�@��}E�ٿq1�����@�^�'�3@�Z��׏!?;�Y�͵@�n��*�ٿr/E�h��@�^�q�3@��,��!?Ї#��@�n��*�ٿr/E�h��@�^�q�3@��,��!?Ї#��@�n��*�ٿr/E�h��@�^�q�3@��,��!?Ї#��@�n��*�ٿr/E�h��@�^�q�3@��,��!?Ї#��@tc��G�ٿ�G��@U�,��3@��N�!?��i>yֵ@.���͐ٿ�f���@{���x�3@��mq�!?Q�(�9	�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@�S�ћ�ٿo��#�#�@{@� �3@ܭ+f�!?�]���B�@/�ƈ`�ٿ{��d�!�@
Z�>�3@&i��V�!?
���C�@/�ƈ`�ٿ{��d�!�@
Z�>�3@&i��V�!?
���C�@�Xö�ٿ�`�T��@�Ky��3@h�2�A�!?߄	P�@�Xö�ٿ�`�T��@�Ky��3@h�2�A�!?߄	P�@���>�ٿ	?N�N�@$�7@�3@�����!?k1[yq�@|�XB��ٿU0xX�@נb���3@*�?���!?������@|�XB��ٿU0xX�@נb���3@*�?���!?������@��Z�ٿ� ~I�@��n��3@�� 1��!?��e0P$�@)ĉQ��ٿ8�Z�a��@+�[}��3@v�� �!?~��Ŵ@)ĉQ��ٿ8�Z�a��@+�[}��3@v�� �!?~��Ŵ@)ĉQ��ٿ8�Z�a��@+�[}��3@v�� �!?~��Ŵ@��@�ٿr�b~�I�@��2��3@\��!?�����j�@��@�ٿr�b~�I�@��2��3@\��!?�����j�@��@�ٿr�b~�I�@��2��3@\��!?�����j�@����>�ٿU�PL�/�@�,��\�3@����ʏ!?����xE�@����>�ٿU�PL�/�@�,��\�3@����ʏ!?����xE�@����>�ٿU�PL�/�@�,��\�3@����ʏ!?����xE�@����>�ٿU�PL�/�@�,��\�3@����ʏ!?����xE�@����>�ٿU�PL�/�@�,��\�3@����ʏ!?����xE�@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@7+d�Z�ٿU�]8��@�f<;��3@��#���!?����ȴ@�1?חٿZ���i��@�(�,]4@����Y�!?G%�Bʴ@�1?חٿZ���i��@�(�,]4@����Y�!?G%�Bʴ@5��ٿ,ʶ�ލ�@]c	E�4@?%W�!?��Bz��@5��ٿ,ʶ�ލ�@]c	E�4@?%W�!?��Bz��@5��ٿ,ʶ�ލ�@]c	E�4@?%W�!?��Bz��@�q7�ٿ�>6�@���L4@�IH>�!?�Bܐn�@�q7�ٿ�>6�@���L4@�IH>�!?�Bܐn�@�q7�ٿ�>6�@���L4@�IH>�!?�Bܐn�@�q7�ٿ�>6�@���L4@�IH>�!?�Bܐn�@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@"p0{�ٿ!��:��@�,6ő4@_b�+��!?[Dt���@���GW�ٿ�x����@g�e��3@�>�Rk�!?�U�󆮴@̉�m�ٿ��G棨�@��O!��3@W�;�#�!?�������@̉�m�ٿ��G棨�@��O!��3@W�;�#�!?�������@̉�m�ٿ��G棨�@��O!��3@W�;�#�!?�������@̉�m�ٿ��G棨�@��O!��3@W�;�#�!?�������@̉�m�ٿ��G棨�@��O!��3@W�;�#�!?�������@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@�lBD��ٿ��,����@Q��ɾ�3@YܡM�!?��~W���@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@��R��ٿ�����@eA�R�3@	3B�}�!?�)�#�3�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@�� _��ٿgԁ
�@t�]���3@���0�!?��Xb$�@a'��-�ٿ������@%�@�3@N���N�!?Q! �@a'��-�ٿ������@%�@�3@N���N�!?Q! �@���ޕٿ;S��K�@T�VM��3@��),}�!?��~2h�@���ޕٿ;S��K�@T�VM��3@��),}�!?��~2h�@���ޕٿ;S��K�@T�VM��3@��),}�!?��~2h�@���ޕٿ;S��K�@T�VM��3@��),}�!?��~2h�@���ޕٿ;S��K�@T�VM��3@��),}�!?��~2h�@i�aP�ٿ`��vE�@��?4@�4�#�!?�5��2�@�8�R�ٿ%��!��@�A��4@����d�!?�~���@����ٿ!�(��c�@����3@�o��m�!?�"�-�@����ٿ!�(��c�@����3@�o��m�!?�"�-�@����ٿ!�(��c�@����3@�o��m�!?�"�-�@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@�A5OM�ٿ_���@\hl�3@\�E,�!?tl=���@<g_4ԓٿ�23��1�@y�����3@�#~T�!?�#�e*J�@<g_4ԓٿ�23��1�@y�����3@�#~T�!?�#�e*J�@<g_4ԓٿ�23��1�@y�����3@�#~T�!?�#�e*J�@<g_4ԓٿ�23��1�@y�����3@�#~T�!?�#�e*J�@>
�7x�ٿl�Ţ!�@�Ev �3@v�E*ُ!?��E�@��zN�ٿ��ه^��@O�ah��3@>��;ޏ!?��aQŴ@�p�٧�ٿ��L�@�M�t�3@��7.�!?�����@�p�٧�ٿ��L�@�M�t�3@��7.�!?�����@�p�٧�ٿ��L�@�M�t�3@��7.�!?�����@�p�٧�ٿ��L�@�M�t�3@��7.�!?�����@�p�٧�ٿ��L�@�M�t�3@��7.�!?�����@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@@���-�ٿ|����*�@.k9���3@s���:�!?� y��=�@Z΅�Ɗٿ�j�:N�@D{.c^�3@�l�-�!?v.�(f�@Z΅�Ɗٿ�j�:N�@D{.c^�3@�l�-�!?v.�(f�@Z΅�Ɗٿ�j�:N�@D{.c^�3@�l�-�!?v.�(f�@�y�X։ٿ�)(��@���Ť�3@���k�!?4�˸o��@�y�X։ٿ�)(��@���Ť�3@���k�!?4�˸o��@gF��ٿw�ē��@���t�3@�+�C��!?}��kl´@gF��ٿw�ē��@���t�3@�+�C��!?}��kl´@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@��gNߖٿY�8U%�@���
�3@c$�6��!?���cuX�@�K�_�ٿ-2�s�@Q����3@��K-v�!?�K�);�@�K�_�ٿ-2�s�@Q����3@��K-v�!?�K�);�@�K�_�ٿ-2�s�@Q����3@��K-v�!?�K�);�@�K�_�ٿ-2�s�@Q����3@��K-v�!?�K�);�@�K�_�ٿ-2�s�@Q����3@��K-v�!?�K�);�@��1�0�ٿ�u�5��@Xl`.�4@�2���!?b�>��ܴ@j�-C��ٿW�1����@���� 4@�/9�!?~[�V;�@j�-C��ٿW�1����@���� 4@�/9�!?~[�V;�@j�-C��ٿW�1����@���� 4@�/9�!?~[�V;�@j�-C��ٿW�1����@���� 4@�/9�!?~[�V;�@���{�ٿR�o����@x.+I��3@B9�W�!?�M�%��@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@��.���ٿ!�Z��(�@�g���3@�I�aM�!?}�����@pb�>�ٿE�Tb}��@�l��3@-<����!?J�8�qK�@����ٿ$R��eU�@Z�g�3@��	�!?|���(��@����ٿ$R��eU�@Z�g�3@��	�!?|���(��@(9E�ٿS�zNp��@�;;�3@e��!L�!?1Sy�Rs�@{� 3��ٿ/�f̗��@�����3@��N�!?��L!�"�@{� 3��ٿ/�f̗��@�����3@��N�!?��L!�"�@{� 3��ٿ/�f̗��@�����3@��N�!?��L!�"�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@L&]cĖٿ9wz�V��@ܐ̄�3@�<d�,�!?J�	�T�@D����ٿ�N#����@9ǻ$��3@'-�R3�!?�`��@D����ٿ�N#����@9ǻ$��3@'-�R3�!?�`��@���}��ٿ���+��@��I*��3@���R�!?�%����@�#N|�ٿ3���ޮ�@�)掞�3@,}9�!?{���S�@�#N|�ٿ3���ޮ�@�)掞�3@,}9�!?{���S�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@��=���ٿ�:|�_��@�jv���3@֕X�!?4��|L7�@H#��ٿ��W�p��@O�����3@.Se}�!?��*n���@tHFd�ٿ�{�E��@U��A�3@.�ն[�!?�Id��<�@`5���ٿ��B���@:S ��3@X�(w�!?;�����@`5���ٿ��B���@:S ��3@X�(w�!?;�����@`5���ٿ��B���@:S ��3@X�(w�!?;�����@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@�u���ٿ��G9:��@	eX�C�3@n�2L�!?d�gAv�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@m���ڕٿy(��<��@��
�d�3@��<��!?�xv�}�@���?P�ٿmn��9|�@ �;�(�3@5M> *�!?��쀛�@�~^�ٿ������@�Ư�	�3@	BfM�!?��x1��@�~^�ٿ������@�Ư�	�3@	BfM�!?��x1��@�~^�ٿ������@�Ư�	�3@	BfM�!?��x1��@ݾ��ٿ�-/��@���g��3@�e��P�!?����@ݾ��ٿ�-/��@���g��3@�e��P�!?����@ݾ��ٿ�-/��@���g��3@�e��P�!?����@ݾ��ٿ�-/��@���g��3@�e��P�!?����@��@�ٿ�@�8��@΁J �3@5>�[�!?���{ |�@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@���᪓ٿ�(;����@��-\��3@"7]��!?���4˴@G6׵��ٿҰfZG�@�ۙެ�3@1Xjt��!?��?��@G6׵��ٿҰfZG�@�ۙެ�3@1Xjt��!?��?��@G6׵��ٿҰfZG�@�ۙެ�3@1Xjt��!?��?��@G6׵��ٿҰfZG�@�ۙެ�3@1Xjt��!?��?��@����ٿ}�� �@� �r�3@��!��!?�-D�3�@����ٿ}�� �@� �r�3@��!��!?�-D�3�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@O��s��ٿ<��&�l�@z#��3@�j�"��!?�-Z_�@@P�T�ٿy;݁-�@�}T?�4@���>�!?���
��@@P�T�ٿy;݁-�@�}T?�4@���>�!?���
��@@P�T�ٿy;݁-�@�}T?�4@���>�!?���
��@3�� �ٿ1�8r���@���4@�CQ���!?��dA�@3�� �ٿ1�8r���@���4@�CQ���!?��dA�@3�� �ٿ1�8r���@���4@�CQ���!?��dA�@3�� �ٿ1�8r���@���4@�CQ���!?��dA�@3�� �ٿ1�8r���@���4@�CQ���!?��dA�@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�_e��ٿ�N�@�9�M{4@�Wx��!?���M��@�����ٿ�5�4��@��V�64@�|d1�!?�_�j�#�@�����ٿ�5�4��@��V�64@�|d1�!?�_�j�#�@�����ٿ�5�4��@��V�64@�|d1�!?�_�j�#�@�����ٿ�5�4��@��V�64@�|d1�!?�_�j�#�@������ٿ�K;�wu�@C��
4@tmg �!?F�+�r��@������ٿ�K;�wu�@C��
4@tmg �!?F�+�r��@�(��ٿ��<@��@k��M�4@����!?�e��H�@�(��ٿ��<@��@k��M�4@����!?�e��H�@�(��ٿ��<@��@k��M�4@����!?�e��H�@�(��ٿ��<@��@k��M�4@����!?�e��H�@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@�^K��ٿ�S����@�ò(�3@�Ր~W�!?�*�p��@��8�H�ٿ݂Ϊ9�@q7����3@þ&g�!?jI_���@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@�Qں�ٿR��VP�@&���p�3@{��N�!?D�3
Vʴ@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@YHwN?�ٿFLమ��@�㸗�3@ZS�?�!?��d���@x$b"��ٿ���qN�@hJ�F.�3@y%W���!?dam�@q�����ٿ������@V�����3@%����!?5H��L��@�̆�ːٿ������@&���i 4@&ݟǸ�!?6NN��b�@�̆�ːٿ������@&���i 4@&ݟǸ�!?6NN��b�@�L�*�ٿ�ӓ���@|S>�Z�3@��~��!?�t�ʹ@�L�*�ٿ�ӓ���@|S>�Z�3@��~��!?�t�ʹ@�L�*�ٿ�ӓ���@|S>�Z�3@��~��!?�t�ʹ@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@�b�ٿ(��	���@f�+ړ�3@|RR��!?�6I�?�@ˢ�Z2�ٿ�xF�2K�@A��Ou�3@�[|!p�!?�ƞR%t�@ˢ�Z2�ٿ�xF�2K�@A��Ou�3@�[|!p�!?�ƞR%t�@ˢ�Z2�ٿ�xF�2K�@A��Ou�3@�[|!p�!?�ƞR%t�@ˢ�Z2�ٿ�xF�2K�@A��Ou�3@�[|!p�!?�ƞR%t�@�(a$�ٿ������@Z|F��3@�`�`'�!?�j7Hд@�(a$�ٿ������@Z|F��3@�`�`'�!?�j7Hд@�(a$�ٿ������@Z|F��3@�`�`'�!?�j7Hд@�zȅ�ٿ��#*aH�@39����3@�U��!?X�לum�@�zȅ�ٿ��#*aH�@39����3@�U��!?X�לum�@��f�֛ٿL 2����@�	F�i�3@(c��6�!?��٩�@��f�֛ٿL 2����@�	F�i�3@(c��6�!?��٩�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@���Γٿn�
SI�@F�k}��3@C�9z	�!?�S��~�@��s2�ٿ�~�͖)�@^���X�3@�:N@j�!?��B�@�l�sٖٿ	�U��@��,km�3@C�+�!?�oةa��@�l�sٖٿ	�U��@��,km�3@C�+�!?�oةa��@�l�sٖٿ	�U��@��,km�3@C�+�!?�oةa��@�l�sٖٿ	�U��@��,km�3@C�+�!?�oةa��@LsG���ٿ�����@,����3@�2H
�!?�ٝA�@LsG���ٿ�����@,����3@�2H
�!?�ٝA�@LsG���ٿ�����@,����3@�2H
�!?�ٝA�@LsG���ٿ�����@,����3@�2H
�!?�ٝA�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@��i�i�ٿV/���@HQ���3@_Oo�!?�[�G7�@9-�3N�ٿ��A4���@�4��3@sG����!?�
�ܫM�@9-�3N�ٿ��A4���@�4��3@sG����!?�
�ܫM�@9-�3N�ٿ��A4���@�4��3@sG����!?�
�ܫM�@9-�3N�ٿ��A4���@�4��3@sG����!?�
�ܫM�@9-�3N�ٿ��A4���@�4��3@sG����!?�
�ܫM�@-���ٿ>��M [�@Ǧ�̩�3@�)#`�!?`��t�@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@f��c9�ٿd���8�@@�#xj�3@<���!?<֥@;���t�ٿJ�S����@��5��4@��^��!?����Ǵ@;���t�ٿJ�S����@��5��4@��^��!?����Ǵ@;���t�ٿJ�S����@��5��4@��^��!?����Ǵ@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@�j�ݞٿrf�'O�@�AP���3@�4]�!?���C˴@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@i�V8�ٿ{_���k�@�6��3@;'� k�!?�ߞ"�@���t��ٿ�~��h�@����3@,+���!?8&��)�@1M����ٿ�B� �@^�Y(��3@�G/���!?�� δ@1M����ٿ�B� �@^�Y(��3@�G/���!?�� δ@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@Ü�:��ٿ�G�ZuK�@���3@�-�L�!?�
����@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@�0��(�ٿ�'>F���@a%���3@�x*E�!?/�?#��@2 ��ٿժ�����@����3@���]G�!?u��,��@2 ��ٿժ�����@����3@���]G�!?u��,��@2 ��ٿժ�����@����3@���]G�!?u��,��@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@�6��ٿ��K��t�@�bxby�3@J�ɏF�!?�l|?!f�@l���ߖٿP8&�@P�����3@>6�"�!?_U�sH{�@l���ߖٿP8&�@P�����3@>6�"�!?_U�sH{�@l���ߖٿP8&�@P�����3@>6�"�!?_U�sH{�@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@�keR�ٿ"	eE�q�@2����4@m_�1I�!?yT��@O���ٿ@��8��@���d��3@���U�!?b�'_�@F�K`D�ٿk�k�K�@IQR��3@�"M�!?�_�¾E�@F�K`D�ٿk�k�K�@IQR��3@�"M�!?�_�¾E�@F�K`D�ٿk�k�K�@IQR��3@�"M�!?�_�¾E�@';�ݯ�ٿ�HSU���@��@�M�3@�� �!?����Ѵ@';�ݯ�ٿ�HSU���@��@�M�3@�� �!?����Ѵ@�B�ė�ٿ�Ev����@��c��3@k<�	D�!?���܎��@�B�ė�ٿ�Ev����@��c��3@k<�	D�!?���܎��@�B�ė�ٿ�Ev����@��c��3@k<�	D�!?���܎��@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@g����ٿ������@������3@���u�!?l���@���W<�ٿ�{j�4�@��I`�3@h��e�!?Vt�.���@�ϵbh�ٿ�:��@�]'�3@���DH�!?G�+�@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@I��w�ٿ$�JA���@���~��3@�.�/�!?���R$��@��W��ٿ�;��K�@�6s{X�3@7�2C�!?1�8E�{�@��W��ٿ�;��K�@�6s{X�3@7�2C�!?1�8E�{�@��W��ٿ�;��K�@�6s{X�3@7�2C�!?1�8E�{�@��W��ٿ�;��K�@�6s{X�3@7�2C�!?1�8E�{�@��W��ٿ�;��K�@�6s{X�3@7�2C�!?1�8E�{�@�S�w��ٿ�r��@�z�$��3@t:��C�!?)��J2:�@�S�w��ٿ�r��@�z�$��3@t:��C�!?)��J2:�@�S�w��ٿ�r��@�z�$��3@t:��C�!?)��J2:�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�Z���ٿ�ز4���@��#��3@;_G�!?�V��b@�@�v�D�ٿ���[D��@��ͻ��3@j��9��!?Y���R�@�v�D�ٿ���[D��@��ͻ��3@j��9��!?Y���R�@�v�D�ٿ���[D��@��ͻ��3@j��9��!?Y���R�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@���z|�ٿnT�#��@�����3@�w@�X�!?��m'�K�@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@E8c��ٿ"�h����@�����3@"��0�!?k'r��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@"C���ٿ�Xt��@�@�8*��3@�I��?�!?[EN��@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@����ٿ�"���B�@����k�3@ѤxX�!?�`FY���@��n�p�ٿXu�^�@�a{#��3@7�wA�!?0FD��+�@��n�p�ٿXu�^�@�a{#��3@7�wA�!?0FD��+�@��n�p�ٿXu�^�@�a{#��3@7�wA�!?0FD��+�@��n�p�ٿXu�^�@�a{#��3@7�wA�!?0FD��+�@i�l�{�ٿ��g�� �@��J-�3@��`�e�!?7���Y�@�L��R�ٿ�O���+�@�w0�?4@񌎕�!?"��'Ŵ@T����ٿ�nCh���@�G׋3�3@֪���!?�p�´@����ٿ�BZ����@�(���3@C��vD�!?�s�lAŴ@����ٿ�BZ����@�(���3@C��vD�!?�s�lAŴ@��j^�ٿ���X��@�o��3@�m��-�!?�] �,Z�@��j^�ٿ���X��@�o��3@�m��-�!?�] �,Z�@��j^�ٿ���X��@�o��3@�m��-�!?�] �,Z�@���ǕٿM���8s�@�*���3@˹�,�!?vW�t�3�@���ǕٿM���8s�@�*���3@˹�,�!?vW�t�3�@���ǕٿM���8s�@�*���3@˹�,�!?vW�t�3�@���ǕٿM���8s�@�*���3@˹�,�!?vW�t�3�@������ٿ�`�F��@��X� 4@̱�B6�!?���.$�@������ٿ�`�F��@��X� 4@̱�B6�!?���.$�@������ٿ�`�F��@��X� 4@̱�B6�!?���.$�@������ٿ�`�F��@��X� 4@̱�B6�!?���.$�@������ٿ�`�F��@��X� 4@̱�B6�!?���.$�@������ٿ�[�N[��@�D��4@\i�A�!?u��|D�@������ٿ�[�N[��@�D��4@\i�A�!?u��|D�@������ٿ�[�N[��@�D��4@\i�A�!?u��|D�@�q�E�ٿl1Mݖ�@C��S�3@��;	B�!?��~�UD�@�q�E�ٿl1Mݖ�@C��S�3@��;	B�!?��~�UD�@�q�E�ٿl1Mݖ�@C��S�3@��;	B�!?��~�UD�@�n�~�ٿP�|40��@A�N���3@�ϣW�!?�v���
�@�n�~�ٿP�|40��@A�N���3@�ϣW�!?�v���
�@�n�~�ٿP�|40��@A�N���3@�ϣW�!?�v���
�@�n�~�ٿP�|40��@A�N���3@�ϣW�!?�v���
�@K$w=�ٿ7���)��@�� Ќ�3@�aAgz�!?+��.�z�@K$w=�ٿ7���)��@�� Ќ�3@�aAgz�!?+��.�z�@K$w=�ٿ7���)��@�� Ќ�3@�aAgz�!?+��.�z�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@(�Z�S�ٿkbc����@�ذ��3@�sZ�!?��!Էj�@ZTm��ٿZ��]j�@��+�v�3@���WI�!?t�GqMf�@&0��6�ٿt-.��`�@�93��3@�nd4%�!?��|�3�@&0��6�ٿt-.��`�@�93��3@�nd4%�!?��|�3�@&0��6�ٿt-.��`�@�93��3@�nd4%�!?��|�3�@J+�Wŕٿ ɏs�@}"�V0�3@�Z�3�!?��^$�n�@J+�Wŕٿ ɏs�@}"�V0�3@�Z�3�!?��^$�n�@J+�Wŕٿ ɏs�@}"�V0�3@�Z�3�!?��^$�n�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@�m���ٿ��G*E�@y�9�3@���
K�!?1ܞ�y�@s�3cזٿ��w8ѡ�@����j�3@)��aL�!?�0��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@T���'�ٿ�̱�&��@ʣN2\�3@���xP�!?����{��@Y�<�p�ٿ�u��@��7���3@Q3�|u�!?��ā"��@����ٿ�̘��@�G>�
�3@j���?�!?��9@�@����ٿ�̘��@�G>�
�3@j���?�!?��9@�@����ٿ�̘��@�G>�
�3@j���?�!?��9@�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@7q����ٿ"-�)ҿ@2�����3@$���Z�!?����P�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@�
jޥ�ٿ�uc:���@�-Ď�3@Io�q�!?����_�@��SG�ٿ64A�F��@�y��4@Y\/\5�!?z�$]��@��SG�ٿ64A�F��@�y��4@Y\/\5�!?z�$]��@��SG�ٿ64A�F��@�y��4@Y\/\5�!?z�$]��@h�BNȘٿ�� ��@�@���w�3@����!?���P�@h�BNȘٿ�� ��@�@���w�3@����!?���P�@h�BNȘٿ�� ��@�@���w�3@����!?���P�@V���m�ٿLѼX�@ٰQ-��3@�/���!?�o�k�@V���m�ٿLѼX�@ٰQ-��3@�/���!?�o�k�@V���m�ٿLѼX�@ٰQ-��3@�/���!?�o�k�@��d�_�ٿ��El$�@ZDVɆ�3@�%k��!?��o��@��뇘ٿ�'�~��@zidX3�3@%�l�!?��^��B�@��뇘ٿ�'�~��@zidX3�3@%�l�!?��^��B�@�Y�O��ٿ�m�����@�*�]��3@k]�#
�!?����@�Y�O��ٿ�m�����@�*�]��3@k]�#
�!?����@�Y�O��ٿ�m�����@�*�]��3@k]�#
�!?����@�Y�O��ٿ�m�����@�*�]��3@k]�#
�!?����@�Y�O��ٿ�m�����@�*�]��3@k]�#
�!?����@�2+�	�ٿX�����@�j�>�3@>d�9�!?C8��@���9j�ٿ��}\x�@�;���3@�J��!?�4����@���9j�ٿ��}\x�@�;���3@�J��!?�4����@iȹFy�ٿ�7�i�@W�T�3@`�|"X�!?�hi�/�@���ٿ���R��@{d_��3@n�
��!?�iG��E�@���ٿ���R��@{d_��3@n�
��!?�iG��E�@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@�T�n�ٿ:o���*�@e��+�3@�zW��!?2nfL��@8����ٿ��ϯ�@�85S�3@������!?,֒E[�@8����ٿ��ϯ�@�85S�3@������!?,֒E[�@8����ٿ��ϯ�@�85S�3@������!?,֒E[�@8����ٿ��ϯ�@�85S�3@������!?,֒E[�@8����ٿ��ϯ�@�85S�3@������!?,֒E[�@�.���ٿ�z"֊w�@-7����3@&��^t�!?���M�@�.���ٿ�z"֊w�@-7����3@&��^t�!?���M�@�2�Q��ٿL1R�r�@�
����3@��S ]�!?R5q �x�@9y���ٿ
5�,���@�����3@�	�|�!?M�7n�m�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@Ӻ5��ٿZP�-�@S}p_��3@u�Pu;�!?u��5�@ז\��ٿ�
��P��@uoLZ�3@�[�(��!?��z^���@ז\��ٿ�
��P��@uoLZ�3@�[�(��!?��z^���@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@z�m���ٿ���~�@������3@�S|"��!?B���r�@�ps�>�ٿ�f�^��@�b@�G�3@%K�T7�!?Xu�l�@Xfɋc�ٿ�Ԛ:^�@���3@b���^�!?�!T ���@Xfɋc�ٿ�Ԛ:^�@���3@b���^�!?�!T ���@��^@�ٿ��:���@w3O��3@Y:sS�!?w�,�@��^@�ٿ��:���@w3O��3@Y:sS�!?w�,�@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@Q�֯��ٿ�ֹ�@���2�3@�VK�b�!?K�Oa��@��&Øٿ�"wO�@�����3@�ج<�!?>A<V�@��&Øٿ�"wO�@�����3@�ج<�!?>A<V�@��&Øٿ�"wO�@�����3@�ج<�!?>A<V�@��&Øٿ�"wO�@�����3@�ج<�!?>A<V�@R^5�ٿ�5���@�/x,��3@�';��!?�6�%�E�@R^5�ٿ�5���@�/x,��3@�';��!?�6�%�E�@R^5�ٿ�5���@�/x,��3@�';��!?�6�%�E�@R^5�ٿ�5���@�/x,��3@�';��!?�6�%�E�@j�Q0�ٿ��C�:��@JK����3@t	�q%�!?03��(�@j�Q0�ٿ��C�:��@JK����3@t	�q%�!?03��(�@&���M�ٿ�i[N7L�@(@�}�3@�1��!?��8q$2�@&���M�ٿ�i[N7L�@(@�}�3@�1��!?��8q$2�@&���M�ٿ�i[N7L�@(@�}�3@�1��!?��8q$2�@᝿Xؓٿ� ��F��@M�{�2�3@S?V=�!?r�ez��@᝿Xؓٿ� ��F��@M�{�2�3@S?V=�!?r�ez��@���ِٿ�Y�Ay��@�����3@͛���!?��7��@���ِٿ�Y�Ay��@�����3@͛���!?��7��@���ِٿ�Y�Ay��@�����3@͛���!?��7��@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@{�/r�ٿ��y�3>�@�Q����3@*V+��!?ӊq�W�@./>=Q�ٿ�@瞔k�@C3=ޔ�3@vU�tp�!?�����"�@./>=Q�ٿ�@瞔k�@C3=ޔ�3@vU�tp�!?�����"�@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@{�_��ٿ �nt^�@bI�s��3@우N1�!?��*�Ĵ@=`�(�ٿ(����&�@�Զv��3@�tBP�!?��l޴@=`�(�ٿ(����&�@�Զv��3@�tBP�!?��l޴@=`�(�ٿ(����&�@�Զv��3@�tBP�!?��l޴@=`�(�ٿ(����&�@�Զv��3@�tBP�!?��l޴@=`�(�ٿ(����&�@�Զv��3@�tBP�!?��l޴@8���Ȝٿ�_Β��@rh���3@Z��BN�!?�'+���@8���Ȝٿ�_Β��@rh���3@Z��BN�!?�'+���@8���Ȝٿ�_Β��@rh���3@Z��BN�!?�'+���@8���Ȝٿ�_Β��@rh���3@Z��BN�!?�'+���@��6��ٿ�^�L���@43�Q�3@�E]�}�!?!N#���@ _{�(�ٿ	Ag�k��@n�.��3@�-,���!?�ۋ.��@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@u�Ƨ��ٿC	�C��@I�3_�3@��n�ԏ!?Ll�1�@(��ۓٿz�9dy��@�vP��3@�Ie�]�!?�Xyw�S�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@����`�ٿ)����@,�v�s�3@ @
)��!?���d9�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@��n�P�ٿ���}�@Ϯ�/��3@�V¬�!?��G<Z:�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@u�N��ٿ�����!�@̢�K�3@�"��R�!?��%�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@�c�ٿ��ٺ09�@�|#��3@xAU_�!?	�o�>�@_J��z�ٿO��l���@���qx�3@>��3�!?ɤ䝝t�@_J��z�ٿO��l���@���qx�3@>��3�!?ɤ䝝t�@-�����ٿԻ���9�@)�b��3@�P�n�!?R���뽵@~`S̔ٿ/�{k���@g"k��3@Y�nf:�!?o5�ɣ�@od@?��ٿ\14g�O�@%CJ
�3@/r���!?k��{b/�@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@>&R =�ٿ��P�%�@�"^w�3@_��
�!?[W�@��@&�{-�ٿ˷�����@ͷ���3@�n�5�!?s��e�h�@&�{-�ٿ˷�����@ͷ���3@�n�5�!?s��e�h�@�(˽�ٿ���H�&�@�����3@?I��?�!?�h�D��@�(˽�ٿ���H�&�@�����3@?I��?�!?�h�D��@��̚ٿ��I)<�@�ʁ��3@q~�R&�!?;���7E�@��̚ٿ��I)<�@�ʁ��3@q~�R&�!?;���7E�@��̚ٿ��I)<�@�ʁ��3@q~�R&�!?;���7E�@��̚ٿ��I)<�@�ʁ��3@q~�R&�!?;���7E�@w=9K/�ٿ,s?�V�@݁��3@7��x�!?�^����@w=9K/�ٿ,s?�V�@݁��3@7��x�!?�^����@u+�|-�ٿ_E�Ph�@"\w�8�3@� >��!?6�4�R$�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@��n�ٿ���crz�@�]�D�3@�yOAJ�!?����ަ�@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@L�PMG�ٿ�ۛ�{�@*?��l�3@sr�o�!?'�S��̵@�#)�ȗٿ�.Bk��@̅~G4@��C�h�!?[j@���@�#)�ȗٿ�.Bk��@̅~G4@��C�h�!?[j@���@�#)�ȗٿ�.Bk��@̅~G4@��C�h�!?[j@���@�#)�ȗٿ�.Bk��@̅~G4@��C�h�!?[j@���@�#)�ȗٿ�.Bk��@̅~G4@��C�h�!?[j@���@u���ǖٿ��v=?�@.�'RD 4@ь��f�!?���ꤵ@u���ǖٿ��v=?�@.�'RD 4@ь��f�!?���ꤵ@u���ǖٿ��v=?�@.�'RD 4@ь��f�!?���ꤵ@u���ǖٿ��v=?�@.�'RD 4@ь��f�!?���ꤵ@u���ǖٿ��v=?�@.�'RD 4@ь��f�!?���ꤵ@�wq��ٿ+e��Ц�@�s�_��3@��}"y�!?����x��@������ٿC}cj}D�@��!�3@��m��!?���>:˴@������ٿC}cj}D�@��!�3@��m��!?���>:˴@������ٿC}cj}D�@��!�3@��m��!?���>:˴@������ٿC}cj}D�@��!�3@��m��!?���>:˴@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@�˪�C�ٿ���l�@&2z�<�3@�vP�7�!?/���ܴ@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@9�p�Ôٿ�v�p�@�ڮ��3@o@�y�!?��;~�O�@)8�3��ٿܣ�r�@�E-�3@��:�)�!?KeD���@)8�3��ٿܣ�r�@�E-�3@��:�)�!?KeD���@�ͦ��ٿ����@� ���3@�_Z�b�!?�
��@,�?�S�ٿ:�Q3;�@Akn��3@
F���!?�H����@�� z5�ٿec6���@��\��3@5o�O\�!?�a�t|��@�� z5�ٿec6���@��\��3@5o�O\�!?�a�t|��@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@�*��əٿzRjæ��@M�����3@�$tOI�!?c����"�@f���͛ٿUq��zx�@��5���3@��V��!?�ұZ��@?eU,A�ٿ�bxa���@rE��k�3@V�8.�!?�T��A��@(*��$�ٿ���H�@����3@��=�e�!?������@(*��$�ٿ���H�@����3@��=�e�!?������@(*��$�ٿ���H�@����3@��=�e�!?������@Jxq�7�ٿR¯�o]�@;�L<��3@��l��!?j�9��@�R�HĔٿ*��}��@GXuY4@e��HK�!?��+�"�@�R�HĔٿ*��}��@GXuY4@e��HK�!?��+�"�@�R�HĔٿ*��}��@GXuY4@e��HK�!?��+�"�@�lƄ�ٿ�4���@�J�� 4@J���!?�\xm%�@Ҁaaؑٿ�=C'�@W�F�^�3@L`R.�!?�b\δ@Ҁaaؑٿ�=C'�@W�F�^�3@L`R.�!?�b\δ@Ҁaaؑٿ�=C'�@W�F�^�3@L`R.�!?�b\δ@Ҁaaؑٿ�=C'�@W�F�^�3@L`R.�!?�b\δ@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@���\�ٿ�*ez��@a�F�c�3@t��Vj�!?BK�@ii���ٿ�Q�[
��@��Ko�3@���"�!?������@ii���ٿ�Q�[
��@��Ko�3@���"�!?������@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@ir7v��ٿ)�52���@}�$���3@�DD[)�!?��ڮ��@���^��ٿi�8.W��@��1Y6�3@&��!?�ݗ���@���^��ٿi�8.W��@��1Y6�3@&��!?�ݗ���@���^��ٿi�8.W��@��1Y6�3@&��!?�ݗ���@���^��ٿi�8.W��@��1Y6�3@&��!?�ݗ���@���^��ٿi�8.W��@��1Y6�3@&��!?�ݗ���@��D5�ٿ�u3��@3��\��3@�����!?ߊ����@�2�/H�ٿ��y�O�@S�(��3@l���!?�p�S޴@�2�/H�ٿ��y�O�@S�(��3@l���!?�p�S޴@�2�/H�ٿ��y�O�@S�(��3@l���!?�p�S޴@fw �ٿ�Υw���@XI�`��3@g8���!?f��Wq�@��I�ٿB�o0!b�@?[��B�3@��$���!?�{3:��@��I�ٿB�o0!b�@?[��B�3@��$���!?�{3:��@��I�ٿB�o0!b�@?[��B�3@��$���!?�{3:��@��I�ٿB�o0!b�@?[��B�3@��$���!?�{3:��@ک�)�ٿ"�/Xf��@����|�3@��{�!?4���a�@ک�)�ٿ"�/Xf��@����|�3@��{�!?4���a�@ک�)�ٿ"�/Xf��@����|�3@��{�!?4���a�@ک�)�ٿ"�/Xf��@����|�3@��{�!?4���a�@��~�ٿ�VG ��@v��	�3@Q�cf�!?6G'p�@��~�ٿ�VG ��@v��	�3@Q�cf�!?6G'p�@��~�ٿ�VG ��@v��	�3@Q�cf�!?6G'p�@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@��dԐٿ�)�C��@���cD�3@�χo�!?쎈��@͝��e�ٿ��m̂��@�O6���3@\� �\�!?���N��@͝��e�ٿ��m̂��@�O6���3@\� �\�!?���N��@͝��e�ٿ��m̂��@�O6���3@\� �\�!?���N��@͝��e�ٿ��m̂��@�O6���3@\� �\�!?���N��@͝��e�ٿ��m̂��@�O6���3@\� �\�!?���N��@�C���ٿ�t,1�7�@�eu��3@�Ð��!?�+㧵�@j֫k�ٿ�X���I�@�k�F�3@_�"췐!?�Jզ��@j֫k�ٿ�X���I�@�k�F�3@_�"췐!?�Jզ��@�rP�ٿ��J^��@o�x~?4@�o�Mv�!?�A����@�rP�ٿ��J^��@o�x~?4@�o�Mv�!?�A����@�rP�ٿ��J^��@o�x~?4@�o�Mv�!?�A����@���1�ٿ���K,��@a����3@j	HA��!?��%�"�@���1�ٿ���K,��@a����3@j	HA��!?��%�"�@8�k��ٿS��	��@��Ļ4@b����!?���RD�@�8��ٿ_a��i�@���W�3@�)�C�!?X3fid�@�8��ٿ_a��i�@���W�3@�)�C�!?X3fid�@�8��ٿ_a��i�@���W�3@�)�C�!?X3fid�@�8��ٿ_a��i�@���W�3@�)�C�!?X3fid�@�L����ٿo�4��@ ���3@�˻`�!?�|���@�L����ٿo�4��@ ���3@�˻`�!?�|���@�L����ٿo�4��@ ���3@�˻`�!?�|���@�L����ٿo�4��@ ���3@�˻`�!?�|���@�L����ٿo�4��@ ���3@�˻`�!?�|���@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@�/�ٿf�#�9��@fQ���3@ܡ�!?*�s�nR�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@��N��ٿP�x��$�@�4�$q�3@��Ώ!?�0�o�@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@

�'�ٿ#���s�@�l�J��3@R!Qm�!?�l����@��R�=�ٿ�W���@}�'i��3@Wc~�!?�lң�=�@��R�=�ٿ�W���@}�'i��3@Wc~�!?�lң�=�@��R�=�ٿ�W���@}�'i��3@Wc~�!?�lң�=�@��R�=�ٿ�W���@}�'i��3@Wc~�!?�lң�=�@�<Cz��ٿ�R-+_>�@���V�3@x��k�!?,?"	�յ@�^}��ٿ��2V���@zJҙ��3@�x�|�!?I���8�@��
�ٿ4�{�=�@Tw.��3@�M�!?���H��@��
�ٿ4�{�=�@Tw.��3@�M�!?���H��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@�IbZ1�ٿ'J��\��@N?M �3@�4��A�!?V|Ee��@^�n��ٿ-Pu	���@������3@��o^%�!?�HP/��@�
�ٿ��!��G�@��ҿ��3@MU�7�!?E?X�FR�@����X�ٿO8�R�@9�F�#�3@�
gS�!?q�Mቴ@����X�ٿO8�R�@9�F�#�3@�
gS�!?q�Mቴ@����X�ٿO8�R�@9�F�#�3@�
gS�!?q�Mቴ@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�u���ٿD=�.���@_���l�3@t6[��!?-��m���@�o��9�ٿ��|�V�@�v^G
�3@�6��!?�*i��!�@�o��9�ٿ��|�V�@�v^G
�3@�6��!?�*i��!�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@Y��t��ٿP���q\�@�^�-�3@��L�!?K�$�@x�/?�ٿ?Q+�`i�@�M�D�3@َ�ip�!?��}}Tb�@���p�ٿk[6��A�@�G�@�3@%=ُN�!?�N�=�3�@���p�ٿk[6��A�@�G�@�3@%=ُN�!?�N�=�3�@���p�ٿk[6��A�@�G�@�3@%=ُN�!?�N�=�3�@���p�ٿk[6��A�@�G�@�3@%=ُN�!?�N�=�3�@���p�ٿk[6��A�@�G�@�3@%=ُN�!?�N�=�3�@��K��ٿ�:�����@G<��3@.�w_�!?@����@��K��ٿ�:�����@G<��3@.�w_�!?@����@r�@˙ٿu�[����@m�g���3@l ����!?�.�O���@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@4��(�ٿT����@ҩ��3@�
�8y�!?�Z�o@Y�@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@ȷ�+H�ٿ���N��@�)�J��3@:�j��!?���;´@��G��ٿ-W�-��@�>
���3@]�
Q�!?AI��R�@��G��ٿ-W�-��@�>
���3@]�
Q�!?AI��R�@��G��ٿ-W�-��@�>
���3@]�
Q�!?AI��R�@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@�cA��ٿ�:��3��@��ZM��3@��P�!?v *A��@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@rD�uI�ٿ���f �@L�I��3@I�����!?*t�}4(�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@��B)b�ٿH�Q���@U�h�3@\*�O'�!?���.^�@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@G��ٿ�z���:�@h���3@��;�w�!?�JK�ȵ@L
,�&�ٿ����.��@B!+�[4@>�Ar�!?�*�G��@�9S�ٿ�1Z=uJ�@b��3@I��f��!?�Ӏ�>/�@�9S�ٿ�1Z=uJ�@b��3@I��f��!?�Ӏ�>/�@�!��B�ٿ������@2����3@�ےd�!?���W�I�@�!��B�ٿ������@2����3@�ےd�!?���W�I�@�!��B�ٿ������@2����3@�ےd�!?���W�I�@�!��B�ٿ������@2����3@�ےd�!?���W�I�@�!��B�ٿ������@2����3@�ےd�!?���W�I�@,��K[�ٿ����<�@���i��3@�z��m�!?�τ�v��@,��K[�ٿ����<�@���i��3@�z��m�!?�τ�v��@,��K[�ٿ����<�@���i��3@�z��m�!?�τ�v��@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@1��?�ٿ��$"��@H�#6�3@�0eu��!?��_�@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@��8��ٿ���ĉ@�@L����3@e�(���!?!�'�=µ@�Ty��ٿv8�Ϡj�@D�1ĭ�3@�
;b�!?�Y"��@�Ty��ٿv8�Ϡj�@D�1ĭ�3@�
;b�!?�Y"��@�Ty��ٿv8�Ϡj�@D�1ĭ�3@�
;b�!?�Y"��@�Ty��ٿv8�Ϡj�@D�1ĭ�3@�
;b�!?�Y"��@�Ty��ٿv8�Ϡj�@D�1ĭ�3@�
;b�!?�Y"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@^ϑ��ٿ�]�$��@g��
~�3@��r���!?q7�"��@6�Wa��ٿZ���?�@�ϜQ��3@�'QY�!?l�?���@6�Wa��ٿZ���?�@�ϜQ��3@�'QY�!?l�?���@6�Wa��ٿZ���?�@�ϜQ��3@�'QY�!?l�?���@6�Wa��ٿZ���?�@�ϜQ��3@�'QY�!?l�?���@6�Wa��ٿZ���?�@�ϜQ��3@�'QY�!?l�?���@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@\w(]�ٿ��;+��@G(�[�3@�"�I�!?p�����@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�����ٿ_��g�@���E�3@�\p�!?�7��"_�@�},#��ٿ�%7����@�a�R��3@�����!?�-n#G�@֠����ٿ�,�����@��p
��3@b�܏�!?/�5�?�@֠����ٿ�,�����@��p
��3@b�܏�!?/�5�?�@֠����ٿ�,�����@��p
��3@b�܏�!?/�5�?�@֠����ٿ�,�����@��p
��3@b�܏�!?/�5�?�@֠����ٿ�,�����@��p
��3@b�܏�!?/�5�?�@yY���ٿ��*����@�=@���3@s��{�!?o��t!�@yY���ٿ��*����@�=@���3@s��{�!?o��t!�@yY���ٿ��*����@�=@���3@s��{�!?o��t!�@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@���m�ٿ:}�"���@ �=.��3@K����!?.v2���@e�&漑ٿ��Kf�@:s��3@�_A��!?y�$�tp�@0�BҔٿC���%�@��gn�3@7}�d�!?Y �X�@���ٿ�JH&�@�uE��3@����~�!?�'�
�@�y+Ё�ٿ��&�ҟ�@x�m��3@��r��!?l�
��@�y+Ё�ٿ��&�ҟ�@x�m��3@��r��!?l�
��@�y+Ё�ٿ��&�ҟ�@x�m��3@��r��!?l�
��@ȕ�ٿm=w&��@�\�eZ�3@D��l�!?�ݺZ�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@�}SY�ٿ|֧�5��@��d�3@��Ư�!?�̿�޲�@"H-�)�ٿ�#))��@1�(��3@��E���!?������@"H-�)�ٿ�#))��@1�(��3@��E���!?������@����ٿ�U�ނ/�@.�C4@�6�F�!?���D��@����ٿ�U�ނ/�@.�C4@�6�F�!?���D��@����ٿ�U�ނ/�@.�C4@�6�F�!?���D��@����ٿ�U�ނ/�@.�C4@�6�F�!?���D��@����ٿ�U�ނ/�@.�C4@�6�F�!?���D��@�����ٿy�����@t$� 4@�J�6׏!?���5M�@�����ٿy�����@t$� 4@�J�6׏!?���5M�@�����ٿy�����@t$� 4@�J�6׏!?���5M�@�-�c��ٿr/�C �@���3@��J&�!?�`\��@�-�c��ٿr/�C �@���3@��J&�!?�`\��@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@N��[�ٿ�0#̄q�@?ʒ���3@r��+�!?��.���@LE�߇�ٿ�	��s��@����3@�ˡ8�!?�Ff�x�@LE�߇�ٿ�	��s��@����3@�ˡ8�!?�Ff�x�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@c;�>^�ٿ�G�U���@�dr�3�3@+�E��!?�BC%
r�@艌h�ٿL���@=��d�3@�֨G�!??�3 `g�@艌h�ٿL���@=��d�3@�֨G�!??�3 `g�@�O�=�ٿ�X��݆�@j�7�4@o
��Z�!?���Gv�@�����ٿ�A�w2��@�ͤ��3@�H�'�!?E-c�b�@�����ٿ�A�w2��@�ͤ��3@�H�'�!?E-c�b�@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@�Aۋ�ٿg���	�@1�:��3@���?4�!?��Z�4��@S����ٿ�}m2��@���4@����!?���ޟ�@S����ٿ�}m2��@���4@����!?���ޟ�@S����ٿ�}m2��@���4@����!?���ޟ�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@��囒ٿ�~G�v#�@�@-+��3@c� V�!?�t|=L�@�/Z�ٿ�������@eN�)$4@�a�#�!?��&ȱR�@�/Z�ٿ�������@eN�)$4@�a�#�!?��&ȱR�@�/Z�ٿ�������@eN�)$4@�a�#�!?��&ȱR�@ˈ�^��ٿҏf)�h�@E�A��	4@����!?����}õ@ˈ�^��ٿҏf)�h�@E�A��	4@����!?����}õ@ �+S�ٿ;��f��@��פ4@WQ4�!?����55�@ �+S�ٿ;��f��@��פ4@WQ4�!?����55�@ �+S�ٿ;��f��@��פ4@WQ4�!?����55�@��/�d�ٿ�.D��@l���3@�\���!?�,��r^�@��/�d�ٿ�.D��@l���3@�\���!?�,��r^�@��/�d�ٿ�.D��@l���3@�\���!?�,��r^�@��/�d�ٿ�.D��@l���3@�\���!?�,��r^�@���1�ٿ��/T]�@�T~��4@̲��!?�����@T�j���ٿ=T���@֝J4@�����!?�rE�o�@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@6T�Ԯ�ٿDf;^2��@�+Z�?4@)^��S�!?���=���@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@FJ�r��ٿH7���p�@�Bt@��3@�=�&��!?�_}Udi�@
��O��ٿt�/p'L�@��p2_�3@� B?�!?Ѐ�2L�@&h�f�ٿ���Ӄ�@�v���3@�U�LX�!?�=\3"�@&h�f�ٿ���Ӄ�@�v���3@�U�LX�!?�=\3"�@&h�f�ٿ���Ӄ�@�v���3@�U�LX�!?�=\3"�@&h�f�ٿ���Ӄ�@�v���3@�U�LX�!?�=\3"�@&h�f�ٿ���Ӄ�@�v���3@�U�LX�!?�=\3"�@�+pu��ٿ������@hZ��}�3@��g��!?AF��~�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@fF�Ee�ٿ�ӭ����@�L'��3@����-�!?~�|1Ǔ�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@u=�>�ٿ���pZ��@���!��3@�d��B�!?kT��K�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@���~�ٿV�/���@NM>5�3@����L�!?ܚ�7�@2�ٿ��4Ka�@(\�A��3@��:��!?��h��@2�ٿ��4Ka�@(\�A��3@��:��!?��h��@D^����ٿ���"���@u�&L�3@��oM��!?^��MӴ@D^����ٿ���"���@u�&L�3@��oM��!?^��MӴ@D^����ٿ���"���@u�&L�3@��oM��!?^��MӴ@D^����ٿ���"���@u�&L�3@��oM��!?^��MӴ@}2��N�ٿ��~�L��@En���3@8h[�]�!?�b~Y�ǵ@�a���ٿ8<H;���@&�q�t�3@+A{�=�!?ۿ_JBT�@OZX��ٿ̮�xv�@�'���3@�VW�!?9oU=8S�@�>��H�ٿ�%F���@��?��4@Kv��u�!?�^_nZ�@�>��H�ٿ�%F���@��?��4@Kv��u�!?�^_nZ�@�>��H�ٿ�%F���@��?��4@Kv��u�!?�^_nZ�@�4)�ٿ�VO���@fS�g�3@���\�!?Zs���/�@�4)�ٿ�VO���@fS�g�3@���\�!?Zs���/�@�4)�ٿ�VO���@fS�g�3@���\�!?Zs���/�@kUQ���ٿ�A�z�/�@�o;��3@C�=�y�!?1W;�s�@kUQ���ٿ�A�z�/�@�o;��3@C�=�y�!?1W;�s�@kUQ���ٿ�A�z�/�@�o;��3@C�=�y�!?1W;�s�@kUQ���ٿ�A�z�/�@�o;��3@C�=�y�!?1W;�s�@kUQ���ٿ�A�z�/�@�o;��3@C�=�y�!?1W;�s�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@=k�V�ٿy#����@QY���3@�s�S�!?�z�LW�@
�8��ٿ���{fC�@vn\�3@Y���!?i�B�P�@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@D4Y3��ٿ�&}Xr�@`wou��3@S|��:�!? �N;��@�n��ٿ\�H̢�@D�/���3@&�i�!?1��S�t�@�n��ٿ\�H̢�@D�/���3@&�i�!?1��S�t�@�n��ٿ\�H̢�@D�/���3@&�i�!?1��S�t�@�n��ٿ\�H̢�@D�/���3@&�i�!?1��S�t�@�!���ٿ�#�	��@J�l�3@ou����!??!h�V�@�!���ٿ�#�	��@J�l�3@ou����!??!h�V�@��ﶒٿn<j[�@e��i�3@�sqK�!?� ����@��ﶒٿn<j[�@e��i�3@�sqK�!?� ����@��ﶒٿn<j[�@e��i�3@�sqK�!?� ����@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@�z%�ٿ�U�׬��@n@�K�3@;���v�!?�>h࿋�@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@[��ٿ�ս���@WB��3@��v`�!?O��+��@� �y�ٿ�:�̘u�@H����3@m���|�!?:f����@|EΪԓٿ��ِ��@I�ܫ��3@�P��ؐ!?��s��@W���ٿխ�FD��@��xG��3@Z�c!?�)��z)�@W���ٿխ�FD��@��xG��3@Z�c!?�)��z)�@W���ٿխ�FD��@��xG��3@Z�c!?�)��z)�@W���ٿխ�FD��@��xG��3@Z�c!?�)��z)�@:�I�ٿ:���^�@gmԴ	�3@�+�!e�!?�頷ȵ@:�I�ٿ:���^�@gmԴ	�3@�+�!e�!?�頷ȵ@dC���ٿ��5��G�@��TZc�3@ ��f�!?��0f�@dC���ٿ��5��G�@��TZc�3@ ��f�!?��0f�@dC���ٿ��5��G�@��TZc�3@ ��f�!?��0f�@dC���ٿ��5��G�@��TZc�3@ ��f�!?��0f�@̎� ĝٿ�$�#��@�$[F��3@'V6�!?�<�=�@̎� ĝٿ�$�#��@�$[F��3@'V6�!?�<�=�@̎� ĝٿ�$�#��@�$[F��3@'V6�!?�<�=�@��tQ�ٿ%��~!�@\�Q�)�3@��� o�!?�!p�馵@��tQ�ٿ%��~!�@\�Q�)�3@��� o�!?�!p�馵@��tQ�ٿ%��~!�@\�Q�)�3@��� o�!?�!p�馵@��tQ�ٿ%��~!�@\�Q�)�3@��� o�!?�!p�馵@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@y��	��ٿQ��u��@��)�3@��ȵ��!?����l�@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@ǻ�?�ٿ��+S_��@��4��3@�(��w�!?�c�?��@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@�9���ٿh��ߧ�@G�ve�3@͖b��!?�\��}�@7P|\�ٿ�9��z�@�YU�y�3@s&3�!?�6e�i�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@��0 �ٿSBK|�E�@e_���3@��z��!?��paғ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@oN���ٿ>E2��@�u?G�3@�*�'@�!?́UƬ�@x&Џ��ٿ�bjz��@��
3��3@�|S���!?��ݽ��@x&Џ��ٿ�bjz��@��
3��3@�|S���!?��ݽ��@x&Џ��ٿ�bjz��@��
3��3@�|S���!?��ݽ��@x&Џ��ٿ�bjz��@��
3��3@�|S���!?��ݽ��@x&Џ��ٿ�bjz��@��
3��3@�|S���!?��ݽ��@@?8��ٿI�6$ո�@��J��3@N�i2R�!?�Q���N�@	]�K�ٿOeZ�Y��@�M@���3@r�b��!?.�T�Fʹ@	]�K�ٿOeZ�Y��@�M@���3@r�b��!?.�T�Fʹ@����Ǔٿ��1�Q�@}N>��3@�Hʚ�!?��q�|�@���g �ٿd%x3��@�,vtt�3@���t�!?9�%wɴ�@���g �ٿd%x3��@�,vtt�3@���t�!?9�%wɴ�@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@-
3կ�ٿ��!o��@���Ӆ�3@�)�_�!?fL%eI̴@�����ٿ2�^�P��@>����3@	��h��!?�A�0y�@�����ٿ2�^�P��@>����3@	��h��!?�A�0y�@�����ٿ2�^�P��@>����3@	��h��!?�A�0y�@�����ٿ2�^�P��@>����3@	��h��!?�A�0y�@�����ٿ2�^�P��@>����3@	��h��!?�A�0y�@ ��K��ٿ��$���@Բ��b�3@�^����!?�G�r1=�@]���ٿ�eѓD�@�c0�E�3@ug����!?�����@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@^)�9ÔٿtWm߾��@`��6�3@~E�!m�!?��k��@lzml�ٿ�L�s�<�@���Cg�3@3��<��!?I���W�@lzml�ٿ�L�s�<�@���Cg�3@3��<��!?I���W�@��W'�ٿ�y�2u�@8?˝R�3@t�ڗ��!?1��0�@��W'�ٿ�y�2u�@8?˝R�3@t�ڗ��!?1��0�@��W'�ٿ�y�2u�@8?˝R�3@t�ڗ��!?1��0�@��W'�ٿ�y�2u�@8?˝R�3@t�ڗ��!?1��0�@��W'�ٿ�y�2u�@8?˝R�3@t�ڗ��!?1��0�@��N<ݗٿ�V= s�@�N��4@8=��!?��0���@��N<ݗٿ�V= s�@�N��4@8=��!?��0���@��N<ݗٿ�V= s�@�N��4@8=��!?��0���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��if4�ٿ	����@��y�3@��y��!?}���@��['i�ٿ���~�N�@XUtj�3@�Y�6��!?L�9|��@��['i�ٿ���~�N�@XUtj�3@�Y�6��!?L�9|��@��['i�ٿ���~�N�@XUtj�3@�Y�6��!?L�9|��@��['i�ٿ���~�N�@XUtj�3@�Y�6��!?L�9|��@÷��ܐٿSҬmqX�@_	d.F 4@�4攕�!?Gw�ʵ��@÷��ܐٿSҬmqX�@_	d.F 4@�4攕�!?Gw�ʵ��@÷��ܐٿSҬmqX�@_	d.F 4@�4攕�!?Gw�ʵ��@÷��ܐٿSҬmqX�@_	d.F 4@�4攕�!?Gw�ʵ��@÷��ܐٿSҬmqX�@_	d.F 4@�4攕�!?Gw�ʵ��@U�v6��ٿ!��U,�@n�R1��3@�wO�Ɛ!?��6NY��@U�v6��ٿ!��U,�@n�R1��3@�wO�Ɛ!?��6NY��@��[��ٿL_��!��@f�i���3@�y�Mw�!?1���z$�@��H�͕ٿ���(�@f,dt)�3@�!d{�!?qD�$�@��H�͕ٿ���(�@f,dt)�3@�!d{�!?qD�$�@��8l�ٿ��ۛ%�@�jՖ��3@�쯈O�!?�#g�>�@��8l�ٿ��ۛ%�@�jՖ��3@�쯈O�!?�#g�>�@��8l�ٿ��ۛ%�@�jՖ��3@�쯈O�!?�#g�>�@��9���ٿ��N�e�@���4@��&�)�!?�;��H�@�k�^k�ٿ�E=���@*|�a� 4@��T��!?�\0J{��@�k�^k�ٿ�E=���@*|�a� 4@��T��!?�\0J{��@�k�^k�ٿ�E=���@*|�a� 4@��T��!?�\0J{��@��e�ٿ��
י��@��ZF��3@�� �!?�h���@��e�ٿ��
י��@��ZF��3@�� �!?�h���@Ďɨ#�ٿ�.��[�@���_�3@�)���!?����ô@Ďɨ#�ٿ�.��[�@���_�3@�)���!?����ô@ނ8��ٿ(�SbI�@/��{=�3@a��!?E����@ނ8��ٿ(�SbI�@/��{=�3@a��!?E����@ނ8��ٿ(�SbI�@/��{=�3@a��!?E����@ނ8��ٿ(�SbI�@/��{=�3@a��!?E����@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@��?ƚٿ��F�M��@�w,Ϲ�3@mZ���!?��n���@i�X9�ٿgї���@*"� A�3@z�B�܏!?.�zG<�@i�X9�ٿgї���@*"� A�3@z�B�܏!?.�zG<�@i�X9�ٿgї���@*"� A�3@z�B�܏!?.�zG<�@�X����ٿ�L���@�����3@��'�!?�+fk �@�X����ٿ�L���@�����3@��'�!?�+fk �@�X����ٿ�L���@�����3@��'�!?�+fk �@�X����ٿ�L���@�����3@��'�!?�+fk �@�X����ٿ�L���@�����3@��'�!?�+fk �@�X����ٿ�L���@�����3@��'�!?�+fk �@����ٿ��QXH�@Z�!���3@Ɔ�d��!?c��9���@����ٿ��QXH�@Z�!���3@Ɔ�d��!?c��9���@����ٿ��QXH�@Z�!���3@Ɔ�d��!?c��9���@�����ٿ��|(5u�@l�%�,4@��l�Ő!?�W�M���@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@��J�ٿ�G�I3��@���q�3@��Ս��!?ȉ,�>�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@�>��:�ٿ��,�$��@XQ�W��3@���R�!?y��x�@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@��!z �ٿ?v0���@�X���3@I�a;�!?E�#wH��@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@G�{#��ٿ�Vg"#�@}�j��3@��b� �!?�G���@V�.�ٿ�}��?K�@�@��4@�[�AZ�!?�h_]��@V�.�ٿ�}��?K�@�@��4@�[�AZ�!?�h_]��@V�.�ٿ�}��?K�@�@��4@�[�AZ�!?�h_]��@H����ٿ֌K��@��k��3@шej�!?E�0��i�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@ͬ^�X�ٿԡH��@���h��3@�ǻ[n�!?E9g�
�@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@y��y�ٿ�g����@o3�jF�3@��
��!?�z��@�M�j�ٿ����@h�c_7 4@,��m|�!?+��'G�@�M�j�ٿ����@h�c_7 4@,��m|�!?+��'G�@�M�j�ٿ����@h�c_7 4@,��m|�!?+��'G�@�M�j�ٿ����@h�c_7 4@,��m|�!?+��'G�@$��ٿ����@���W}�3@kjE�1�!?)�\�F�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@�����ٿI���|�@�ǀ?k�3@�b���!?��z�a�@wB��l�ٿpMV�=��@94��4@�6�e��!?U�[��@wB��l�ٿpMV�=��@94��4@�6�e��!?U�[��@wB��l�ٿpMV�=��@94��4@�6�e��!?U�[��@��A��ٿ�R_���@�M�`@�3@0#��!?�f���@��A��ٿ�R_���@�M�`@�3@0#��!?�f���@��A��ٿ�R_���@�M�`@�3@0#��!?�f���@�x�/��ٿ�]�L�?�@�/���3@K����!?R"�%p��@�x�/��ٿ�]�L�?�@�/���3@K����!?R"�%p��@)�r��ٿ�ck/w�@ ��1��3@����u�!?��fD��@)�r��ٿ�ck/w�@ ��1��3@����u�!?��fD��@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@����ٿ���1��@�'Qa�3@)V�Q~�!? ��e�@� �ٿ`�b����@�P�3@��`�!?�t�>^ص@� �ٿ`�b����@�P�3@��`�!?�t�>^ص@>��゛ٿ�����@D����3@*q �!?�P,�(��@�-�{�ٿ�_5�FH�@[�^-84@oTP���!?������@�-�{�ٿ�_5�FH�@[�^-84@oTP���!?������@�-�{�ٿ�_5�FH�@[�^-84@oTP���!?������@�-�{�ٿ�_5�FH�@[�^-84@oTP���!?������@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@I���ٿ���A�@����3@�1��|�!?=��ju�@;{����ٿ�3���Z�@wcb�3@�ޛ��!?�Py�
?�@;{����ٿ�3���Z�@wcb�3@�ޛ��!?�Py�
?�@�l�z�ٿ+"�v���@��<�B�3@$�K��!?+77O:�@��b�y�ٿ�j�c���@���|��3@RO��!?���1T��@�[љٿ��=d��@x�d��3@�X��}�!?T������@�[љٿ��=d��@x�d��3@�X��}�!?T������@�[љٿ��=d��@x�d��3@�X��}�!?T������@�[љٿ��=d��@x�d��3@�X��}�!?T������@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�| ��ٿ�!f�m�@�95��3@+=N�g�!?��iC䷵@�xo�ٿ�� _Y�@�0ʗQ�3@���Y�!?(��~�*�@�xo�ٿ�� _Y�@�0ʗQ�3@���Y�!?(��~�*�@,B۔ٿn�a2'��@&g���3@��˧Y�!?�N���@;���ٿ@������@.��p��3@f���!?;Cg��ǵ@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@lY;�u�ٿًn"��@���K�3@���Y�!?���?��@��w�ٿLvM�;�@��9���3@�ԡ�i�!?��	5O"�@Q� � �ٿ]ͼ�Y��@|dG6��3@��8<o�!?sIE2�@Q� � �ٿ]ͼ�Y��@|dG6��3@��8<o�!?sIE2�@��1�i�ٿ�R�^L��@6�;�$�3@>���Z�!?�i-x�Ӵ@��1�i�ٿ�R�^L��@6�;�$�3@>���Z�!?�i-x�Ӵ@��1�i�ٿ�R�^L��@6�;�$�3@>���Z�!?�i-x�Ӵ@�,9V �ٿ9���')�@��J�3@�UM\�!?�̇@Z�@�,9V �ٿ9���')�@��J�3@�UM\�!?�̇@Z�@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@E��u�ٿ����@w��~�3@�'�0�!?�~=����@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@�Kk�ٿj�^����@BMAI�3@�)�Jt�!?��
�_�@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���>�ٿ�(�W��@'V�sJ�3@��ڹD�!?���I���@���Ƒٿ�wuf��@���3@���r�!?���$��@���Ƒٿ�wuf��@���3@���r�!?���$��@���Ƒٿ�wuf��@���3@���r�!?���$��@���Ƒٿ�wuf��@���3@���r�!?���$��@���Ƒٿ�wuf��@���3@���r�!?���$��@���Ƒٿ�wuf��@���3@���r�!?���$��@�A���ٿ7�S��@IK
6��3@O��I�!?J)�\��@�A���ٿ7�S��@IK
6��3@O��I�!?J)�\��@�A���ٿ7�S��@IK
6��3@O��I�!?J)�\��@�A���ٿ7�S��@IK
6��3@O��I�!?J)�\��@�}���ٿ��OT��@�9ikr�3@�ۤ �!?�C��vɵ@�}���ٿ��OT��@�9ikr�3@�ۤ �!?�C��vɵ@�}���ٿ��OT��@�9ikr�3@�ۤ �!?�C��vɵ@�����ٿ�L��l�@(%�X�3@([芐!?�N~�@�����ٿ�L��l�@(%�X�3@([芐!?�N~�@�����ٿ�L��l�@(%�X�3@([芐!?�N~�@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@3i�V�ٿ$�V��@OE���3@����F�!?>x���̴@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@"�@-��ٿ���KW��@d�����3@�2_*�!?L��ƴ@�ғv̓ٿP��2A2�@;�ei��3@|�5��!?PQGn���@�ғv̓ٿP��2A2�@;�ei��3@|�5��!?PQGn���@�6�ٿ!_���L�@ҁ$4�3@e4��!?t�%ٍ��@��A@ۓٿs�G�\�@[+ekB�3@*��f�!?C	�[�`�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@D��ґٿy,���}�@7�ݵ~�3@V�}P�!?�g�@�͒ٿQp��k�@�����3@�#�!?�_s��o�@�͒ٿQp��k�@�����3@�#�!?�_s��o�@4Kᩉ�ٿ�n:�@)C��s�3@�?�v��!?������@4Kᩉ�ٿ�n:�@)C��s�3@�?�v��!?������@4Kᩉ�ٿ�n:�@)C��s�3@�?�v��!?������@�@��%�ٿ�~�����@E���P�3@(���5�!?g��M�@�@��%�ٿ�~�����@E���P�3@(���5�!?g��M�@�@��%�ٿ�~�����@E���P�3@(���5�!?g��M�@�5�]�ٿ :��G�@r�7���3@ nAi,�!?�g�WzA�@��WD�ٿ�T ��@sU^
��3@1na�!?� �Ѵ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@ӡ��ٿ�Wͩj�@�m�4>�3@������!?�2�'�ٴ@Yy?�ٿ�l�{J�@�ɦ��4@�Z�֐!?U����l�@Yy?�ٿ�l�{J�@�ɦ��4@�Z�֐!?U����l�@Yy?�ٿ�l�{J�@�ɦ��4@�Z�֐!?U����l�@Yy?�ٿ�l�{J�@�ɦ��4@�Z�֐!?U����l�@Yy?�ٿ�l�{J�@�ɦ��4@�Z�֐!?U����l�@�_bsW�ٿvЮkҼ�@JP^|	4@��Nj��!?��m�@&��;�ٿ���w�W�@	�Ehf�3@�	|�W�!?h�"[
ܴ@�wSs��ٿ�"�gp7�@[FS!E4@̮�M��!?"���d��@0�;a�ٿ��Uq$7�@��;�3@���f��!?b�B��x�@0�;a�ٿ��Uq$7�@��;�3@���f��!?b�B��x�@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@�o�Ƙٿ1�+aP�@�B8@L�3@���E��!?		����@m��C8�ٿ\�����@uo	��3@9��n�!?�l�r��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@ś{IZ�ٿ��z(���@eViP��3@PM�\L�!?3�To��@�AZϚٿڋۍ���@��:��3@L?�ee�!?��R����@�p����ٿ������@�)���3@�{�6�!?G���+F�@�p����ٿ������@�)���3@�{�6�!?G���+F�@�p����ٿ������@�)���3@�{�6�!?G���+F�@�p����ٿ������@�)���3@�{�6�!?G���+F�@�/�P�ٿ�ӽ�l��@��N?S�3@,���^�!?.���@KIr�ǘٿ��Z
A��@GpR"^�3@���O�!?Dw��@KIr�ǘٿ��Z
A��@GpR"^�3@���O�!?Dw��@KIr�ǘٿ��Z
A��@GpR"^�3@���O�!?Dw��@KIr�ǘٿ��Z
A��@GpR"^�3@���O�!?Dw��@�E8?�ٿ������@k&��3@K�c��!?3�����@�E8?�ٿ������@k&��3@K�c��!?3�����@�E8?�ٿ������@k&��3@K�c��!?3�����@�E8?�ٿ������@k&��3@K�c��!?3�����@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@h񋄇�ٿ��B�^�@/Iޑ�3@B�����!?Su���@�^��ٿ
.kz��@�N����3@��5��!?ma���@�^��ٿ
.kz��@�N����3@��5��!?ma���@�^��ٿ
.kz��@�N����3@��5��!?ma���@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�t��j�ٿ��Ǎ)��@�� 4��3@8��jz�!?�HX8��@�N��n�ٿNz��@ۯ�k��3@�i���!?�U���@#�y��ٿL�ͣ��@���3@Gi1��!?hw�6-H�@&����ٿQ�(����@Q�-F�3@��QDP�!?pL�0�@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@�R&1�ٿl#����@5��
��3@�����!?�bU�ô@|T���ٿ��"��g�@3ׁ�% 4@��q��!?��a�~�@|T���ٿ��"��g�@3ׁ�% 4@��q��!?��a�~�@�qՒ��ٿP���@��d��3@V�dS�!?��^��S�@�qՒ��ٿP���@��d��3@V�dS�!?��^��S�@>���a�ٿ�!�|&�@b�J�#�3@U{�G�!?X��b��@>���a�ٿ�!�|&�@b�J�#�3@U{�G�!?X��b��@>���a�ٿ�!�|&�@b�J�#�3@U{�G�!?X��b��@>���a�ٿ�!�|&�@b�J�#�3@U{�G�!?X��b��@>���a�ٿ�!�|&�@b�J�#�3@U{�G�!?X��b��@�#y�ٿ(��8ڣ�@o�	�3@�	q��!?�>3�U��@�#y�ٿ(��8ڣ�@o�	�3@�	q��!?�>3�U��@�#y�ٿ(��8ڣ�@o�	�3@�	q��!?�>3�U��@�#y�ٿ(��8ڣ�@o�	�3@�	q��!?�>3�U��@�#y�ٿ(��8ڣ�@o�	�3@�	q��!?�>3�U��@AG��=�ٿL�·V�@򋒯W�3@��eW�!?�C&�@AG��=�ٿL�·V�@򋒯W�3@��eW�!?�C&�@u�Ӝz�ٿ�(�44�@Ո�T*�3@[���B�!?��7�0F�@u�Ӝz�ٿ�(�44�@Ո�T*�3@[���B�!?��7�0F�@7&�A��ٿi��sr�@�^0�'�3@
��I+�!?�bՋ��@7&�A��ٿi��sr�@�^0�'�3@
��I+�!?�bՋ��@7&�A��ٿi��sr�@�^0�'�3@
��I+�!?�bՋ��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@HZΨؔٿy�3$�N�@o�i[�3@�8���!?�+S��@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@ٍ���ٿ-��擱�@U���3@G6N/�!?�T4�]q�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@|��`��ٿ5I]Y_w�@�wr��3@���=�!?G��8�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@���<5�ٿ����5�@�)�s��3@m��{w�!?0?,�m�@�@��ٿd���� �@HZ���3@u�ȗ�!?E�)��@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@��R��ٿ��E�߅�@���|{�3@QN�v�!?���讴@x��ٿ��^(���@[�V��3@��~��!?q�f���@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@�3��C�ٿ�H���@��RR��3@���f�!?6G�b�@vΒ�Øٿ~Ż�@S�1"�3@��U���!?����Ӵ@7�g���ٿ�WX�/t�@u�r�3@.яً�!?l�}:5�@7�g���ٿ�WX�/t�@u�r�3@.яً�!?l�}:5�@{�5���ٿ�ʪ��K�@�?� �3@�E�3�!?B�$�r{�@{�5���ٿ�ʪ��K�@�?� �3@�E�3�!?B�$�r{�@{�5���ٿ�ʪ��K�@�?� �3@�E�3�!?B�$�r{�@{�5���ٿ�ʪ��K�@�?� �3@�E�3�!?B�$�r{�@� C:�ٿ���,�@�����3@Oi�6d�!?�{O����@� C:�ٿ���,�@�����3@Oi�6d�!?�{O����@� C:�ٿ���,�@�����3@Oi�6d�!?�{O����@� C:�ٿ���,�@�����3@Oi�6d�!?�{O����@mOI(�ٿ���>U�@)Cv�F�3@���8W�!?s���.4�@�8k�S�ٿ~%��7�@�B�#��3@�h�/H�!?�H*�q�@�8k�S�ٿ~%��7�@�B�#��3@�h�/H�!?�H*�q�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@S����ٿL��y�j�@�{&�{�3@������!?' 3襰�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@��am�ٿ4ko��@�>r��3@����f�!?�Z*��-�@�n�%�ٿ���a�@��Dg�3@P�H"8�!??�x��@�n�%�ٿ���a�@��Dg�3@P�H"8�!??�x��@�n�%�ٿ���a�@��Dg�3@P�H"8�!??�x��@��<��ٿ$��^��@��Т<�3@��2��!?yX����@��<��ٿ$��^��@��Т<�3@��2��!?yX����@��<��ٿ$��^��@��Т<�3@��2��!?yX����@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@q�x��ٿ	�����@'	���3@�zCr�!?b~�e���@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@���~�ٿHc;��@@Hh�G�3@R~`V��!?����@�@g��+��ٿ�#ś"�@5I��J�3@'�0��!?���9�@g��+��ٿ�#ś"�@5I��J�3@'�0��!?���9�@g��+��ٿ�#ś"�@5I��J�3@'�0��!?���9�@]����ٿq����@��j�3@ʋ"�#�!?|��4�
�@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@�
�XY�ٿ�����@\V|��3@�,��=�!?�u�W�Ҵ@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@p�����ٿ�;�t���@VVe���3@�>�8�!?%ꥩ�@�G.�ٿ-�?C�/�@�C�]�3@^3|�G�!?9���*�@�G.�ٿ-�?C�/�@�C�]�3@^3|�G�!?9���*�@�G.�ٿ-�?C�/�@�C�]�3@^3|�G�!?9���*�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@$F����ٿ?ON^j�@*_B9��3@�at���!?�]��V�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@|�M���ٿ��Gl��@�+�Q��3@>��D�!?F�nBJl�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@Vf�)�ٿ/���>�@�w@�o�3@�)3%&�!?��Fq�@4�L�ٿ��2C�@wdq��3@��(�$�!?�����@4�L�ٿ��2C�@wdq��3@��(�$�!?�����@4�L�ٿ��2C�@wdq��3@��(�$�!?�����@4�L�ٿ��2C�@wdq��3@��(�$�!?�����@4�L�ٿ��2C�@wdq��3@��(�$�!?�����@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@벍œٿU��H�]�@ҍE���3@��--�!?9������@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@5��!��ٿ0�yX�6�@h�U��3@�;���!?�U}�A3�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@(���ٿ�䌍���@���y��3@���Q*�!?��>M�@�j,��ٿV�Ff��@�HC'�3@�aq�P�!?�`K�Xܴ@�j,��ٿV�Ff��@�HC'�3@�aq�P�!?�`K�Xܴ@�j,��ٿV�Ff��@�HC'�3@�aq�P�!?�`K�Xܴ@�p� �ٿ�Rs3gC�@D�J��3@0�i��!?��9h�t�@�p� �ٿ�Rs3gC�@D�J��3@0�i��!?��9h�t�@�p� �ٿ�Rs3gC�@D�J��3@0�i��!?��9h�t�@�p� �ٿ�Rs3gC�@D�J��3@0�i��!?��9h�t�@D,cw�ٿ��GN��@�(��3@���O�!?22�_R(�@����o�ٿ������@t�
�z4@��|���!?�ה�h��@����o�ٿ������@t�
�z4@��|���!?�ה�h��@l��ٿ�������@���4@픵&�!?=�Xu�@�]��ٿ�7t����@e�Y	�
4@�y1~(�!?9�W�h�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@0��ћٿp����@[3Yc�4@���"��!?)?�1Ns�@@�bdD�ٿ�X`oM�@��w�k4@TA��{�!?;i:����@@�bdD�ٿ�X`oM�@��w�k4@TA��{�!?;i:����@�P]lL�ٿn}G{*��@d���1�3@�ya g�!?'_��k�@����ٿ�x4��@���:�3@���(�!?�|X�@����ٿ�x4��@���:�3@���(�!?�|X�@����ٿ�x4��@���:�3@���(�!?�|X�@����ٿ�x4��@���:�3@���(�!?�|X�@����ٿ�x4��@���:�3@���(�!?�|X�@ФIRT�ٿ�.�B6��@�^G��3@Zu��!?=t��w�@ФIRT�ٿ�.�B6��@�^G��3@Zu��!?=t��w�@ФIRT�ٿ�.�B6��@�^G��3@Zu��!?=t��w�@ФIRT�ٿ�.�B6��@�^G��3@Zu��!?=t��w�@ФIRT�ٿ�.�B6��@�^G��3@Zu��!?=t��w�@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@�C�b�ٿ^�z��@+���3@u�[�!?\ȕÖ��@��Ϙp�ٿ��"I{��@� ����3@�ki��!?�/{g�ݴ@��Ϙp�ٿ��"I{��@� ����3@�ki��!?�/{g�ݴ@��Ϙp�ٿ��"I{��@� ����3@�ki��!?�/{g�ݴ@i6%�ٿ۹���v�@����3@{�q�!?�.˭�@�@i6%�ٿ۹���v�@����3@{�q�!?�.˭�@�@i6%�ٿ۹���v�@����3@{�q�!?�.˭�@�@i6%�ٿ۹���v�@����3@{�q�!?�.˭�@�@-�����ٿZ��p���@�s:,��3@�Q(��!?[�k$˵@��ؚ;�ٿ{H�����@�F[��3@]D��Ր!?f��	�L�@e�螄�ٿ�V�O}Z�@aB/�z�3@�+
��!?����|�@e�螄�ٿ�V�O}Z�@aB/�z�3@�+
��!?����|�@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@��Ώ��ٿ��(��K�@�;&�G�3@�W�F�!?/�(z��@EţW�ٿ���2Y��@�R��3@����!?�0
�ϟ�@EţW�ٿ���2Y��@�R��3@����!?�0
�ϟ�@EţW�ٿ���2Y��@�R��3@����!?�0
�ϟ�@EţW�ٿ���2Y��@�R��3@����!?�0
�ϟ�@EţW�ٿ���2Y��@�R��3@����!?�0
�ϟ�@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@�͑S�ٿu�:~F��@؃�%�3@�35�&�!?�$$aӴ@��F_őٿr��5�@5k.r6�3@���eU�!?b��\�@��F_őٿr��5�@5k.r6�3@���eU�!?b��\�@�uq�ٿ��t�d��@���b4�3@C� w]�!??+��[�@�uq�ٿ��t�d��@���b4�3@C� w]�!??+��[�@�uq�ٿ��t�d��@���b4�3@C� w]�!??+��[�@�uq�ٿ��t�d��@���b4�3@C� w]�!??+��[�@�uq�ٿ��t�d��@���b4�3@C� w]�!??+��[�@���\l�ٿBu�!3�@�3�W�3@��Y�!?T���5*�@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@(��O�ٿ"2 <�
�@�P9��3@#b}ky�!?c<B(��@�4v��ٿ�d���@K�DE�3@ȋsa^�!?�|��B�@�4v��ٿ�d���@K�DE�3@ȋsa^�!?�|��B�@>9�>��ٿ>%�Q�U�@"X�sh�3@.�l\��!?�e��L�@>9�>��ٿ>%�Q�U�@"X�sh�3@.�l\��!?�e��L�@VW�Ȇ�ٿ�S��)��@���/�3@�� 6�!?�K�*y�@VW�Ȇ�ٿ�S��)��@���/�3@�� 6�!?�K�*y�@VW�Ȇ�ٿ�S��)��@���/�3@�� 6�!?�K�*y�@VW�Ȇ�ٿ�S��)��@���/�3@�� 6�!?�K�*y�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@Ȩ����ٿ@���D�@9��!�3@4�$(Z�!?�yӀd�@�f(�$�ٿ
�����@F�����3@q/JX[�!?-rA��@�f(�$�ٿ
�����@F�����3@q/JX[�!?-rA��@�f(�$�ٿ
�����@F�����3@q/JX[�!?-rA��@L�ѭ�ٿK��O��@S����3@#l7�<�!?��p��@L�ѭ�ٿK��O��@S����3@#l7�<�!?��p��@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@#�pXϖٿC��H���@ش�'�3@>y[EG�!?��;��R�@b[KE��ٿ��ԉ��@O�`��3@���V�!?�lN��G�@b[KE��ٿ��ԉ��@O�`��3@���V�!?�lN��G�@�#���ٿ�k�����@�
x��3@�˕�6�!?O��0õ@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@x�&�G�ٿx���5�@��]'�3@��(3��!?4���@��`��ٿ���`j�@��qgy�3@	#b���!?*�)E�@��`��ٿ���`j�@��qgy�3@	#b���!?*�)E�@��`��ٿ���`j�@��qgy�3@	#b���!?*�)E�@��`��ٿ���`j�@��qgy�3@	#b���!?*�)E�@jċђ�ٿ�{(Y���@�e ��3@�{��p�!?65�����@jċђ�ٿ�{(Y���@�e ��3@�{��p�!?65�����@jċђ�ٿ�{(Y���@�e ��3@�{��p�!?65�����@jċђ�ٿ�{(Y���@�e ��3@�{��p�!?65�����@_n�ٿ[HXe6�@|��X$�3@J㶠��!?�i<D��@_n�ٿ[HXe6�@|��X$�3@J㶠��!?�i<D��@��w�7�ٿ��S���@���/�3@C�uD�!? �@A�״@��w�7�ٿ��S���@���/�3@C�uD�!? �@A�״@��w�7�ٿ��S���@���/�3@C�uD�!? �@A�״@x�,̈�ٿ¿��
=�@�i%�F�3@��^�!?Q����@x�,̈�ٿ¿��
=�@�i%�F�3@��^�!?Q����@x�,̈�ٿ¿��
=�@�i%�F�3@��^�!?Q����@x�,̈�ٿ¿��
=�@�i%�F�3@��^�!?Q����@x�,̈�ٿ¿��
=�@�i%�F�3@��^�!?Q����@�D�E��ٿ!���i]�@F{�N��3@Ư�7�!?�B[a��@�D�E��ٿ!���i]�@F{�N��3@Ư�7�!?�B[a��@���n�ٿ�6E�S'�@	|�_��3@`_��!?|t�R�@̵����ٿ{�yA�e�@H�3�4@��d�!?�,��ύ�@̵����ٿ{�yA�e�@H�3�4@��d�!?�,��ύ�@̵����ٿ{�yA�e�@H�3�4@��d�!?�,��ύ�@̵����ٿ{�yA�e�@H�3�4@��d�!?�,��ύ�@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�:�-��ٿ��P5��@�Qj |4@h.|1�!?�k�P���@�e��<�ٿ=�cw;�@X7�Z4@��x�P�!?
�M0�@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@�8��ٿO�/ԋ�@M�b_�3@=��HP�!?#?~#��@���;�ٿ�]�b���@�`
�3@��F	�!?�+t*�9�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@CM���ٿjs����@���^��3@��W�!?��Q7wx�@Q�}��ٿ�b�	[�@M7�r�4@��]�!?���K�´@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�����ٿy�ZH���@��4Ӕ 4@�6�!?�0�ٛ�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�,�ĘٿX>
�@�@��*?x�3@Ż���!?A�F�N�@�;&�ٿ2���@s|N��3@wj��5�!?Y��2r�@��L!�ٿ�Z
f�@����4@S=�#B�!?���@�K�Q�ٿ+�B���@x�9B'�3@�-��!?�=�@�u�@����ٿ$jGk�@��Mș4@ �|�!?�'�,��@����ٿ$jGk�@��Mș4@ �|�!?�'�,��@����ٿ$jGk�@��Mș4@ �|�!?�'�,��@v��r�ٿ2���@n�4@L70�0�!?	�����@��eq�ٿTQ#��@l��Z 4@1���l�!?�\v:P�@��eq�ٿTQ#��@l��Z 4@1���l�!?�\v:P�@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@̥�!�ٿ��P���@RT��14@=�-��!?���۴@1Sm��ٿ+�x~ea�@�V��3@EZ�<P�!?_��Fwʹ@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@�I��P�ٿ�l3�/�@�Ҩ,J�3@h;�m�!?;%�7Ǟ�@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@��B���ٿΛ�F��@�pZ���3@աo|Z�!?�d�lݴ@
�ߴ�ٿ��)h˛�@1��H�3@ֱ�J�!?�l�ķ(�@
�ߴ�ٿ��)h˛�@1��H�3@ֱ�J�!?�l�ķ(�@����ٿ�:c�.�@�B�4*�3@�,� �!?��p���@����ٿ�:c�.�@�B�4*�3@�,� �!?��p���@����ٿ�:c�.�@�B�4*�3@�,� �!?��p���@��!���ٿ��AYT�@a~�P��3@A+�,n�!?V�"��@��!���ٿ��AYT�@a~�P��3@A+�,n�!?V�"��@��!���ٿ��AYT�@a~�P��3@A+�,n�!?V�"��@��!���ٿ��AYT�@a~�P��3@A+�,n�!?V�"��@��!���ٿ��AYT�@a~�P��3@A+�,n�!?V�"��@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@�-�@јٿ�Wjy��@U��0�3@~�["��!?�uTy�@`fz�ٿ���).9�@���)��3@*���!?�uPg�@`fz�ٿ���).9�@���)��3@*���!?�uPg�@`fz�ٿ���).9�@���)��3@*���!?�uPg�@`fz�ٿ���).9�@���)��3@*���!?�uPg�@�b	��ٿښ��{m�@AY�J��3@�&Q�!?������@�b	��ٿښ��{m�@AY�J��3@�&Q�!?������@�b	��ٿښ��{m�@AY�J��3@�&Q�!?������@�b	��ٿښ��{m�@AY�J��3@�&Q�!?������@/خ@��ٿP��}���@�sȍ�3@� ��?�!?.�g�<��@�(�.��ٿ���Yt�@Q��c�3@U:��$�!?����p�@�(�.��ٿ���Yt�@Q��c�3@U:��$�!?����p�@ܑ~ 0�ٿQ�\��|�@*�ZX�3@�!J�2�!?r�vih��@ܑ~ 0�ٿQ�\��|�@*�ZX�3@�!J�2�!?r�vih��@ܑ~ 0�ٿQ�\��|�@*�ZX�3@�!J�2�!?r�vih��@ܑ~ 0�ٿQ�\��|�@*�ZX�3@�!J�2�!?r�vih��@���Q��ٿ�SD���@*��#A�3@����<�!?]N�i��@���Q��ٿ�SD���@*��#A�3@����<�!?]N�i��@+��vǒٿ\]|#���@Q�9��3@��G1�!?�$NA��@+��vǒٿ\]|#���@Q�9��3@��G1�!?�$NA��@+��vǒٿ\]|#���@Q�9��3@��G1�!?�$NA��@UԸy�ٿ�DEDA�@[g�\\4@ʼ���!?
o�X�@UԸy�ٿ�DEDA�@[g�\\4@ʼ���!?
o�X�@�N~�3�ٿM�^�H��@��2��3@i�.a�!?����%�@�N~�3�ٿM�^�H��@��2��3@i�.a�!?����%�@�N~�3�ٿM�^�H��@��2��3@i�.a�!?����%�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@nv��ٿ�p�,�@iA#O��3@��AMd�!?��`J�@�xAU!�ٿ�3��F��@�Y���4@�/�a�!?d�C�R�@�xAU!�ٿ�3��F��@�Y���4@�/�a�!?d�C�R�@�xAU!�ٿ�3��F��@�Y���4@�/�a�!?d�C�R�@�xAU!�ٿ�3��F��@�Y���4@�/�a�!?d�C�R�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@�+��ٿ��"J�@�R1F��3@�rd�J�!?�*�ΐ�@��΢�ٿ��7�O �@�[0,�3@��g�!?������@��΢�ٿ��7�O �@�[0,�3@��g�!?������@��΢�ٿ��7�O �@�[0,�3@��g�!?������@�_P>Ԛٿ'yo]�@W���3@�sgY�!?a����@�_P>Ԛٿ'yo]�@W���3@�sgY�!?a����@�_P>Ԛٿ'yo]�@W���3@�sgY�!?a����@�j�L�ٿB>R4$�@��Vv�3@�-�8�!?~Q����@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@!�x`��ٿ������@gո���3@P�-?Q�!?�`��Dz�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@��g��ٿ�eC���@�����4@�hIY�!?I�a�R�@�hx�ٿ[�Z�Y�@��-Pg�3@r��o�!?&I����@�hx�ٿ[�Z�Y�@��-Pg�3@r��o�!?&I����@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@g���ٿ��c�J��@�Dگe�3@�A=��!?��t8�@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@����%�ٿ����Du�@�)�ľ4@���G�!?=TO���@`���
�ٿyQ�@�(�@��4@,!��C�!?:J�j|�@`���
�ٿyQ�@�(�@��4@,!��C�!?:J�j|�@`���
�ٿyQ�@�(�@��4@,!��C�!?:J�j|�@`���
�ٿyQ�@�(�@��4@,!��C�!?:J�j|�@�ٿ�m0���@���4@������!?��mb�@�@�ٿ�m0���@���4@������!?��mb�@�@��-�ٿ��$����@$0R��3@y?�zs�!?w� ©�@�G��}�ٿZ�B����@ny��4@+��Ej�!?_��dS�@�G��}�ٿZ�B����@ny��4@+��Ej�!?_��dS�@��8��ٿ��Y���@{�F�3@�fm�!?�~v��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@�l�V�ٿU'�	�>�@�X�/�3@���؁�!?�g&��@F��YΠٿKXK>B0�@(ؗ/c�3@��ZvQ�!?����^�@F��YΠٿKXK>B0�@(ؗ/c�3@��ZvQ�!?����^�@F��YΠٿKXK>B0�@(ؗ/c�3@��ZvQ�!?����^�@F��YΠٿKXK>B0�@(ؗ/c�3@��ZvQ�!?����^�@�36�ٿd.s�0�@�}@��3@�QSz�!?a7�	̴@�D0�ٿ���]SE�@���i�3@SD��F�!?3*��S�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�?d_�ٿ�U2���@��3A1�3@�����!?��Y�D�@�H�/7�ٿ)�|�Q��@�3�l� 4@��y�!?��uU�.�@�H�/7�ٿ)�|�Q��@�3�l� 4@��y�!?��uU�.�@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@�p��A�ٿ�Դ%_�@�4�: 4@��\�9�!?ϴ�M�״@u$��?�ٿ��A�2��@���l�3@���N�!?���@u$��?�ٿ��A�2��@���l�3@���N�!?���@u$��?�ٿ��A�2��@���l�3@���N�!?���@u$��?�ٿ��A�2��@���l�3@���N�!?���@u$��?�ٿ��A�2��@���l�3@���N�!?���@u$��?�ٿ��A�2��@���l�3@���N�!?���@�);�ٿd����@/,N��3@1؉`-�!?�uM����@�);�ٿd����@/,N��3@1؉`-�!?�uM����@B���^�ٿ�;`���@A!��3@���j�!?9�����@���4�ٿ��3����@~��o�3@]�,p!�!?1o�o̴@���4�ٿ��3����@~��o�3@]�,p!�!?1o�o̴@���4�ٿ��3����@~��o�3@]�,p!�!?1o�o̴@���5�ٿvN��j�@�q[���3@��s�!?�7�B���@���5�ٿvN��j�@�q[���3@��s�!?�7�B���@���5�ٿvN��j�@�q[���3@��s�!?�7�B���@���5�ٿvN��j�@�q[���3@��s�!?�7�B���@���5�ٿvN��j�@�q[���3@��s�!?�7�B���@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@u���ٿc�l�@���>�3@76U��!?���`q�@����ٿu�H���@K_�7��3@8���!?Z�
AC1�@B4�9ܘٿ�P83K-�@VූD�3@\�$F��!?v�_�aٴ@B4�9ܘٿ�P83K-�@VූD�3@\�$F��!?v�_�aٴ@B4�9ܘٿ�P83K-�@VූD�3@\�$F��!?v�_�aٴ@B4�9ܘٿ�P83K-�@VූD�3@\�$F��!?v�_�aٴ@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@'v2^�ٿ��B���@�V����3@e�T�)�!?*�V��$�@?���ٿ8T���@�վ��3@����h�!?�@r�Ӵ@g9rT�ٿ{H�|C��@̇�q��3@WÊl@�!?��c5O��@g9rT�ٿ{H�|C��@̇�q��3@WÊl@�!?��c5O��@g9rT�ٿ{H�|C��@̇�q��3@WÊl@�!?��c5O��@g9rT�ٿ{H�|C��@̇�q��3@WÊl@�!?��c5O��@g9rT�ٿ{H�|C��@̇�q��3@WÊl@�!?��c5O��@�rP��ٿ�Ȝ(8��@�s�8�3@u�T�!?~A��a�@�rP��ٿ�Ȝ(8��@�s�8�3@u�T�!?~A��a�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@�f�2��ٿ�י]��@`0㬨�3@�m!j�!?MҀь\�@
���ٿ�n$�qg�@Aә���3@���e�!?�w����@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@�ꔋ��ٿ�܈��@��'�3@R��&�!?R����H�@d
(��ٿ^�b���@HpH��3@�D((ޏ!?}��8��@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@(�����ٿ�O�[�@k=�o�3@#[���!?�a��闵@8!|�ؗٿ�y���@��o4@�w�܏!?"�]�@8!|�ؗٿ�y���@��o4@�w�܏!?"�]�@8!|�ؗٿ�y���@��o4@�w�܏!?"�]�@��l��ٿ�r��#�@��5�3@(��9�!?O���E�@��l��ٿ�r��#�@��5�3@(��9�!?O���E�@���/�ٿd�}�|)�@��OØ�3@p��\��!?F�*.��@���/�ٿd�}�|)�@��OØ�3@p��\��!?F�*.��@���/�ٿd�}�|)�@��OØ�3@p��\��!?F�*.��@���/�ٿd�}�|)�@��OØ�3@p��\��!?F�*.��@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@��J�ϒٿ�To���@>�w���3@��5a��!?�o�ᵵ@���ٿ��7�̓�@̍Ƿ*�3@�M;G�!?H!ݑ�h�@?�=j�ٿ�Z�v�_�@nr���3@�>�5P�!?ҔiV��@?�=j�ٿ�Z�v�_�@nr���3@�>�5P�!?ҔiV��@?�=j�ٿ�Z�v�_�@nr���3@�>�5P�!?ҔiV��@69J��ٿ�Ej#3��@b�a{�3@�7��!?O�d��d�@69J��ٿ�Ej#3��@b�a{�3@�7��!?O�d��d�@;Su�ٿ�2��@�����3@r]���!?5�*(1z�@;Su�ٿ�2��@�����3@r]���!?5�*(1z�@;Su�ٿ�2��@�����3@r]���!?5�*(1z�@;Su�ٿ�2��@�����3@r]���!?5�*(1z�@;Su�ٿ�2��@�����3@r]���!?5�*(1z�@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@y��ࠕٿ��$v�@'� ���3@���^�!?[4o�O޵@#!t�"�ٿg���L�@]\}֮�3@��!�!?F��o��@���z�ٿ�#�h8��@����3@Y �!�!?�<>D`�@���z�ٿ�#�h8��@����3@Y �!�!?�<>D`�@���z�ٿ�#�h8��@����3@Y �!�!?�<>D`�@�`�}2�ٿ�N��*��@�8�?��3@�l\�U�!?o�qd�@�`�}2�ٿ�N��*��@�8�?��3@�l\�U�!?o�qd�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@�>��ٿ�Fq����@�����3@������!?b�s�gC�@n���ٿ�g���@h��\��3@I3$�l�!?�7;D�z�@n���ٿ�g���@h��\��3@I3$�l�!?�7;D�z�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@t�,N�ٿ�'��c��@��U�t�3@��w���!?���6�@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@�r�bT�ٿc�t��@O4L4�3@��ģl�!?�a3��@��l��ٿ�z*���@=�s���3@�x F��!?�X�����@��l��ٿ�z*���@=�s���3@�x F��!?�X�����@��l��ٿ�z*���@=�s���3@�x F��!?�X�����@�����ٿ"xp���@�Ξ�3@w#�$�!?��Gi��@�����ٿ"xp���@�Ξ�3@w#�$�!?��Gi��@�����ٿ"xp���@�Ξ�3@w#�$�!?��Gi��@�����ٿ"xp���@�Ξ�3@w#�$�!?��Gi��@�����ٿ"xp���@�Ξ�3@w#�$�!?��Gi��@�$s��ٿZ���]o�@�n%{��3@�R��b�!?(����@Wh��j�ٿg%{���@ֲ���3@���!?�cP´@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@�r݅4�ٿ����#�@�#��s�3@�V�F_�!?[��
�@��<�ٿ���p���@0!"�3@��IFJ�!?����ߴ@��<�ٿ���p���@0!"�3@��IFJ�!?����ߴ@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@v�c�<�ٿryP"�@c�˿+�3@�,�H��!?1;F��@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��my�ٿaT����@�,m��3@03ʠ�!?4�n�dٴ@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@��e�ٿ����@�S�3@�1V�!?z��*5�@)r"��ٿ�x�6�D�@\��+��3@l^F:ߐ!?�Z�֦�@)r"��ٿ�x�6�D�@\��+��3@l^F:ߐ!?�Z�֦�@��d��ٿ�f��W�@�͜��3@8dڐ!?b���c��@X^�ۓٿ�wtkM�@����3@
��e�!?-u��G�@��j�[�ٿM�>�!�@0�t��4@�@�wא!?7RI�`�@��j�[�ٿM�>�!�@0�t��4@�@�wא!?7RI�`�@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@]XAB,�ٿ�����`�@�j$N�3@C�̤��!?/e��"��@D��ٿ��j���@�0n�3@mXt�!?��h�@D��ٿ��j���@�0n�3@mXt�!?��h�@D��ٿ��j���@�0n�3@mXt�!?��h�@D��ٿ��j���@�0n�3@mXt�!?��h�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@�#��&�ٿ"�O8�@~���3@��j�_�!?�o���<�@����ٿ������@Q�}$M�3@� �r/�!?U*��w��@����ٿ������@Q�}$M�3@� �r/�!?U*��w��@����ٿ������@Q�}$M�3@� �r/�!?U*��w��@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@`v���ٿ���A��@-[c�3@@��5'�!?z��T�{�@&��5�ٿ]��,m�@��9~4@į���!?�"o߀�@AX��@�ٿ.PP�<�@��]��3@V�z|�!?&��MtJ�@AX��@�ٿ.PP�<�@��]��3@V�z|�!?&��MtJ�@�����ٿc��߰�@I�M���3@z��	s�!?��Ǎ ��@�����ٿc��߰�@I�M���3@z��	s�!?��Ǎ ��@Xn��%�ٿ�����G�@�7	���3@�	n�e�!?�'C�)�@J����ٿL�l!.��@���8�3@�`E���!?�+6A)�@J����ٿL�l!.��@���8�3@�`E���!?�+6A)�@J����ٿL�l!.��@���8�3@�`E���!?�+6A)�@J����ٿL�l!.��@���8�3@�`E���!?�+6A)�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@�zO��ٿ��Q�h�@��M+3�3@�]o��!?�	
p�@��\���ٿ�"��؜�@6��4@9��c(�!?���`�:�@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@\�n�b�ٿ/��i>�@�1�]��3@��a���!?̮ȁGɴ@Qto��ٿp�����@
!��*�3@B��D�!?��I!��@Qto��ٿp�����@
!��*�3@B��D�!?��I!��@Qto��ٿp�����@
!��*�3@B��D�!?��I!��@���;�ٿôf6r��@���BS�3@�kiHJ�!?r��OEC�@���;�ٿôf6r��@���BS�3@�kiHJ�!?r��OEC�@�ܷ!6�ٿ�f�E�@�m��o�3@^a�5�!?C��,�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@��e�ٿ���?.��@bl���3@��?�@�!?��<C8�@7Bvd�ٿ�pz �@c�Qk��3@;�l�X�!?���K�@7Bvd�ٿ�pz �@c�Qk��3@;�l�X�!?���K�@7Bvd�ٿ�pz �@c�Qk��3@;�l�X�!?���K�@7Bvd�ٿ�pz �@c�Qk��3@;�l�X�!?���K�@7Bvd�ٿ�pz �@c�Qk��3@;�l�X�!?���K�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@�n�ι�ٿlx߸���@������3@�<F.�!?��0R9�@���P��ٿ�L��B��@-�^1�3@��=�O�!?�
L��x�@���P��ٿ�L��B��@-�^1�3@��=�O�!?�
L��x�@`�|e�ٿӧᠡ\�@��Y�3@�&X��!?��wvc�@�9%��ٿ��7y9��@v×#C�3@�h�m��!?{f��g�@�9%��ٿ��7y9��@v×#C�3@�h�m��!?{f��g�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@�����ٿ�#���@�d�.�3@ZZ>)��!?e�v��N�@Iۏs��ٿ!��@3v+`��3@�ԥ��!?g/Z��@Iۏs��ٿ!��@3v+`��3@�ԥ��!?g/Z��@Iۏs��ٿ!��@3v+`��3@�ԥ��!?g/Z��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@G�hE��ٿڨ2���@���i�3@���3\�!?Ժ�Hp��@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@1&�ٿpʩ`��@�O��z�3@�<����!?�a�S�@-��֔ٿ��1���@b^��J�3@��5I�!?�}�$I6�@��Hx�ٿ�����0�@�k8j��3@����!? *���@?u�cƔٿ��g�P�@�;<��3@L�Sj��!?$Y���S�@�@k!��ٿ�f?8��@T�Κ��3@���M��!?F#h �@���Q�ٿ�a�����@�Ӭ!Q�3@[����!?(\��&�@���Q�ٿ�a�����@�Ӭ!Q�3@[����!?(\��&�@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@���%
�ٿ�������@�$�y��3@�I���!?�s�&~��@�t���ٿq?���N�@���m 4@�`w�,�!?_���!�@�t���ٿq?���N�@���m 4@�`w�,�!?_���!�@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�6)��ٿ�5�P"�@���4�3@�B7�@�!?X�g�C��@�d5b�ٿ�e��@��U<�3@�7]-�!?/��l�ʹ@�d5b�ٿ�e��@��U<�3@�7]-�!?/��l�ʹ@�d5b�ٿ�e��@��U<�3@�7]-�!?/��l�ʹ@1	�;��ٿ��,��x�@͸�Z��3@w��M�!?�jb�vմ@1	�;��ٿ��,��x�@͸�Z��3@w��M�!?�jb�vմ@1	�;��ٿ��,��x�@͸�Z��3@w��M�!?�jb�vմ@1	�;��ٿ��,��x�@͸�Z��3@w��M�!?�jb�vմ@���<�ٿ5Y%?�@�6�֖�3@��tV?�!?�́8
�@���<�ٿ5Y%?�@�6�֖�3@��tV?�!?�́8
�@���<�ٿ5Y%?�@�6�֖�3@��tV?�!?�́8
�@��p��ٿ����r�@�>��3@>�R)�!?�z8f�̴@��p��ٿ����r�@�>��3@>�R)�!?�z8f�̴@��p��ٿ����r�@�>��3@>�R)�!?�z8f�̴@��p��ٿ����r�@�>��3@>�R)�!?�z8f�̴@9�vm��ٿ%م�&�@�]�#�3@�C�"�!?1)k�Ci�@9�vm��ٿ%م�&�@�]�#�3@�C�"�!?1)k�Ci�@9�vm��ٿ%م�&�@�]�#�3@�C�"�!?1)k�Ci�@9�vm��ٿ%م�&�@�]�#�3@�C�"�!?1)k�Ci�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@.�=�E�ٿކZ�)��@2ӮZ�3@I����!?�'�=�I�@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@Z�-���ٿ�Y��.��@-��3@/��!?�_��@݆Ԗi�ٿ��X\��@i�Z�3@:����!?AX����@݆Ԗi�ٿ��X\��@i�Z�3@:����!?AX����@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@Ahz�ٿ�^��R&�@���ak�3@>�g��!?̼��K�@�JS8��ٿ�P ���@�Y����3@Tb8ER�!?;6�pǊ�@�JS8��ٿ�P ���@�Y����3@Tb8ER�!?;6�pǊ�@�JS8��ٿ�P ���@�Y����3@Tb8ER�!?;6�pǊ�@�JS8��ٿ�P ���@�Y����3@Tb8ER�!?;6�pǊ�@�JS8��ٿ�P ���@�Y����3@Tb8ER�!?;6�pǊ�@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@6}ޡ�ٿjb���)�@Q�I��3@��y�!?��Lx暵@���q,�ٿ�QȘ��@灜�o�3@����y�!?E�'ݢ��@���q,�ٿ�QȘ��@灜�o�3@����y�!?E�'ݢ��@���q,�ٿ�QȘ��@灜�o�3@����y�!?E�'ݢ��@���q,�ٿ�QȘ��@灜�o�3@����y�!?E�'ݢ��@���q,�ٿ�QȘ��@灜�o�3@����y�!?E�'ݢ��@����U�ٿ=К�He�@h&�֮�3@�*=�/�!?B�~}j�@*\z�ٿ�_d}l0�@��'��3@�d͢�!?�W��)�@*\z�ٿ�_d}l0�@��'��3@�d͢�!?�W��)�@*\z�ٿ�_d}l0�@��'��3@�d͢�!?�W��)�@*\z�ٿ�_d}l0�@��'��3@�d͢�!?�W��)�@�d�ٿ��/�
��@l)l6�3@q(ܫ�!?0ap�IV�@�d�ٿ��/�
��@l)l6�3@q(ܫ�!?0ap�IV�@����s�ٿ_+9��0�@���Wa4@Ȋ� p�!?�����@����s�ٿ_+9��0�@���Wa4@Ȋ� p�!?�����@Tcl1��ٿ��>��~�@�F�$4@�>R��!?C(���@Tcl1��ٿ��>��~�@�F�$4@�>R��!?C(���@E�|��ٿ�0���@${��4@H-��q�!?f!�ޡ�@E�|��ٿ�0���@${��4@H-��q�!?f!�ޡ�@�WG+�ٿ��K�0�@��o��3@=D�\��!?��<wܴ@�)��	�ٿ��%DY��@j5����3@���.�!?��@7>r�@�)��	�ٿ��%DY��@j5����3@���.�!?��@7>r�@�g57'�ٿ��[Y"�@[dپ�3@U厙*�!?۟`j�@�Q�վ�ٿGT�2��@�x�Y4@��<�`�!?=;.�B��@�Q�վ�ٿGT�2��@�x�Y4@��<�`�!?=;.�B��@�Q�վ�ٿGT�2��@�x�Y4@��<�`�!?=;.�B��@�Q�վ�ٿGT�2��@�x�Y4@��<�`�!?=;.�B��@B�TL}�ٿI�}ŏH�@b��4@KO�K�!?c���͵@�!:^��ٿ���=	�@�a|�54@��}�3�!?��r�m�@�!:^��ٿ���=	�@�a|�54@��}�3�!?��r�m�@�!:^��ٿ���=	�@�a|�54@��}�3�!?��r�m�@�!:^��ٿ���=	�@�a|�54@��}�3�!?��r�m�@�!:^��ٿ���=	�@�a|�54@��}�3�!?��r�m�@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@��z
ϓٿpn�ʊr�@��8++�3@�W>��!?����@���ٿpD�HO�@���`4@�%:���!?�m��� �@���ٿpD�HO�@���`4@�%:���!?�m��� �@�VE�^�ٿs����@ų}O�4@�D`�!?;�N���@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@��4r�ٿe�2���@W���4@TG�Y��!?H��z�Ӵ@�c!��ٿ
[�f��@{>s��4@�I9�!?h5�!�@�c!��ٿ
[�f��@{>s��4@�I9�!?h5�!�@
"���ٿb���@�SvE4@���w�!?b���쨴@
"���ٿb���@�SvE4@���w�!?b���쨴@
"���ٿb���@�SvE4@���w�!?b���쨴@wU�Ѡ�ٿ�� ^]�@&��P��3@f�/��!?��0���@wU�Ѡ�ٿ�� ^]�@&��P��3@f�/��!?��0���@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@����.�ٿn
�,��@V����4@w�p���!?�w(�W"�@2����ٿ�*�;�@5춆��3@599�4�!?��n�x�@2����ٿ�*�;�@5춆��3@599�4�!?��n�x�@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@Í��r�ٿ��	���@^F?���3@����U�!?�/��4��@vǖ�d�ٿ��X�>��@�_ ��3@n�u�!?^��rP�@vǖ�d�ٿ��X�>��@�_ ��3@n�u�!?^��rP�@vǖ�d�ٿ��X�>��@�_ ��3@n�u�!?^��rP�@vǖ�d�ٿ��X�>��@�_ ��3@n�u�!?^��rP�@!x,cO�ٿ�L4���@�?�\��3@�v:�R�!?�``��_�@!x,cO�ٿ�L4���@�?�\��3@�v:�R�!?�``��_�@!x,cO�ٿ�L4���@�?�\��3@�v:�R�!?�``��_�@!x,cO�ٿ�L4���@�?�\��3@�v:�R�!?�``��_�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@��qv�ٿd.��C��@V`�t�3@R*!|��!?�}�/�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@(!�s�ٿ} �sR��@�ƈh�3@���m��!?D��,�@�i��|�ٿGD;�C��@��Ёb�3@�:�䶐!?�������@�i��|�ٿGD;�C��@��Ёb�3@�:�䶐!?�������@�i��|�ٿGD;�C��@��Ёb�3@�:�䶐!?�������@�%��ٿ0pI���@���:�3@wE����!?|��@�%��ٿ0pI���@���:�3@wE����!?|��@�%��ٿ0pI���@���:�3@wE����!?|��@�%��ٿ0pI���@���:�3@wE����!?|��@�%��ٿ0pI���@���:�3@wE����!?|��@���o�ٿB�tqW�@�˶��3@nt�q�!?�yZ�ƴ@���o�ٿB�tqW�@�˶��3@nt�q�!?�yZ�ƴ@d��Vٿ%U=�
��@IV[�3@mE��!?f��vQ�@�M����ٿcl%-���@S��9��3@>��t�!? �eqA�@�M����ٿcl%-���@S��9��3@>��t�!? �eqA�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@[�i� �ٿ��yZ�@<s�5��3@uM/�!?��v`+(�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@�CE��ٿ�1xψ�@�(��, 4@�r@�!?Ǵ��%�@v<B6y�ٿ�ԫ���@�4@]�@��!?@_��C�@v<B6y�ٿ�ԫ���@�4@]�@��!?@_��C�@��J]D�ٿ�����@��IQm�3@��w���!?;��Q�I�@��J]D�ٿ�����@��IQm�3@��w���!?;��Q�I�@��J]D�ٿ�����@��IQm�3@��w���!?;��Q�I�@���ӕٿ̓�����@Y�ޥ	 4@�~�ۏ!?�+����@���ӕٿ̓�����@Y�ޥ	 4@�~�ۏ!?�+����@���ӕٿ̓�����@Y�ޥ	 4@�~�ۏ!?�+����@���ӕٿ̓�����@Y�ޥ	 4@�~�ۏ!?�+����@��ă�ٿ_]�2X�@X���4@��.�!?H��_Ɔ�@�?0���ٿC�B� ��@�wt��3@۰�V�!?�ѵx>�@�?0���ٿC�B� ��@�wt��3@۰�V�!?�ѵx>�@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@�?wn�ٿ�#�qߵ�@��|��3@�`!8�!?w~����@���[�ٿ�R:��@�(M'�3@�Y2�!?��s�z�@���[�ٿ�R:��@�(M'�3@�Y2�!?��s�z�@���[�ٿ�R:��@�(M'�3@�Y2�!?��s�z�@���[�ٿ�R:��@�(M'�3@�Y2�!?��s�z�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@Dŕ�E�ٿDHP��@U�jc�3@���~!�!?��{�q�@-NLZ8�ٿ+kY9;�@�D���3@�"��,�!?��1m.J�@b�,���ٿ�R���@��6���3@�^�"��!?Y�/�4G�@b�,���ٿ�R���@��6���3@�^�"��!?Y�/�4G�@
(s�o�ٿ 7u���@�0���3@��.�ǐ!?P�vT?�@
(s�o�ٿ 7u���@�0���3@��.�ǐ!?P�vT?�@
(s�o�ٿ 7u���@�0���3@��.�ǐ!?P�vT?�@
(s�o�ٿ 7u���@�0���3@��.�ǐ!?P�vT?�@
(s�o�ٿ 7u���@�0���3@��.�ǐ!?P�vT?�@dV���ٿ�n/8�P�@B�X���3@A��J��!?�L�T���@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@0L~7��ٿFt6[��@退�~�3@%����!?��I�:��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�U�n"�ٿ�<�t#r�@�i2�3@��I�!?r��6	��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@�ZE"�ٿ��{1Y��@x=�b��3@983�O�!?'�)��@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@wNa��ٿDhQ��@�~�/��3@P�[��!?urڈ�Ǵ@sA��L�ٿ����`J�@�	����3@m��*��!?�U·��@sA��L�ٿ����`J�@�	����3@m��*��!?�U·��@sA��L�ٿ����`J�@�	����3@m��*��!?�U·��@sA��L�ٿ����`J�@�	����3@m��*��!?�U·��@+.��w�ٿa$�qLv�@Tƕ*�3@oS�	e�!?��v��@+.��w�ٿa$�qLv�@Tƕ*�3@oS�	e�!?��v��@+.��w�ٿa$�qLv�@Tƕ*�3@oS�	e�!?��v��@+.��w�ٿa$�qLv�@Tƕ*�3@oS�	e�!?��v��@+.��w�ٿa$�qLv�@Tƕ*�3@oS�	e�!?��v��@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@L�ZX�ٿ|���I��@���A)�3@��X���!?�L���̴@F����ٿ&EZ|o��@���3@���^E�!?�߆�� �@��$
M�ٿ��|�N��@���D��3@�&m{�!?>��
E�@��$
M�ٿ��|�N��@���D��3@�&m{�!?>��
E�@��$
M�ٿ��|�N��@���D��3@�&m{�!?>��
E�@��$
M�ٿ��|�N��@���D��3@�&m{�!?>��
E�@������ٿ����k�@�=
���3@E���0�!?e
�fqH�@KQɿ_�ٿU�,W�9�@̺�n��3@�}"(b�!?s�-Te�@KQɿ_�ٿU�,W�9�@̺�n��3@�}"(b�!?s�-Te�@KQɿ_�ٿU�,W�9�@̺�n��3@�}"(b�!?s�-Te�@KQɿ_�ٿU�,W�9�@̺�n��3@�}"(b�!?s�-Te�@KQɿ_�ٿU�,W�9�@̺�n��3@�}"(b�!?s�-Te�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@t�˚�ٿJ*���}�@�����3@F��T^�!?.=e�$�@�':�ٿ�ף49��@!2��3@��w�!?<�.�E�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�����ٿ�tU���@}�8��4@�
�:�!?QL{��3�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@�H�G�ٿF�;�^�@����T	4@��M�E�!?�Ň��5�@F^�Q�ٿ�_0�Y�@�?w�x4@���i�!?y���JŴ@F^�Q�ٿ�_0�Y�@�?w�x4@���i�!?y���JŴ@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@e&�"דٿAM|����@feo�T�3@��Ш��!?�L��n�@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@b����ٿJ���9��@� t>� 4@� ��L�!?�K��QӴ@����ٿ��t,���@Jڳ���3@f?.g[�!?%�>�S�@����ٿ��t,���@Jڳ���3@f?.g[�!?%�>�S�@����ٿ��t,���@Jڳ���3@f?.g[�!?%�>�S�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@�zc��ٿy�S)���@�.U���3@������!?���Os�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@ث`��ٿxZ�&E!�@��o	o�3@�J�Є�!?�nԥaI�@���F��ٿ��6d�;�@��z*��3@�;��Z�!?O�n?�@���F��ٿ��6d�;�@��z*��3@�;��Z�!?O�n?�@���F��ٿ��6d�;�@��z*��3@�;��Z�!?O�n?�@9iM|:�ٿ�s���@<��~��3@���k�!?�5=\��@9iM|:�ٿ�s���@<��~��3@���k�!?�5=\��@z��A�ٿ��R?�@�����3@�$9�f�!?$[`��L�@���Q�ٿ��t��g�@'L{��3@0?T7��!?��'e�@;�R��ٿ��^c	�@���U�3@��&[�!?���É�@;�R��ٿ��^c	�@���U�3@��&[�!?���É�@*3v��ٿ��쏣�@�M���3@R���5�!?/я�-�@�`x]�ٿ|�*a4�@bE���3@_��J:�!?-�r���@�`x]�ٿ|�*a4�@bE���3@_��J:�!?-�r���@��3�ȗٿod��@��G�-�3@\�w9�!?J��y.c�@=�m{��ٿ �B�Zi�@�^)��3@\Q�e�!?3ڟ5��@i[��p�ٿ�8��	�@ˮr��3@ؓ��S�!?A���/�@�>B~�ٿs�&i6�@��Jw9�3@U��q=�!?1�!:�@�=)r�ٿ�._S���@p��b �3@A��Y�!?��&ѥ��@�=)r�ٿ�._S���@p��b �3@A��Y�!?��&ѥ��@�=)r�ٿ�._S���@p��b �3@A��Y�!?��&ѥ��@�=)r�ٿ�._S���@p��b �3@A��Y�!?��&ѥ��@�=)r�ٿ�._S���@p��b �3@A��Y�!?��&ѥ��@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@�x�Вٿ�,}��@�ބ�3@o�6<Z�!?�I��c�@ �6��ٿ����t�@b���3@�q��0�!?��aJ?��@����a�ٿ�Z�n ;�@G6��^�3@�9C��!?�*D��Y�@��iȐٿO��Զ��@v��?�3@ĉ�O��!?�}8���@��iȐٿO��Զ��@v��?�3@ĉ�O��!?�}8���@A��a��ٿt������@�XU�#�3@��ؽ�!?X�&v���@A��a��ٿt������@�XU�#�3@��ؽ�!?X�&v���@A��a��ٿt������@�XU�#�3@��ؽ�!?X�&v���@A��a��ٿt������@�XU�#�3@��ؽ�!?X�&v���@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@|�A�ٿ7D�����@Eu�?�3@ͼ*���!?����,�@�ݲ;�ٿ��\'�@_�[���3@�i�F/�!? |�e6�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@��!�ٿ��1�@�<��3@udX�!?���@"�@�\��ٿ'x^�C��@j
~���3@ІC�(�!?��:��@c�
�ٿuɬ��^�@�Q�6�3@�'"�8�!?��V8�@c�
�ٿuɬ��^�@�Q�6�3@�'"�8�!?��V8�@c�
�ٿuɬ��^�@�Q�6�3@�'"�8�!?��V8�@c�
�ٿuɬ��^�@�Q�6�3@�'"�8�!?��V8�@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@����ٿj,ͱ��@#�5��3@�A���!?���8��@���(�ٿP���@�$.y�3@�_�!?�(:��3�@$̙�ٿ��um��@�%m�R�3@�����!?�U�]�@$̙�ٿ��um��@�%m�R�3@�����!?�U�]�@$̙�ٿ��um��@�%m�R�3@�����!?�U�]�@$̙�ٿ��um��@�%m�R�3@�����!?�U�]�@p11ր�ٿ�}�5/��@#�/^�3@ k�,p�!?2�B�(�@���?-�ٿ]p���4�@@r�I�3@9/ ~��!?~տqK�@���?-�ٿ]p���4�@@r�I�3@9/ ~��!?~տqK�@���?-�ٿ]p���4�@@r�I�3@9/ ~��!?~տqK�@�ӧz��ٿ��G4��@�p����3@y;�9�!?Rژcش@�ӧz��ٿ��G4��@�p����3@y;�9�!?Rژcش@�aL�8�ٿ�k�.�@Neh&�3@�H��!?{�{=|E�@�aL�8�ٿ�k�.�@Neh&�3@�H��!?{�{=|E�@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@H��6�ٿ�QIw��@���%E�3@�q��	�!?�-���@���.՗ٿ��`M��@6���_�3@�K�#��!?.yZN���@���.՗ٿ��`M��@6���_�3@�K�#��!?.yZN���@���.՗ٿ��`M��@6���_�3@�K�#��!?.yZN���@���.՗ٿ��`M��@6���_�3@�K�#��!?.yZN���@WR���ٿN;kD�K�@0(�3�3@�#pH�!?�|�D0�@�R���ٿh�[�J�@i��jQ�3@��f�)�!?P&�"�@l��'�ٿ��=VS��@d8;=��3@/�o"[�!?1�x��@l��'�ٿ��=VS��@d8;=��3@/�o"[�!?1�x��@ ����ٿ&��!��@;�Y4@>�Şj�!?N�|@r�@ ����ٿ&��!��@;�Y4@>�Şj�!?N�|@r�@ ����ٿ&��!��@;�Y4@>�Şj�!?N�|@r�@ ����ٿ&��!��@;�Y4@>�Şj�!?N�|@r�@ ����ٿ&��!��@;�Y4@>�Şj�!?N�|@r�@Vݎ��ٿҰyu���@������3@@�ʐ!?m��}�[�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@5ϷVȚٿ{X��4�@^����3@C���F�!?ۇ��G�@��r=P�ٿ�\�2�-�@��ڋ��3@GpLvq�!?�����@��r=P�ٿ�\�2�-�@��ڋ��3@GpLvq�!?�����@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@P֏1͙ٿk�	7|��@F�4��3@;4q��!?��wL�@5<�ٿ���ػ��@�x�5,�3@&��!a�!?�4}�:�@5<�ٿ���ػ��@�x�5,�3@&��!a�!?�4}�:�@5<�ٿ���ػ��@�x�5,�3@&��!a�!?�4}�:�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@t�H��ٿ��ہ9�@���3@d�@�S�!?�B�}�@ݶ���ٿ*�z q��@~���3@A��;]�!?��	,���@ݶ���ٿ*�z q��@~���3@A��;]�!?��	,���@ݶ���ٿ*�z q��@~���3@A��;]�!?��	,���@ݶ���ٿ*�z q��@~���3@A��;]�!?��	,���@u����ٿ��bc S�@33���3@���V��!?�'�ǭ�@u����ٿ��bc S�@33���3@���V��!?�'�ǭ�@u����ٿ��bc S�@33���3@���V��!?�'�ǭ�@u����ٿ��bc S�@33���3@���V��!?�'�ǭ�@u����ٿ��bc S�@33���3@���V��!?�'�ǭ�@.Ѿ5I�ٿ4g�7��@,Cw�3@���T�!?�
EB�l�@.Ѿ5I�ٿ4g�7��@,Cw�3@���T�!?�
EB�l�@.Ѿ5I�ٿ4g�7��@,Cw�3@���T�!?�
EB�l�@.Ѿ5I�ٿ4g�7��@,Cw�3@���T�!?�
EB�l�@.Ѿ5I�ٿ4g�7��@,Cw�3@���T�!?�
EB�l�@%k;+^�ٿ���J~��@�yf*T�3@�nϏ!?2wO���@%k;+^�ٿ���J~��@�yf*T�3@�nϏ!?2wO���@%k;+^�ٿ���J~��@�yf*T�3@�nϏ!?2wO���@%k;+^�ٿ���J~��@�yf*T�3@�nϏ!?2wO���@%k;+^�ٿ���J~��@�yf*T�3@�nϏ!?2wO���@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@]����ٿ��A��:�@P����3@���ҏ!?:y�lK��@!��m��ٿ��fsu�@�/�=p�3@7����!?�"��۵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@[
�<m�ٿ��:�F��@�����3@8��'�!?/���켵@��	�!�ٿ��XG��@c��3@���$�!?�ee��@�@�n���ٿ�:/ ��@QΉd��3@�E���!?fiL\��@�n���ٿ�:/ ��@QΉd��3@�E���!?fiL\��@�n���ٿ�:/ ��@QΉd��3@�E���!?fiL\��@<�xl�ٿN�P��@Վ���3@f�gN�!?��Ng��@<�xl�ٿN�P��@Վ���3@f�gN�!?��Ng��@<�xl�ٿN�P��@Վ���3@f�gN�!?��Ng��@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@GU~,��ٿAh� y�@�|���3@x71*Ə!?������@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@G�$��ٿ�>�=Y�@nŴ���3@O��܏!?�g���@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@ b`�N�ٿ{�w���@��s(M4@o�Bϑ�!?^$7��@Z��?`�ٿ��y����@�2h�<4@~n��!?f	��Ǵ@Z��?`�ٿ��y����@�2h�<4@~n��!?f	��Ǵ@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@hť��ٿ�s�.�u�@�i�q��3@.yN��!?)�}��@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��Yf��ٿ�������@�^ 1��3@���2i�!?���D�3�@��!Ƙٿ�$��	%�@>�@���3@�]^��!?f�3|�@��!Ƙٿ�$��	%�@>�@���3@�]^��!?f�3|�@7G��@�ٿ��qI{h�@�@���3@\�6�1�!?_�3��@7G��@�ٿ��qI{h�@�@���3@\�6�1�!?_�3��@�!��ٿ�Y��3��@����Z4@��
Fx�!?6˳��0�@�!��ٿ�Y��3��@����Z4@��
Fx�!?6˳��0�@�!��ٿ�Y��3��@����Z4@��
Fx�!?6˳��0�@�!��ٿ�Y��3��@����Z4@��
Fx�!?6˳��0�@P���J�ٿ <mjZ�@U.�`��3@�)�v�!?+���~ִ@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@X4�	�ٿ�A0��@�$9*T�3@��cb�!?��?<�@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@ y���ٿC���i��@����3@��#�%�!?@���?׵@�7���ٿ,[�C&d�@*��<L�3@s�ɐ�!?��6YV�@�7���ٿ,[�C&d�@*��<L�3@s�ɐ�!?��6YV�@�4>��ٿ�A]z�:�@�n����3@4(��H�!?,Aq�ǵ@�4>��ٿ�A]z�:�@�n����3@4(��H�!?,Aq�ǵ@���ۜٿ�@����@�Aƴ�3@�b3!>�!?�|
���@���ۜٿ�@����@�Aƴ�3@�b3!>�!?�|
���@���ۜٿ�@����@�Aƴ�3@�b3!>�!?�|
���@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@��+N?�ٿi繋�J�@�����3@�7V+0�!?�t��4�@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@�6�ٿ��qWk�@O*���3@�� =�!?:�śKҵ@��-%�ٿ
�|��@����B�3@$��)�!?h�5��r�@��-%�ٿ
�|��@����B�3@$��)�!?h�5��r�@��-%�ٿ
�|��@����B�3@$��)�!?h�5��r�@�SA��ٿ}�L����@�����3@����K�!?v&��i�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��Js��ٿ���R��@�T�
��3@�C	��!?��?��=�@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@��w"��ٿ��{��@��v�3@��� �!?�cE����@H����ٿ�̩M�[�@�'��1�3@�-�{�!?�
_Wz�@H����ٿ�̩M�[�@�'��1�3@�-�{�!?�
_Wz�@H����ٿ�̩M�[�@�'��1�3@�-�{�!?�
_Wz�@H����ٿ�̩M�[�@�'��1�3@�-�{�!?�
_Wz�@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@��.:��ٿ�#J>�+�@V��h�3@
�vZ�!?No��N��@�����ٿ|rE�,�@y�tgp�3@���!?��wxŵ@ ����ٿ��2){��@�Ol��4@�����!?w�\ �@ ����ٿ��2){��@�Ol��4@�����!?w�\ �@ ����ٿ��2){��@�Ol��4@�����!?w�\ �@ ����ٿ��2){��@�Ol��4@�����!?w�\ �@ ����ٿ��2){��@�Ol��4@�����!?w�\ �@�j�ʈ�ٿv��`*��@��� r�3@�O��!?�R���@�j�ʈ�ٿv��`*��@��� r�3@�O��!?�R���@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@�?m�ٿAކ_�@�@�e�J��3@�T����!?4֟eK�@V����ٿM� W��@1�����3@t�����!?ze����@V����ٿM� W��@1�����3@t�����!?ze����@���ᥖٿ�8�"o<�@QJ̬�3@��R��!?__�0��@���ᥖٿ�8�"o<�@QJ̬�3@��R��!?__�0��@���ᥖٿ�8�"o<�@QJ̬�3@��R��!?__�0��@���ᥖٿ�8�"o<�@QJ̬�3@��R��!?__�0��@��mM��ٿ>C,Ĝ�@+�u��3@�Pw�0�!?P�����@5�6ϣ�ٿF(��@��m�3@���u	�!?U�:�C�@5�6ϣ�ٿF(��@��m�3@���u	�!?U�:�C�@#s�Fߞٿ�u�{�@jk����3@˨<��!?W�E�&�@�*`��ٿ����I�@ӫ�r<�3@��Iq2�!?*�Kw�@uq	�ٿȽR-4��@k����4@�����!?(�>G���@uq	�ٿȽR-4��@k����4@�����!?(�>G���@uq	�ٿȽR-4��@k����4@�����!?(�>G���@uq	�ٿȽR-4��@k����4@�����!?(�>G���@�y��ٿZ�'�Ĥ�@v�R_�3@k:
��!?X�LB�=�@�y��ٿZ�'�Ĥ�@v�R_�3@k:
��!?X�LB�=�@�y��ٿZ�'�Ĥ�@v�R_�3@k:
��!?X�LB�=�@��؀��ٿ�q-1b�@�r>>|�3@�Q(r�!?�eʞ���@r`dΖٿ~��@=���3@L�nD�!?�}��iԵ@r`dΖٿ~��@=���3@L�nD�!?�}��iԵ@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�穖ٿ��8]�@	�N���3@V�RU�!?ӽ�����@�	a#��ٿ�d�V�@�r���3@M� ��!?���Z>z�@�	a#��ٿ�d�V�@�r���3@M� ��!?���Z>z�@�	a#��ٿ�d�V�@�r���3@M� ��!?���Z>z�@�O�)��ٿ�����@#�)�m�3@��/̎�!?=ځ ��@�O�)��ٿ�����@#�)�m�3@��/̎�!?=ځ ��@�����ٿ�ځ�Ձ�@��5�3@��q��!?֦s��@��y���ٿ�{����@��\4@���IP�!?����⁵@��y���ٿ�{����@��\4@���IP�!?����⁵@��y���ٿ�{����@��\4@���IP�!?����⁵@��y���ٿ�{����@��\4@���IP�!?����⁵@5��X��ٿ'��9Zh�@�-}Z+4@��:X�!?��\��@5��X��ٿ'��9Zh�@�-}Z+4@��:X�!?��\��@5��X��ٿ'��9Zh�@�-}Z+4@��:X�!?��\��@5��X��ٿ'��9Zh�@�-}Z+4@��:X�!?��\��@�r�m��ٿ��َ��@�@<�I4@�,��!?����I�@��셡ٿ�fQ�@"8�Z�3@\F�-4�!?7Τ����@��셡ٿ�fQ�@"8�Z�3@\F�-4�!?7Τ����@��셡ٿ�fQ�@"8�Z�3@\F�-4�!?7Τ����@��셡ٿ�fQ�@"8�Z�3@\F�-4�!?7Τ����@�<60z�ٿD�
��@��f͒�3@,>�V �!?n���+�@����ޘٿ�c�P�@��"��3@.�S�w�!?�}�y�=�@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@L��ٿ�[!W��@:���3@���c<�!?T%6�qԴ@�JJ���ٿ�p�Ǧ��@7@��a�3@�L��V�!?3$+1ώ�@��k�?�ٿ<EѺ#�@��]�n�3@�u��!?VjA�c%�@��k�?�ٿ<EѺ#�@��]�n�3@�u��!?VjA�c%�@:��~��ٿ���G7�@�UD��3@2:�^�!?�h}�b�@:��~��ٿ���G7�@�UD��3@2:�^�!?�h}�b�@:��~��ٿ���G7�@�UD��3@2:�^�!?�h}�b�@:��~��ٿ���G7�@�UD��3@2:�^�!?�h}�b�@:��~��ٿ���G7�@�UD��3@2:�^�!?�h}�b�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@�|��ٿ��-Lw�@�ⴗ��3@�"i}�!?q��MI�@('���ٿ)�buY�@+�+��3@`���!?��qHz��@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@����ٿI�3�+�@܇��M 4@%���j�!?�+�\�
�@�=��ٿ���jY�@S8V���3@���:�!?��y�r״@U�U���ٿ�ի�[�@d^���3@V��Mo�!?`c;����@U�U���ٿ�ի�[�@d^���3@V��Mo�!?`c;����@U�U���ٿ�ի�[�@d^���3@V��Mo�!?`c;����@U�U���ٿ�ի�[�@d^���3@V��Mo�!?`c;����@:�)��ٿ3km�<�@@����3@]��ߥ�!?%Za�@�@:�)��ٿ3km�<�@@����3@]��ߥ�!?%Za�@�@:�)��ٿ3km�<�@@����3@]��ߥ�!?%Za�@�@�U��E�ٿ�`E�+<�@�k��3@@�UꞐ!?" ���@�U��E�ٿ�`E�+<�@�k��3@@�UꞐ!?" ���@��F�ٿ�Xs���@���3@*`�8&�!?�vߎ�@�c��Θٿؤ�>���@����3@�Xa��!?zu��)�@�c��Θٿؤ�>���@����3@�Xa��!?zu��)�@�c��Θٿؤ�>���@����3@�Xa��!?zu��)�@�c��Θٿؤ�>���@����3@�Xa��!?zu��)�@�c��Θٿؤ�>���@����3@�Xa��!?zu��)�@[L�d�ٿ�����@yD�4@@�R'�!?�5(+>+�@[L�d�ٿ�����@yD�4@@�R'�!?�5(+>+�@[L�d�ٿ�����@yD�4@@�R'�!?�5(+>+�@[L�d�ٿ�����@yD�4@@�R'�!?�5(+>+�@l�C��ٿ�>&o��@}�����3@��!?�)g�)�@l�C��ٿ�>&o��@}�����3@��!?�)g�)�@}��ٿG�qh�;�@K��o4@�oT?�!?�D+k�@�<n�8�ٿ�^v��@`Cp��3@��u�!?R�>�@�<n�8�ٿ�^v��@`Cp��3@��u�!?R�>�@�<n�8�ٿ�^v��@`Cp��3@��u�!?R�>�@�<n�8�ٿ�^v��@`Cp��3@��u�!?R�>�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@��-�ٿV����@t��Q�3@`h��!?�!��n�@8"`���ٿ�ߗ��s�@��V�3@a]��Ï!?����@8"`���ٿ�ߗ��s�@��V�3@a]��Ï!?����@8"`���ٿ�ߗ��s�@��V�3@a]��Ï!?����@8"`���ٿ�ߗ��s�@��V�3@a]��Ï!?����@jl�Țٿ �|��@_�
�3@�n�ԏ!?�ƽE܎�@jl�Țٿ �|��@_�
�3@�n�ԏ!?�ƽE܎�@jl�Țٿ �|��@_�
�3@�n�ԏ!?�ƽE܎�@jl�Țٿ �|��@_�
�3@�n�ԏ!?�ƽE܎�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@�:��ٿ���@B5�%��3@�
�XI�!?�mDƣ�@[�}�U�ٿ��V�ߧ�@�ؖv��3@�Fh�!?���f3 �@[�}�U�ٿ��V�ߧ�@�ؖv��3@�Fh�!?���f3 �@[�}�U�ٿ��V�ߧ�@�ؖv��3@�Fh�!?���f3 �@[�}�U�ٿ��V�ߧ�@�ؖv��3@�Fh�!?���f3 �@[�}�U�ٿ��V�ߧ�@�ؖv��3@�Fh�!?���f3 �@5�R��ٿ-A|j��@��e���3@�N�e��!?��罸B�@;N��L�ٿ�|�UT�@:�XW�3@��'@֏!?CdL-�ٴ@;N��L�ٿ�|�UT�@:�XW�3@��'@֏!?CdL-�ٴ@;N��L�ٿ�|�UT�@:�XW�3@��'@֏!?CdL-�ٴ@;N��L�ٿ�|�UT�@:�XW�3@��'@֏!?CdL-�ٴ@,�v�K�ٿ�*O�D�@�~jA]4@~!�\�!?����˴@�����ٿz�3~��@���4@����_�!?�Y_�ˈ�@�����ٿz�3~��@���4@����_�!?�Y_�ˈ�@�����ٿz�3~��@���4@����_�!?�Y_�ˈ�@	q|}ݔٿ�Ǫ6C��@�"��	4@�g�8�!?4�X�е@	q|}ݔٿ�Ǫ6C��@�"��	4@�g�8�!?4�X�е@�,Ɓ�ٿ֕G�R.�@��Q4@.��h/�!?jJ���Ƶ@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@4�`�ٿϲ��E�@��Z���3@�U�-�!?Q"�!�@�o���ٿK�[�@D�h�3@L�2>K�!?��V�jD�@�o���ٿK�[�@D�h�3@L�2>K�!?��V�jD�@�o���ٿK�[�@D�h�3@L�2>K�!?��V�jD�@�o���ٿK�[�@D�h�3@L�2>K�!?��V�jD�@�o���ٿK�[�@D�h�3@L�2>K�!?��V�jD�@��ٜٿ�p^&�\�@{�`�$4@�7�!?':��$�@��ٜٿ�p^&�\�@{�`�$4@�7�!?':��$�@��ٜٿ�p^&�\�@{�`�$4@�7�!?':��$�@��n��ٿl״Y��@+�^�[�3@^����!?�;����@��n��ٿl״Y��@+�^�[�3@^����!?�;����@��@���ٿ2@� X�@x|���3@����!?r��f�[�@��@���ٿ2@� X�@x|���3@����!?r��f�[�@��@���ٿ2@� X�@x|���3@����!?r��f�[�@��@���ٿ2@� X�@x|���3@����!?r��f�[�@���Bg�ٿ�Jw���@Z���3@c���-�!?�
��@���Bg�ٿ�Jw���@Z���3@c���-�!?�
��@�f��ٿ��='���@Q͆���3@��[o�!?�|���@�f��ٿ��='���@Q͆���3@��[o�!?�|���@�f��ٿ��='���@Q͆���3@��[o�!?�|���@�f��ٿ��='���@Q͆���3@��[o�!?�|���@�f��ٿ��='���@Q͆���3@��[o�!?�|���@���O�ٿk�F���@�Ѽ ��3@��;��!?Rm-��@���O�ٿk�F���@�Ѽ ��3@��;��!?Rm-��@�6hA�ٿ�l��j��@��)�3@:Tj�8�!?c���e�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@��v���ٿ�"��f��@����a�3@FU�0�!?���q!Z�@����[�ٿk��1��@L��$V�3@���ֈ�!?"uz%2�@����[�ٿk��1��@L��$V�3@���ֈ�!?"uz%2�@����[�ٿk��1��@L��$V�3@���ֈ�!?"uz%2�@����ٿ�`G�м�@�FG~��3@U�}^�!?�Rdf��@����ٿ�`G�м�@�FG~��3@U�}^�!?�Rdf��@����ٿ�`G�м�@�FG~��3@U�}^�!?�Rdf��@�i�H�ٿE$�#��@&:X�1�3@[�=�u�!?FZ,��@2�x�ٿcP|�@�餐��3@�� 8�!?�,k�I��@�9���ٿW
.��@�c��`�3@D/�1�!?E?��b�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@^[��ٿKx���@ԫ��?�3@{Aʂ�!?wZg_H�@j���ٿ�	�Ƹ��@+�yy�3@C�nڜ�!?�i����@܃���ٿ��_%$*�@ ���3@-���!?c�ȹ�@܃���ٿ��_%$*�@ ���3@-���!?c�ȹ�@܃���ٿ��_%$*�@ ���3@-���!?c�ȹ�@܃���ٿ��_%$*�@ ���3@-���!?c�ȹ�@܃���ٿ��_%$*�@ ���3@-���!?c�ȹ�@tsՕٿp���tM�@��-�f�3@̡���!?�[qj`�@������ٿi{���@
���d�3@u�����!?������@������ٿi{���@
���d�3@u�����!?������@������ٿi{���@
���d�3@u�����!?������@������ٿi{���@
���d�3@u�����!?������@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@��@�M�ٿ���h��@ẕ���3@��vb��!?�%g�@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@߳荎�ٿ!�[�=�@f%�
�3@}��!?�K�s	ߴ@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�7L�r�ٿy��|��@��p���3@;��	�!?�m�C�t�@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�w�iG�ٿ�J��.��@$����3@�dP i�!?Z'`7P��@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�ߜ���ٿ4�v}��@�dG�3@t1R�&�!?��:j�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@�=ۉ�ٿ�H��`A�@�HN!R�3@c
��!?4p��Q�@��~�ٿ|��0D,�@���3@l�^���!? $mC*�@q�{�ސٿ��Q�s�@YȖi��3@H�e�<�!?�F�^E[�@8���ݓٿ�A�K�_�@#s��&�3@N�i��!?�긡���@8���ݓٿ�A�K�_�@#s��&�3@N�i��!?�긡���@8���ݓٿ�A�K�_�@#s��&�3@N�i��!?�긡���@8���ݓٿ�A�K�_�@#s��&�3@N�i��!?�긡���@8���ݓٿ�A�K�_�@#s��&�3@N�i��!?�긡���@c�A��ٿ3"ə�@V�����3@�o��*�!?R��#�@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�X�8�ٿ��/痵�@� %��3@zOF�]�!?�ū��ĵ@�[k[�ٿ|ev	}�@�V����3@�Yu�q�!?�kR� P�@�[k[�ٿ|ev	}�@�V����3@�Yu�q�!?�kR� P�@�[k[�ٿ|ev	}�@�V����3@�Yu�q�!?�kR� P�@�[k[�ٿ|ev	}�@�V����3@�Yu�q�!?�kR� P�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@:G��ٿ#Ӟ`��@s�����3@w��c�!?LP��W�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@!&m�ٿ��u����@�
,:.�3@4��c��!?|��<�@��MJ-�ٿwzc'�@c)UA�3@�u v��!?6N���@��MJ-�ٿwzc'�@c)UA�3@�u v��!?6N���@��MJ-�ٿwzc'�@c)UA�3@�u v��!?6N���@��MJ-�ٿwzc'�@c)UA�3@�u v��!?6N���@��MJ-�ٿwzc'�@c)UA�3@�u v��!?6N���@k���ٿGi�8j��@4��#6�3@|`pKv�!?�sRѡ+�@k���ٿGi�8j��@4��#6�3@|`pKv�!?�sRѡ+�@�'���ٿd�.�u�@��
W��3@h����!?q���Դ@�'���ٿd�.�u�@��
W��3@h����!?q���Դ@�'���ٿd�.�u�@��
W��3@h����!?q���Դ@���]��ٿ�M'����@��@�i4@�2e<�!?S��Q�@���]��ٿ�M'����@��@�i4@�2e<�!?S��Q�@���]��ٿ�M'����@��@�i4@�2e<�!?S��Q�@���]��ٿ�M'����@��@�i4@�2e<�!?S��Q�@���]��ٿ�M'����@��@�i4@�2e<�!?S��Q�@!G���ٿ��S���@C�����3@��H�!?�,�����@!G���ٿ��S���@C�����3@��H�!?�,�����@!G���ٿ��S���@C�����3@��H�!?�,�����@!G���ٿ��S���@C�����3@��H�!?�,�����@�9,��ٿ�>�B��@�%=/m�3@��9�!?]a�S��@�9,��ٿ�>�B��@�%=/m�3@��9�!?]a�S��@�9,��ٿ�>�B��@�%=/m�3@��9�!?]a�S��@�9,��ٿ�>�B��@�%=/m�3@��9�!?]a�S��@�9,��ٿ�>�B��@�%=/m�3@��9�!?]a�S��@J͐�ٿ�l0ųD�@6�C��3@�4����!?��E��@J͐�ٿ�l0ųD�@6�C��3@�4����!?��E��@J͐�ٿ�l0ųD�@6�C��3@�4����!?��E��@J͐�ٿ�l0ųD�@6�C��3@�4����!?��E��@�S�?��ٿ��� I�@p��T�4@9Sr��!?IҌ=c�@i��#�ٿ<T=�G�@Aǥg!4@�,}Ɛ!?�di�gU�@i��#�ٿ<T=�G�@Aǥg!4@�,}Ɛ!?�di�gU�@i��#�ٿ<T=�G�@Aǥg!4@�,}Ɛ!?�di�gU�@�R�`9�ٿ拭C8��@��^Y�3@��;߀�!?3�k��@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@���|ӑٿ��-H�@��)��3@e�Ξ�!?&�ۑ�@�kl���ٿpe�U
�@�k�'��3@Mxk�\�!?����ʹ@�kl���ٿpe�U
�@�k�'��3@Mxk�\�!?����ʹ@ALv��ٿ�O<�C��@�e���3@�/���!?r�ԫ��@ALv��ٿ�O<�C��@�e���3@�/���!?r�ԫ��@ALv��ٿ�O<�C��@�e���3@�/���!?r�ԫ��@ALv��ٿ�O<�C��@�e���3@�/���!?r�ԫ��@ALv��ٿ�O<�C��@�e���3@�/���!?r�ԫ��@�g�@�ٿ*(�� �@��=�?�3@��%�!?���kx�@�g�@�ٿ*(�� �@��=�?�3@��%�!?���kx�@�g�@�ٿ*(�� �@��=�?�3@��%�!?���kx�@�g�@�ٿ*(�� �@��=�?�3@��%�!?���kx�@�g�@�ٿ*(�� �@��=�?�3@��%�!?���kx�@t�+�\�ٿ���W"�@�E����3@���# �!?��,����@t�+�\�ٿ���W"�@�E����3@���# �!?��,����@���x��ٿ�~�8��@d׎w�3@�W+�!?!��/,��@�ӑ��ٿ���0�Z�@ҫ���3@=�<I�!?7�?B?�@�ӑ��ٿ���0�Z�@ҫ���3@=�<I�!?7�?B?�@�ӑ��ٿ���0�Z�@ҫ���3@=�<I�!?7�?B?�@�ӑ��ٿ���0�Z�@ҫ���3@=�<I�!?7�?B?�@�ӑ��ٿ���0�Z�@ҫ���3@=�<I�!?7�?B?�@x���	�ٿUZe�n�@?���3@����o�!?a�/�8�@���7�ٿ�8��R��@��~�3@#q�=�!?�m�Aት@~�/��ٿ�'B#��@�r�^��3@�w� �!?R^(��z�@~�/��ٿ�'B#��@�r�^��3@�w� �!?R^(��z�@~�/��ٿ�'B#��@�r�^��3@�w� �!?R^(��z�@~�/��ٿ�'B#��@�r�^��3@�w� �!?R^(��z�@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@7���"�ٿ�����@�R�v4@�v7 �!?����Z��@b6ZG��ٿ 	6Oe��@ ����3@��ؓa�!?�V��#*�@t�O?R�ٿ��Yo�@�*��U�3@H�}ɐ!?X�+��z�@t�O?R�ٿ��Yo�@�*��U�3@H�}ɐ!?X�+��z�@t�O?R�ٿ��Yo�@�*��U�3@H�}ɐ!?X�+��z�@t�O?R�ٿ��Yo�@�*��U�3@H�}ɐ!?X�+��z�@t�O?R�ٿ��Yo�@�*��U�3@H�}ɐ!?X�+��z�@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@���8m�ٿG�����@�h�>4@S��U�!?��UG �@w^��ٿW�
X!�@~�)��3@c��pz�!?�b�N�P�@w^��ٿW�
X!�@~�)��3@c��pz�!?�b�N�P�@w^��ٿW�
X!�@~�)��3@c��pz�!?�b�N�P�@w^��ٿW�
X!�@~�)��3@c��pz�!?�b�N�P�@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@�����ٿ�t�_��@TL��B�3@�)j��!?[����@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@ś�ǟ�ٿ�MZ�@?�"�3@�
5�T�!?:�Tm1�@�dgˑٿ�����@\oa�3@�UFp�!?��W��#�@�dgˑٿ�����@\oa�3@�UFp�!?��W��#�@�dgˑٿ�����@\oa�3@�UFp�!?��W��#�@�dgˑٿ�����@\oa�3@�UFp�!?��W��#�@��s
��ٿ��a,�$�@�A���4@�gR��!?�*e��=�@��s
��ٿ��a,�$�@�A���4@�gR��!?�*e��=�@�t"�p�ٿ�p�j�@IAܧ�3@R�%Gg�!?�$]�x�@�t"�p�ٿ�p�j�@IAܧ�3@R�%Gg�!?�$]�x�@�t"�p�ٿ�p�j�@IAܧ�3@R�%Gg�!?�$]�x�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@[Bj%�ٿ��.CB��@����4@Q����!?I�"0G�@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@��e���ٿ��9-��@/�qu��3@K#��.�!?�؅I� �@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@X�_ݕٿ�Aw���@M����3@�ZtX�!?�//r.�@ǵ�+�ٿ����@Z���$�3@R��9�!?v�
=G�@u*�o��ٿ��=�O�@��-�	�3@�a�
~�!?*e{u5(�@u*�o��ٿ��=�O�@��-�	�3@�a�
~�!?*e{u5(�@�(��s�ٿ����@�eC���3@>!?'�{�д@�:��E�ٿ�24���@)F1�J�3@��[&�!?��fq?�@)�|��ٿ-�ie5[�@���$�3@GGZk�!?ޚI����@F:�1�ٿ��p��@���3@?`�'��!?,V�	�@F:�1�ٿ��p��@���3@?`�'��!?,V�	�@F:�1�ٿ��p��@���3@?`�'��!?,V�	�@MA�5��ٿ�(�����@6[~�K�3@y�oȇ�!?���մ@MA�5��ٿ�(�����@6[~�K�3@y�oȇ�!?���մ@MA�5��ٿ�(�����@6[~�K�3@y�oȇ�!?���մ@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@���M��ٿ2�����@[�~�3@�Nu
�!?�cAʹ��@)��;�ٿBƲm��@v�����3@&�1�?�!?����D�@)��;�ٿBƲm��@v�����3@&�1�?�!?����D�@��B��ٿ��Q����@m^|�3@�&h	�!?�kC> �@В�(ؗٿ4<xO|�@u��V��3@9|���!?]�y�W�@В�(ؗٿ4<xO|�@u��V��3@9|���!?]�y�W�@В�(ؗٿ4<xO|�@u��V��3@9|���!?]�y�W�@>gE��ٿG2P���@Q1�3@���m�!?��P���@>gE��ٿG2P���@Q1�3@���m�!?��P���@>gE��ٿG2P���@Q1�3@���m�!?��P���@"mE�ٿ�BGK�@�R�t��3@2�[?�!?�*g��@���s�ٿ#�֚E��@�^}�3@u�R�I�!?��1��@���s�ٿ#�֚E��@�^}�3@u�R�I�!?��1��@���s�ٿ#�֚E��@�^}�3@u�R�I�!?��1��@���s�ٿ#�֚E��@�^}�3@u�R�I�!?��1��@���s�ٿ#�֚E��@�^}�3@u�R�I�!?��1��@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@�A���ٿt/�PiA�@o�t��3@�E"���!?ҵ3�42�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@� V�ٿ�yTXi��@�����3@�9�k�!?�ŉ�*�@#�퉐�ٿ^j����@�Z��3@���C�!?�4k�@#�퉐�ٿ^j����@�Z��3@���C�!?�4k�@#�퉐�ٿ^j����@�Z��3@���C�!?�4k�@#�퉐�ٿ^j����@�Z��3@���C�!?�4k�@  [P�ٿ�s����@�)���3@�I�k�!?w��?YU�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@=�s2_�ٿ��4���@(�����3@�^o�!?�rQQ	U�@�.붚ٿ;�k#�@�,Ĩ}�3@�� ��!?���A�@��RgK�ٿ�Xh4��@�$�%��3@8;�U�!?�M��p�@��RgK�ٿ�Xh4��@�$�%��3@8;�U�!?�M��p�@"v@���ٿ��N/P�@�X'r�3@�R�~�!?��̀��@7z;ɜٿ��Ce���@���3@*I�!?���@x?�ٿ���~<��@�#95�3@7�.�!?���\�z�@m��e�ٿ�6H8*"�@n> � 4@L�6�#�!?�3
I��@m��e�ٿ�6H8*"�@n> � 4@L�6�#�!?�3
I��@m��e�ٿ�6H8*"�@n> � 4@L�6�#�!?�3
I��@X+�0�ٿ����P�@��7z�3@{����!?zԌ��ִ@X+�0�ٿ����P�@��7z�3@{����!?zԌ��ִ@X+�0�ٿ����P�@��7z�3@{����!?zԌ��ִ@E���}�ٿ,e�5� �@[i�N 4@x�?�F�!?��a�Ƈ�@E���}�ٿ,e�5� �@[i�N 4@x�?�F�!?��a�Ƈ�@E���}�ٿ,e�5� �@[i�N 4@x�?�F�!?��a�Ƈ�@*��ߓٿT]k���@F��W�4@�g홁�!?��`!�G�@*��ߓٿT]k���@F��W�4@�g홁�!?��`!�G�@*��ߓٿT]k���@F��W�4@�g홁�!?��`!�G�@*��ߓٿT]k���@F��W�4@�g홁�!?��`!�G�@�� $r�ٿq�D�<M�@�}���3@�QV�9�!?u��� �@���ߓٿ��>���@�;�:��3@��oD�!?� 
�#�@���ߓٿ��>���@�;�:��3@��oD�!?� 
�#�@g�+��ٿg�I�f��@s?b�A�3@g�1/7�!?�k��Ե@+|����ٿI��'�@hŚް�3@1���[�!?�i�X�N�@+|����ٿI��'�@hŚް�3@1���[�!?�i�X�N�@+|����ٿI��'�@hŚް�3@1���[�!?�i�X�N�@8{.G��ٿ�~V��@��b�3@���?o�!?�a�0��@���ٿ��Ј��@���_S�3@�˭���!?2�E��@���ٿ��Ј��@���_S�3@�˭���!?2�E��@[�`���ٿ��^�S�@9�����3@�נ<w�!?H+�Xx�@[�`���ٿ��^�S�@9�����3@�נ<w�!?H+�Xx�@[�`���ٿ��^�S�@9�����3@�נ<w�!?H+�Xx�@�~$�
�ٿ0�*P'�@b�q�l�3@�=�ƍ�!?SaX�o�@�~$�
�ٿ0�*P'�@b�q�l�3@�=�ƍ�!?SaX�o�@�~$�
�ٿ0�*P'�@b�q�l�3@�=�ƍ�!?SaX�o�@���@�ٿ���O�R�@�"v�E�3@�	�Iv�!??<�T$�@���@�ٿ���O�R�@�"v�E�3@�	�Iv�!??<�T$�@���@�ٿ���O�R�@�"v�E�3@�	�Iv�!??<�T$�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@̥���ٿX��
&�@�f�HV�3@*8a�!?YZ�UW�@N�ƒ=�ٿB�x�@�]v�3@ &�sI�!?kc�9s�@N�ƒ=�ٿB�x�@�]v�3@ &�sI�!?kc�9s�@v[
�ٿ��w�ϛ�@�#��4@7"�@�!?��s��@v[
�ٿ��w�ϛ�@�#��4@7"�@�!?��s��@�)�L$�ٿ�eˍ�@��8���3@z��!?!@F�(1�@�)�L$�ٿ�eˍ�@��8���3@z��!?!@F�(1�@�)�L$�ٿ�eˍ�@��8���3@z��!?!@F�(1�@��H�4�ٿNŲ���@b0�E�3@�F2��!?�ի�!�@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@WWT:��ٿOUH�i�@�����3@���d�!?�2�Y��@5Y��(�ٿ���j2�@�:���3@�K,|�!?�R�v;�@5Y��(�ٿ���j2�@�:���3@�K,|�!?�R�v;�@��� �ٿ��{�%��@������3@fNL�!?��}g��@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@����ٿ_@����@�q{�3@ 8�!�!?� ��l
�@��I�F�ٿ��o�%��@y�M���3@D�m�X�!?VI��@��I�F�ٿ��o�%��@y�M���3@D�m�X�!?VI��@��I�F�ٿ��o�%��@y�M���3@D�m�X�!?VI��@���t��ٿDNJ��%�@���*k�3@uK��Q�!?��i���@���t��ٿDNJ��%�@���*k�3@uK��Q�!?��i���@���t��ٿDNJ��%�@���*k�3@uK��Q�!?��i���@���t��ٿDNJ��%�@���*k�3@uK��Q�!?��i���@���t��ٿDNJ��%�@���*k�3@uK��Q�!?��i���@��H��ٿ��¢~=�@7��=��3@�?"=�!?�9����@��H��ٿ��¢~=�@7��=��3@�?"=�!?�9����@�KK�"�ٿ��,�]�@�8�H�3@B��6�!?���*�@�KK�"�ٿ��,�]�@�8�H�3@B��6�!?���*�@�KK�"�ٿ��,�]�@�8�H�3@B��6�!?���*�@.��e��ٿ�|��@�=}��3@f�T@�!?��޿Z^�@7��J�ٿ�=#3��@��T"2�3@b}�=�!?X��@7��J�ٿ�=#3��@��T"2�3@b}�=�!?X��@^ജ�ٿF����@��L��3@�6E�1�!?&�C�@^ജ�ٿF����@��L��3@�6E�1�!?&�C�@^ജ�ٿF����@��L��3@�6E�1�!?&�C�@7]3��ٿI2�9S�@�́t��3@��ھI�!?ý,y��@7]3��ٿI2�9S�@�́t��3@��ھI�!?ý,y��@7]3��ٿI2�9S�@�́t��3@��ھI�!?ý,y��@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@��
p��ٿ��/</�@~�K��3@��
���!?�{VJѴ@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@�NLHҒٿ{��Yy�@�A���3@WK�e��!?�x�Ѓ��@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@���zٿ_"�����@u�_D��3@��b�W�!?@�3~䡴@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@V�!hܔٿ=
D�c1�@Q~y��3@,���c�!?P�->��@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@E{_�p�ٿ+�_���@uo�R"�3@K/v�a�!?nK2ᱴ@�x�U�ٿJ^,�Bk�@&��sc�3@Ŋ�H�!?Mj!�'��@�x�U�ٿJ^,�Bk�@&��sc�3@Ŋ�H�!?Mj!�'��@�x�U�ٿJ^,�Bk�@&��sc�3@Ŋ�H�!?Mj!�'��@�x�U�ٿJ^,�Bk�@&��sc�3@Ŋ�H�!?Mj!�'��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@��q��ٿ�(�Y�@�u�W�3@�X�h�!?{wu��@�s��ٿ��@?�@�CG���3@�t� 6�!?0��O��@�s��ٿ��@?�@�CG���3@�t� 6�!?0��O��@�s��ٿ��@?�@�CG���3@�t� 6�!?0��O��@����ٿ߇W���@��vU��3@�\gᩐ!?ɖ���`�@����ٿ߇W���@��vU��3@�\gᩐ!?ɖ���`�@�Vޤ	�ٿS9�J�!�@Jv3��3@��"���!?
���z�@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�w�gV�ٿ�G��A~�@�pM���3@�^P��!?�&"�.��@�~c�ٿ�Q�Y��@�k����3@��זl�!?]��;@�@�~c�ٿ�Q�Y��@�k����3@��זl�!?]��;@�@�~c�ٿ�Q�Y��@�k����3@��זl�!?]��;@�@�~c�ٿ�Q�Y��@�k����3@��זl�!?]��;@�@�~c�ٿ�Q�Y��@�k����3@��זl�!?]��;@�@D��N�ٿ��H�p�@�]���3@.��?��!?���<��@D��N�ٿ��H�p�@�]���3@.��?��!?���<��@D��N�ٿ��H�p�@�]���3@.��?��!?���<��@D��N�ٿ��H�p�@�]���3@.��?��!?���<��@bl"�K�ٿkJ�x���@��ox�3@���Ǡ�!?�I|�&�@Xx7�ٿ��z����@��q�3@>~*�А!?�D�8µ@Xx7�ٿ��z����@��q�3@>~*�А!?�D�8µ@Xx7�ٿ��z����@��q�3@>~*�А!?�D�8µ@Xx7�ٿ��z����@��q�3@>~*�А!?�D�8µ@���#o�ٿ�F�YW[�@�d�%h4@�a 
��!?����۵@���#o�ٿ�F�YW[�@�d�%h4@�a 
��!?����۵@���6%�ٿ�? �s�@�o����3@�hĥ}�!?D��_�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@�{O�ٿ��2�RZ�@���K�3@���M�!?���e�"�@��``��ٿ��'a�@v����3@��	�&�!?L:����@��``��ٿ��'a�@v����3@��	�&�!?L:����@=�q��ٿĸ���g�@ �#`�3@����!?�i�HԴ@=�q��ٿĸ���g�@ �#`�3@����!?�i�HԴ@�����ٿ��A�Nn�@����3@9�z^O�!?t�F�]��@�����ٿ��A�Nn�@����3@9�z^O�!?t�F�]��@�����ٿ��A�Nn�@����3@9�z^O�!?t�F�]��@Ӟ�VO�ٿⓝ��a�@��w��3@8��(�!?�հ	���@Ӟ�VO�ٿⓝ��a�@��w��3@8��(�!?�հ	���@Ӟ�VO�ٿⓝ��a�@��w��3@8��(�!?�հ	���@Ӟ�VO�ٿⓝ��a�@��w��3@8��(�!?�հ	���@Ӟ�VO�ٿⓝ��a�@��w��3@8��(�!?�հ	���@P����ٿ�q��@��+6b�3@8��V�!?�U ����@P����ٿ�q��@��+6b�3@8��V�!?�U ����@P����ٿ�q��@��+6b�3@8��V�!?�U ����@P����ٿ�q��@��+6b�3@8��V�!?�U ����@P����ٿ�q��@��+6b�3@8��V�!?�U ����@{'�Břٿ{�k�W�@�Ŗ��3@X�}�!?Ѳ:�� �@{'�Břٿ{�k�W�@�Ŗ��3@X�}�!?Ѳ:�� �@���+�ٿ�D/�.�@K���v�3@`h�|�!?�W�q�{�@�1_��ٿC���@�iہ!�3@H����!?���\H��@�1_��ٿC���@�iہ!�3@H����!?���\H��@�1_��ٿC���@�iہ!�3@H����!?���\H��@�1_��ٿC���@�iہ!�3@H����!?���\H��@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@ͺ8Hܖٿ���rY��@D
�I�3@�/��j�!?̽��b�@<��ٿZO�y|�@u��f	�3@����F�!?8�x�@���ᦔٿ:P)�/�@K�יK�3@�����!?m�QP�2�@���ᦔٿ:P)�/�@K�יK�3@�����!?m�QP�2�@���ᦔٿ:P)�/�@K�יK�3@�����!?m�QP�2�@���ᦔٿ:P)�/�@K�יK�3@�����!?m�QP�2�@�)jV�ٿ�^v_��@�G�j�3@9a,J�!?�E�ӻ�@�)jV�ٿ�^v_��@�G�j�3@9a,J�!?�E�ӻ�@�)jV�ٿ�^v_��@�G�j�3@9a,J�!?�E�ӻ�@�)jV�ٿ�^v_��@�G�j�3@9a,J�!?�E�ӻ�@��F�ٿ)��5��@��
4@�%�m�!?�ЭzK{�@��F�ٿ)��5��@��
4@�%�m�!?�ЭzK{�@v�o��ٿI��T�@m�� ��3@8Y��!?��h�9�@v�o��ٿI��T�@m�� ��3@8Y��!?��h�9�@���ٿ4���<m�@��n��3@I����!?������@�;>���ٿ^kiߡd�@&�v!�3@�$�?��!?/��,/~�@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ٿ�]uN\��@��ϻ�3@�����!?�����@���ޔٿ��B���@��4~�3@�/yR�!?푟���@&��7��ٿ���yz��@%j��Z�3@�3��!�!?�"���<�@&��7��ٿ���yz��@%j��Z�3@�3��!�!?�"���<�@�?�? �ٿ#	)Ek�@�=]u�4@���� �!?�|̞��@�?�? �ٿ#	)Ek�@�=]u�4@���� �!?�|̞��@�?�? �ٿ#	)Ek�@�=]u�4@���� �!?�|̞��@�?�? �ٿ#	)Ek�@�=]u�4@���� �!?�|̞��@�F��D�ٿ_��Y�@/L���3@!����!?����@�F��D�ٿ_��Y�@/L���3@!����!?����@�ȁ�ٿ�;S!Tl�@X�Co��3@G9#J�!?I��А�@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@�w]Q�ٿXW�����@��?��3@S��J\�!?=����@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@'�A}��ٿ��?���@�ڗ��3@��i�;�!?��X­w�@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@ڐ �ݓٿ�(f��m�@�Cx���3@&�]"&�!?�d%p��@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@�5�Y�ٿ������@��g_�3@�YO/�!?��N�Xx�@E�f�c�ٿ�m\I�	�@��'��3@��xD-�!?�+��ڴ@E�f�c�ٿ�m\I�	�@��'��3@��xD-�!?�+��ڴ@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@OJ%A��ٿ�Rq���@��>Co�3@�s�i{�!?�g"��0�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@)H�-�ٿ	����@��Z�D�3@MXa+t�!?��(�"
�@�y�ژٿ}@@ʱ�@{�C�o�3@���!?�����(�@�y�ژٿ}@@ʱ�@{�C�o�3@���!?�����(�@�y�ژٿ}@@ʱ�@{�C�o�3@���!?�����(�@�y�ژٿ}@@ʱ�@{�C�o�3@���!?�����(�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@�v���ٿ߼��~:�@�q";�3@^�x�^�!?�Q#.R�@��h뗑ٿs{L���@�
����3@��V_�!?�O}��@��h뗑ٿs{L���@�
����3@��V_�!?�O}��@>�=���ٿlx�G���@E����3@}x����!?�!�ñ�@>�=���ٿlx�G���@E����3@}x����!?�!�ñ�@>�=���ٿlx�G���@E����3@}x����!?�!�ñ�@>�=���ٿlx�G���@E����3@}x����!?�!�ñ�@f�z�i�ٿ���\���@e4�3��3@dHd.��!?|����@,seLB�ٿ�����=�@8��<8�3@'E�F�!?��C�ڴ@,seLB�ٿ�����=�@8��<8�3@'E�F�!?��C�ڴ@,seLB�ٿ�����=�@8��<8�3@'E�F�!?��C�ڴ@wyw��ٿǫ��ο@h12+�3@ADa�>�!?u㨟�\�@wyw��ٿǫ��ο@h12+�3@ADa�>�!?u㨟�\�@wyw��ٿǫ��ο@h12+�3@ADa�>�!?u㨟�\�@wyw��ٿǫ��ο@h12+�3@ADa�>�!?u㨟�\�@wyw��ٿǫ��ο@h12+�3@ADa�>�!?u㨟�\�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@�~���ٿ��2D)��@
�0���3@_�ЍP�!?�:]�nP�@���ٿN�`��@�}،�3@򎽊�!?�٢Fs�@�^��ٿ~V�V���@�<YPg�3@����E�!?�/�nd�@�^��ٿ~V�V���@�<YPg�3@����E�!?�/�nd�@]���ٿ�8��3.�@����3@D&�2�!?���Fs�@��u��ٿ-�	�PU�@
��n��3@R�Fz!�!?;��P���@��u��ٿ-�	�PU�@
��n��3@R�Fz!�!?;��P���@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@�;�\��ٿ�w��}��@���3@��Ǜ;�!?�_3��R�@+O�+֚ٿ	��n��@ͼ��3@��w\�!?��3� �@+O�+֚ٿ	��n��@ͼ��3@��w\�!?��3� �@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@�E�I=�ٿ67����@�*j�3@�y�ϳ�!?~�G��@ʩ�ٿ�����@�Iu�G�3@�oI!?�[�_t�@ʩ�ٿ�����@�Iu�G�3@�oI!?�[�_t�@B�����ٿ�n�{U��@��0���3@dzd�_�!?.$T<~�@B�����ٿ�n�{U��@��0���3@dzd�_�!?.$T<~�@B�����ٿ�n�{U��@��0���3@dzd�_�!?.$T<~�@B�����ٿ�n�{U��@��0���3@dzd�_�!?.$T<~�@B�����ٿ�n�{U��@��0���3@dzd�_�!?.$T<~�@;���ٿ���\��@�΢���3@JC�0�!?��.��/�@������ٿWl��n�@.SE��3@)';�M�!?��
��Ҵ@������ٿWl��n�@.SE��3@)';�M�!?��
��Ҵ@������ٿWl��n�@.SE��3@)';�M�!?��
��Ҵ@������ٿWl��n�@.SE��3@)';�M�!?��
��Ҵ@������ٿWl��n�@.SE��3@)';�M�!?��
��Ҵ@fu�_�ٿ�iT3S��@���+�3@.���|�!?3"U
ܽ�@�Z;��ٿ�ɊLml�@�����3@�Z�"!�!?��1�wӴ@�Z;��ٿ�ɊLml�@�����3@�Z�"!�!?��1�wӴ@�Z;��ٿ�ɊLml�@�����3@�Z�"!�!?��1�wӴ@�z��s�ٿ��텫��@}�kޝ�3@!tQJG�!?��+�ɵ@�z��s�ٿ��텫��@}�kޝ�3@!tQJG�!?��+�ɵ@�|49��ٿm���0V�@�{§�3@.}�sk�!?p�����@�|49��ٿm���0V�@�{§�3@.}�sk�!?p�����@�|49��ٿm���0V�@�{§�3@.}�sk�!?p�����@�|49��ٿm���0V�@�{§�3@.}�sk�!?p�����@�|49��ٿm���0V�@�{§�3@.}�sk�!?p�����@��ꃞٿ$�Q�w��@�����3@o�~�!?r1D_�;�@��ꃞٿ$�Q�w��@�����3@o�~�!?r1D_�;�@��ꃞٿ$�Q�w��@�����3@o�~�!?r1D_�;�@�h|'��ٿC�v�@���v��3@lv�k�!?���.ߴ@�h|'��ٿC�v�@���v��3@lv�k�!?���.ߴ@�h|'��ٿC�v�@���v��3@lv�k�!?���.ߴ@�h|'��ٿC�v�@���v��3@lv�k�!?���.ߴ@�h|'��ٿC�v�@���v��3@lv�k�!?���.ߴ@$_�Y�ٿuݪ�}��@��t[�3@��_�!?�,F�д@$_�Y�ٿuݪ�}��@��t[�3@��_�!?�,F�д@$_�Y�ٿuݪ�}��@��t[�3@��_�!?�,F�д@�e6}��ٿy.tQ�@+mQ�3@{���$�!?�0rsK��@�e6}��ٿy.tQ�@+mQ�3@{���$�!?�0rsK��@�e6}��ٿy.tQ�@+mQ�3@{���$�!?�0rsK��@�e6}��ٿy.tQ�@+mQ�3@{���$�!?�0rsK��@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@��	菔ٿ*�VE
�@�oR6�3@�3�x�!?��4� �@ffg���ٿ���(�@R��5�3@�=�|F�!?s�'Y�&�@ffg���ٿ���(�@R��5�3@�=�|F�!?s�'Y�&�@ffg���ٿ���(�@R��5�3@�=�|F�!?s�'Y�&�@ffg���ٿ���(�@R��5�3@�=�|F�!?s�'Y�&�@ffg���ٿ���(�@R��5�3@�=�|F�!?s�'Y�&�@@\�ܙ�ٿ4 ���@�M���3@�z�9]�!?m�dw��@U�6!��ٿ�]���R�@z��d�3@]��)�!?/��ߺϴ@U�6!��ٿ�]���R�@z��d�3@]��)�!?/��ߺϴ@U�6!��ٿ�]���R�@z��d�3@]��)�!?/��ߺϴ@U�6!��ٿ�]���R�@z��d�3@]��)�!?/��ߺϴ@U�6!��ٿ�]���R�@z��d�3@]��)�!?/��ߺϴ@����ٿk�#��@a����3@!���$�!?R�aú�@����ٿk�#��@a����3@!���$�!?R�aú�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@Y��?��ٿ$4����@y�(]��3@'˩�D�!?�CE;�@2���ٿWԒJ��@��M�3@���/�!?�	F=�@2���ٿWԒJ��@��M�3@���/�!?�	F=�@2���ٿWԒJ��@��M�3@���/�!?�	F=�@�&��:�ٿ���L���@�����3@
�9�6�!?Cu��zڵ@�y���ٿ-��$��@�ű���3@���Ŏ�!?�I�Ƶ@�y���ٿ-��$��@�ű���3@���Ŏ�!?�I�Ƶ@Z>�H~�ٿ����@����B4@ҩ��b�!?K�Dp�t�@Z>�H~�ٿ����@����B4@ҩ��b�!?K�Dp�t�@Z>�H~�ٿ����@����B4@ҩ��b�!?K�Dp�t�@Z>�H~�ٿ����@����B4@ҩ��b�!?K�Dp�t�@Z>�H~�ٿ����@����B4@ҩ��b�!?K�Dp�t�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@�h+��ٿ�%�@���@�5�4@�A .t�!?f�f/�@&Tn.�ٿ����S��@!EBY�	4@��`Da�!?�1..�@&Tn.�ٿ����S��@!EBY�	4@��`Da�!?�1..�@&Tn.�ٿ����S��@!EBY�	4@��`Da�!?�1..�@�X��ٿ�y-k�@�3(��3@�"nt�!?ɞ���@�X��ٿ�y-k�@�3(��3@�"nt�!?ɞ���@�X��ٿ�y-k�@�3(��3@�"nt�!?ɞ���@�X��ٿ�y-k�@�3(��3@�"nt�!?ɞ���@�u��ٿ��i`S|�@�$�v:�3@�W'e�!?�]��v��@D`���ٿ���f_I�@�U�74@% �J�!?w-�2��@D`���ٿ���f_I�@�U�74@% �J�!?w-�2��@��D��ٿh&�?�@B|M��4@(�-�Y�!?�|���R�@��D��ٿh&�?�@B|M��4@(�-�Y�!?�|���R�@��D��ٿh&�?�@B|M��4@(�-�Y�!?�|���R�@!�逯�ٿ���2p�@�K�R�3@/"[Ň�!?m�lN��@!�逯�ٿ���2p�@�K�R�3@/"[Ň�!?m�lN��@!�逯�ٿ���2p�@�K�R�3@/"[Ň�!?m�lN��@	�ٙٿ�,���@B��ڐ�3@�}��^�!?������@	�ٙٿ�,���@B��ڐ�3@�}��^�!?������@ځ�
��ٿ�پjcJ�@Q-Y�3@��{a�!?*8;��Ѵ@ځ�
��ٿ�پjcJ�@Q-Y�3@��{a�!?*8;��Ѵ@ځ�
��ٿ�پjcJ�@Q-Y�3@��{a�!?*8;��Ѵ@ځ�
��ٿ�پjcJ�@Q-Y�3@��{a�!?*8;��Ѵ@���掕ٿ��@"O�@��fA��3@�=)�9�!?)�$��@���掕ٿ��@"O�@��fA��3@�=)�9�!?)�$��@:��(٘ٿ@*�H0�@���N�3@LitU�!?�I5���@:��(٘ٿ@*�H0�@���N�3@LitU�!?�I5���@:��(٘ٿ@*�H0�@���N�3@LitU�!?�I5���@:��(٘ٿ@*�H0�@���N�3@LitU�!?�I5���@:��(٘ٿ@*�H0�@���N�3@LitU�!?�I5���@�c���ٿ!6�.}�@�'���3@��mWk�!?qy���@�c���ٿ!6�.}�@�'���3@��mWk�!?qy���@d�,1I�ٿ�x�����@5��]%�3@;s�0H�!?aM��G��@d�,1I�ٿ�x�����@5��]%�3@;s�0H�!?aM��G��@d�,1I�ٿ�x�����@5��]%�3@;s�0H�!?aM��G��@OӋ��ٿ#�V�:�@�!� 4@�*�-7�!?>ʏ�s�@OӋ��ٿ#�V�:�@�!� 4@�*�-7�!?>ʏ�s�@)y�fu�ٿ@��F[6�@����k�3@��ff<�!?l�>�h��@)y�fu�ٿ@��F[6�@����k�3@��ff<�!?l�>�h��@)y�fu�ٿ@��F[6�@����k�3@��ff<�!?l�>�h��@"r(��ٿ��+P=[�@�枚64@����!?�R#j�@"r(��ٿ��+P=[�@�枚64@����!?�R#j�@��Ȑٿ���
=�@�#�Pg4@���ZG�!?Cþ#�@��Ȑٿ���
=�@�#�Pg4@���ZG�!?Cþ#�@��Ȑٿ���
=�@�#�Pg4@���ZG�!?Cþ#�@��Ȑٿ���
=�@�#�Pg4@���ZG�!?Cþ#�@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@�?�΢�ٿ1(͌�"�@@�Y�.�3@� /�A�!?}�c����@%��V�ٿ<e��W�@?����3@뻣�f�!?]rs_�@%��V�ٿ<e��W�@?����3@뻣�f�!?]rs_�@%��V�ٿ<e��W�@?����3@뻣�f�!?]rs_�@%��V�ٿ<e��W�@?����3@뻣�f�!?]rs_�@%��V�ٿ<e��W�@?����3@뻣�f�!?]rs_�@��
��ٿ��Ȋ�@ℌpg�3@+���k�!?z���lQ�@��
��ٿ��Ȋ�@ℌpg�3@+���k�!?z���lQ�@��
��ٿ��Ȋ�@ℌpg�3@+���k�!?z���lQ�@��
��ٿ��Ȋ�@ℌpg�3@+���k�!?z���lQ�@�)d/P�ٿ6�F6O��@�[�,�3@U�W )�!?�2�i�@�)d/P�ٿ6�F6O��@�[�,�3@U�W )�!?�2�i�@�)d/P�ٿ6�F6O��@�[�,�3@U�W )�!?�2�i�@�}���ٿ�;�y[w�@v#a��3@��g��!?+��>�@�}���ٿ�;�y[w�@v#a��3@��g��!?+��>�@�}���ٿ�;�y[w�@v#a��3@��g��!?+��>�@�2881�ٿ8� ù��@�&���3@ܸ�`�!?n�Õ۴@�2881�ٿ8� ù��@�&���3@ܸ�`�!?n�Õ۴@�2881�ٿ8� ù��@�&���3@ܸ�`�!?n�Õ۴@�2881�ٿ8� ù��@�&���3@ܸ�`�!?n�Õ۴@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@���j��ٿ�l���2�@*)+���3@4:o=�!?��p���@����ٿ���Y)�@9��Ѱ�3@O��Y`�!?l;D=��@����ٿ���Y)�@9��Ѱ�3@O��Y`�!?l;D=��@����ٿ���Y)�@9��Ѱ�3@O��Y`�!?l;D=��@ʮݦ��ٿ*^���B�@8��)c�3@��Xs�!?A��ㄊ�@}CMt7�ٿ6d[NX�@j�R�L4@`v�~��!?����`�@}CMt7�ٿ6d[NX�@j�R�L4@`v�~��!?����`�@�E�).�ٿY�Mq���@�D�P>4@��y���!?��Z�Z��@(O�&��ٿ��Vh��@�<�4@C8��!?8+�LHR�@(O�&��ٿ��Vh��@�<�4@C8��!?8+�LHR�@(O�&��ٿ��Vh��@�<�4@C8��!?8+�LHR�@�;߱��ٿ>AWlK�@�lE4@ؿ.�k�!?��W
�H�@�;߱��ٿ>AWlK�@�lE4@ؿ.�k�!?��W
�H�@�;߱��ٿ>AWlK�@�lE4@ؿ.�k�!?��W
�H�@N�Z�ٿ���I��@������3@-�
��!?��&&ܴ@Ƣ���ٿӞ�i��@.B��3@ W���!?M���5�@Ƣ���ٿӞ�i��@.B��3@ W���!?M���5�@,N��f�ٿ.�K�Y�@[y����3@��ᤁ�!?X�խ[�@,N��f�ٿ.�K�Y�@[y����3@��ᤁ�!?X�խ[�@,N��f�ٿ.�K�Y�@[y����3@��ᤁ�!?X�խ[�@K��{�ٿE�f_�G�@&�#��3@��
Ӑ!?�:>�@K��{�ٿE�f_�G�@&�#��3@��
Ӑ!?�:>�@N�"��ٿ?�o��R�@���b��3@�O͐!?���ڴ@N�"��ٿ?�o��R�@���b��3@�O͐!?���ڴ@�g�߶�ٿ
�����@���>m�3@j���А!?/�o��l�@�g�߶�ٿ
�����@���>m�3@j���А!?/�o��l�@�g�߶�ٿ
�����@���>m�3@j���А!?/�o��l�@�g�߶�ٿ
�����@���>m�3@j���А!?/�o��l�@��f���ٿ������@Ԋ��3@���!?����|�@��f���ٿ������@Ԋ��3@���!?����|�@��f���ٿ������@Ԋ��3@���!?����|�@K�Q��ٿ�t��%G�@.E.�3@>}�֞�!?�����@K�Q��ٿ�t��%G�@.E.�3@>}�֞�!?�����@K�Q��ٿ�t��%G�@.E.�3@>}�֞�!?�����@K�Q��ٿ�t��%G�@.E.�3@>}�֞�!?�����@K�Q��ٿ�t��%G�@.E.�3@>}�֞�!?�����@�:�A�ٿ��[�K�@ǐ���3@8�Ow�!?e�l1��@�:�A�ٿ��[�K�@ǐ���3@8�Ow�!?e�l1��@�i\�j�ٿ��g���@�64K��3@��U��!?��1׭�@�i\�j�ٿ��g���@�64K��3@��U��!?��1׭�@�i\�j�ٿ��g���@�64K��3@��U��!?��1׭�@W;�z;�ٿ�� ��@� ����3@o#Ab��!?I�RP��@��&��ٿ�Z��)��@m�14@]rj�v�!?���6�@��&��ٿ�Z��)��@m�14@]rj�v�!?���6�@��&��ٿ�Z��)��@m�14@]rj�v�!?���6�@��&��ٿ�Z��)��@m�14@]rj�v�!?���6�@X�Q:ٿ��k�j��@>��74@Z*�&��!?6o��*�@X�Q:ٿ��k�j��@>��74@Z*�&��!?6o��*�@X�Q:ٿ��k�j��@>��74@Z*�&��!?6o��*�@X�Q:ٿ��k�j��@>��74@Z*�&��!?6o��*�@X�Q:ٿ��k�j��@>��74@Z*�&��!?6o��*�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@Ԩ�h�ٿ���[
M�@��o�3@]1%���!?<�F�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@���ٿ��J���@�Eʬ��3@^hz&�!?�|�C�@~�7j�ٿH���m>�@��a%�3@�p!�4�!?&�Oc]�@~�7j�ٿH���m>�@��a%�3@�p!�4�!?&�Oc]�@�CU:B�ٿ�,��@���xx�3@x:J��!?��c���@�CU:B�ٿ�,��@���xx�3@x:J��!?��c���@�CU:B�ٿ�,��@���xx�3@x:J��!?��c���@T��U�ٿ}�Dg
��@xٹ��3@W�� �!?3���DԴ@T��U�ٿ}�Dg
��@xٹ��3@W�� �!?3���DԴ@T��U�ٿ}�Dg
��@xٹ��3@W�� �!?3���DԴ@T��U�ٿ}�Dg
��@xٹ��3@W�� �!?3���DԴ@T��U�ٿ}�Dg
��@xٹ��3@W�� �!?3���DԴ@�u�}�ٿq�N�(B�@k�$O4�3@ކG�я!? �@�M(�@�u�}�ٿq�N�(B�@k�$O4�3@ކG�я!? �@�M(�@�Gb��ٿ+5͈�@?2*�3@����5�!?5�Np�@�Gb��ٿ+5͈�@?2*�3@����5�!?5�Np�@�Gb��ٿ+5͈�@?2*�3@����5�!?5�Np�@�Gb��ٿ+5͈�@?2*�3@����5�!?5�Np�@2���d�ٿ�ڴ��S�@`v�5�3@�vN�!? ��V�ϴ@2���d�ٿ�ڴ��S�@`v�5�3@�vN�!? ��V�ϴ@2���d�ٿ�ڴ��S�@`v�5�3@�vN�!? ��V�ϴ@��'M�ٿ���y��@�ϸ�G�3@����V�!?�ԳK5�@��'M�ٿ���y��@�ϸ�G�3@����V�!?�ԳK5�@��'M�ٿ���y��@�ϸ�G�3@����V�!?�ԳK5�@��'M�ٿ���y��@�ϸ�G�3@����V�!?�ԳK5�@��'M�ٿ���y��@�ϸ�G�3@����V�!?�ԳK5�@j�=D/�ٿ؜�����@�b*�4@�	��+�!?y�oE_�@j�=D/�ٿ؜�����@�b*�4@�	��+�!?y�oE_�@h�^���ٿ��oia�@�&@���3@�cx�[�!?�~9]<i�@h�^���ٿ��oia�@�&@���3@�cx�[�!?�~9]<i�@h�^���ٿ��oia�@�&@���3@�cx�[�!?�~9]<i�@h�^���ٿ��oia�@�&@���3@�cx�[�!?�~9]<i�@h�^���ٿ��oia�@�&@���3@�cx�[�!?�~9]<i�@�+�e�ٿp�A̞b�@�,��4@E�h�'�!?���nk�@�+�e�ٿp�A̞b�@�,��4@E�h�'�!?���nk�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�M�az�ٿ�������@�M����3@���%�!?Y��L[�@�fXk�ٿ4�1+��@���C�4@�{��@�!?��r.h��@�fXk�ٿ4�1+��@���C�4@�{��@�!?��r.h��@�fXk�ٿ4�1+��@���C�4@�{��@�!?��r.h��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@4�z��ٿ���!���@�)���3@*�6�!?�$��@ [�(בٿe͑����@��r���3@�f=�!?�����B�@ [�(בٿe͑����@��r���3@�f=�!?�����B�@6GS$�ٿa����@p����3@0�I*�!?���h�@6GS$�ٿa����@p����3@0�I*�!?���h�@��A-�ٿ<i�8��@����4@���2�!?8p��z��@��qu�ٿ*?�v���@�yO�:�3@���I؏!?[]�RU;�@��qu�ٿ*?�v���@�yO�:�3@���I؏!?[]�RU;�@��qu�ٿ*?�v���@�yO�:�3@���I؏!?[]�RU;�@��qu�ٿ*?�v���@�yO�:�3@���I؏!?[]�RU;�@}j�h9�ٿXy�R��@�޸��3@>�9P9�!?��״@}j�h9�ٿXy�R��@�޸��3@>�9P9�!?��״@#�}��ٿ�����@���Q�3@s=5�P�!?v$+^���@#�}��ٿ�����@���Q�3@s=5�P�!?v$+^���@#�}��ٿ�����@���Q�3@s=5�P�!?v$+^���@=���ٿ�[��@j���'�3@+�}�f�!?��!&���@=���ٿ�[��@j���'�3@+�}�f�!?��!&���@=���ٿ�[��@j���'�3@+�}�f�!?��!&���@�p�זٿy���W�@4A��3@���G�!?� 0��!�@�p�זٿy���W�@4A��3@���G�!?� 0��!�@�p�זٿy���W�@4A��3@���G�!?� 0��!�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@6�=�7�ٿcE`��@�s�4@#��/�!?��եqb�@�7���ٿ'4�;�1�@�j��5�3@�c䞗�!?�� ����@�7���ٿ'4�;�1�@�j��5�3@�c䞗�!?�� ����@�7���ٿ'4�;�1�@�j��5�3@�c䞗�!?�� ����@�7���ٿ'4�;�1�@�j��5�3@�c䞗�!?�� ����@�7���ٿ'4�;�1�@�j��5�3@�c䞗�!?�� ����@X�eс�ٿ��'v���@�Km�J�3@�V	�!?;eK����@X�eс�ٿ��'v���@�Km�J�3@�V	�!?;eK����@X�eс�ٿ��'v���@�Km�J�3@�V	�!?;eK����@�k˳1�ٿ`ĺg��@���D�4@��u���!?�N(��@�k˳1�ٿ`ĺg��@���D�4@��u���!?�N(��@�k˳1�ٿ`ĺg��@���D�4@��u���!?�N(��@='��ٿ��v@p��@����3@�{�ZI�!?�2�6�ô@='��ٿ��v@p��@����3@�{�ZI�!?�2�6�ô@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@
c�n�ٿ!�k�L�@�]8��3@�&��+�!?�أ��@_̜���ٿ�d�����@�#Uy�3@39��!?�eb�q�@_̜���ٿ�d�����@�#Uy�3@39��!?�eb�q�@����ٿ�˪�K��@��G��3@�^ᅏ!?�9�D�@����ٿ�˪�K��@��G��3@�^ᅏ!?�9�D�@pK��ٿT���(�@�����3@C��L�!?��h�խ�@f+�]�ٿ�gys��@�0�7��3@�B�!?ơ/��1�@f+�]�ٿ�gys��@�0�7��3@�B�!?ơ/��1�@f+�]�ٿ�gys��@�0�7��3@�B�!?ơ/��1�@f+�]�ٿ�gys��@�0�7��3@�B�!?ơ/��1�@k�PZ�ٿ[�㒊�@��<6�3@�>�J3�!?w�$�\�@k�PZ�ٿ[�㒊�@��<6�3@�>�J3�!?w�$�\�@k�PZ�ٿ[�㒊�@��<6�3@�>�J3�!?w�$�\�@k�PZ�ٿ[�㒊�@��<6�3@�>�J3�!?w�$�\�@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@@�°��ٿ�&�1���@�A���3@`�{s�!? ɇ��ߴ@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@�Z�S��ٿ��e�@:��l�3@�Bx[�!?h�M���@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@bBf�g�ٿ�·���@<���2�3@2P��-�!?J�V	�Y�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@1�s���ٿ��Vk��@ҧ)�3@Vb�q�!?�X�:�@	»��ٿ��o���@�#���3@L!?��?��-�@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@�n���ٿm}� E�@D79�4@R�?R�!?�3|Nٴ@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����[�ٿEվ2:�@�����3@�ۯbQ�!?)~V���@����ΔٿI�����@��e5��3@�Rǃ3�!?Ez��2�@����ΔٿI�����@��e5��3@�Rǃ3�!?Ez��2�@����ΔٿI�����@��e5��3@�Rǃ3�!?Ez��2�@����ΔٿI�����@��e5��3@�Rǃ3�!?Ez��2�@����ΔٿI�����@��e5��3@�Rǃ3�!?Ez��2�@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@��hٙٿ���(T�@t,K��3@����!?�If�2��@�
��X�ٿ
}�-���@��_F��3@����7�!?ګ& !�@�
��X�ٿ
}�-���@��_F��3@����7�!?ګ& !�@KL9�ٿ�Q:����@� 4c�3@����D�!?�pG��@KL9�ٿ�Q:����@� 4c�3@����D�!?�pG��@KL9�ٿ�Q:����@� 4c�3@����D�!?�pG��@KL9�ٿ�Q:����@� 4c�3@����D�!?�pG��@=�]�˗ٿ�V�7�p�@ԫ��3@�Vw�!?��a�(P�@�̉B��ٿ��P:Ҿ�@[��t��3@�y�p#�!?/��Was�@�̉B��ٿ��P:Ҿ�@[��t��3@�y�p#�!?/��Was�@�̉B��ٿ��P:Ҿ�@[��t��3@�y�p#�!?/��Was�@�̉B��ٿ��P:Ҿ�@[��t��3@�y�p#�!?/��Was�@��ߒx�ٿg���p��@��w�3@;\k�'�!?��"�%J�@t��[c�ٿXx��{�@㬈2u�3@�G��!�!?���d6�@t��[c�ٿXx��{�@㬈2u�3@�G��!�!?���d6�@t��[c�ٿXx��{�@㬈2u�3@�G��!�!?���d6�@t��[c�ٿXx��{�@㬈2u�3@�G��!�!?���d6�@��4���ٿB�E�ӳ�@�����3@��1��!?v3�&Ǵ@�+Y��ٿ;Y�=ڨ�@fB��/�3@6u<N�!?�ś/x��@)���ٿn����@@����3@(�.�!?W�dR�@)���ٿn����@@����3@(�.�!?W�dR�@)���ٿn����@@����3@(�.�!?W�dR�@)���ٿn����@@����3@(�.�!?W�dR�@)���ٿn����@@����3@(�.�!?W�dR�@)���ٿn����@@����3@(�.�!?W�dR�@31���ٿN�vn��@'��x0�3@�^oX�!?�2��l��@Q9M%��ٿ�dH���@6�+��3@���w�!?�:5�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@��փ=�ٿ��)����@�?b�3@�����!?��J��4�@@=>��ٿl���p�@�-�d��3@�骹��!?%���+�@@=>��ٿl���p�@�-�d��3@�骹��!?%���+�@@=>��ٿl���p�@�-�d��3@�骹��!?%���+�@@=>��ٿl���p�@�-�d��3@�骹��!?%���+�@@=>��ٿl���p�@�-�d��3@�骹��!?%���+�@z'�2�ٿ��$��@��Q��3@�<1Th�!?�8m����@z'�2�ٿ��$��@��Q��3@�<1Th�!?�8m����@z'�2�ٿ��$��@��Q��3@�<1Th�!?�8m����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@��V���ٿ7^���@�@D�^�#�3@����!?Z�����@ʰS��ٿ�^I���@Āg��3@v2�!?������@8	Sz$�ٿ1��3�@�����3@����!?��`�_j�@��a4�ٿO��#�j�@c��o�3@׋���!?���'��@���]M�ٿ4�^s�@J�T�3@Z��,�!?�RK�'�@���]M�ٿ4�^s�@J�T�3@Z��,�!?�RK�'�@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@7���ѕٿ�aܠp��@�ID��3@���M�!?>O��n��@GzPZ�ٿ�JN
��@��b��3@��
�[�!?ĤX��E�@e�O�J�ٿ���>��@~�`U�3@�4�fD�!?>>wb�@e�O�J�ٿ���>��@~�`U�3@�4�fD�!?>>wb�@e�O�J�ٿ���>��@~�`U�3@�4�fD�!?>>wb�@e�O�J�ٿ���>��@~�`U�3@�4�fD�!?>>wb�@�lc{ �ٿ4u�U�E�@��0���3@w|�_��!?X��6�	�@�lc{ �ٿ4u�U�E�@��0���3@w|�_��!?X��6�	�@b�I�u�ٿ�ȵ�t�@��j5��3@� _W�!?���'�@��?T�ٿ���%�@�b�vO�3@E\�X�!?�=ю���@��?T�ٿ���%�@�b�vO�3@E\�X�!?�=ю���@��?T�ٿ���%�@�b�vO�3@E\�X�!?�=ю���@5���F�ٿ�p�/���@`#ܘ�3@�
SH)�!?�$��Dִ@5���F�ٿ�p�/���@`#ܘ�3@�
SH)�!?�$��Dִ@5���F�ٿ�p�/���@`#ܘ�3@�
SH)�!?�$��Dִ@5���F�ٿ�p�/���@`#ܘ�3@�
SH)�!?�$��Dִ@�̦��ٿc����@��=T�3@.��R�!?����
�@�̦��ٿc����@��=T�3@.��R�!?����
�@�̦��ٿc����@��=T�3@.��R�!?����
�@�̦��ٿc����@��=T�3@.��R�!?����
�@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�<s�"�ٿɁ�~�@��E�G�3@�tHd}�!?4F�D�ϴ@�@i'�ٿ�hs�5�@����3@���p�!?��Иa.�@��(�ٿLsM�H�@����3@�P��!?+�=4�L�@��(�ٿLsM�H�@����3@�P��!?+�=4�L�@�����ٿ23�#)��@�����3@�����!?�cGRb��@�����ٿ23�#)��@�����3@�����!?�cGRb��@�����ٿ23�#)��@�����3@�����!?�cGRb��@�����ٿ23�#)��@�����3@�����!?�cGRb��@Z/9�ٿ>�]�@����3@�O]�!?%���@Z/9�ٿ>�]�@����3@�O]�!?%���@Z/9�ٿ>�]�@����3@�O]�!?%���@�C�P��ٿ��o5%�@'�6r4@/��J�!?�P3�}�@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@�#�Vv�ٿ�t~���@`X��3@��w�t�!?J�jq#��@܉p��ٿF �-A��@*O?� 4@�=`��!?<w�?M�@܉p��ٿF �-A��@*O?� 4@�=`��!?<w�?M�@܉p��ٿF �-A��@*O?� 4@�=`��!?<w�?M�@܉p��ٿF �-A��@*O?� 4@�=`��!?<w�?M�@܉p��ٿF �-A��@*O?� 4@�=`��!?<w�?M�@!�����ٿ1��O��@c/Y?��3@N��t��!?�Uh����@!�����ٿ1��O��@c/Y?��3@N��t��!?�Uh����@\����ٿ4�����@�S�"p�3@Ռ�5��!?@���Jߴ@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@�o�hΔٿ:o3��@u
	��3@5b҉��!?U{߼9�@^rp9��ٿ���	���@��&���3@�D����!?\8J�D?�@^rp9��ٿ���	���@��&���3@�D����!?\8J�D?�@^rp9��ٿ���	���@��&���3@�D����!?\8J�D?�@a���ٿw�%Yh_�@-�w�p�3@��6���!?���b-�@a���ٿw�%Yh_�@-�w�p�3@��6���!?���b-�@��7C�ٿ+]<�+�@��+�3@��Ϲ��!?��t�ʹ@��7C�ٿ+]<�+�@��+�3@��Ϲ��!?��t�ʹ@��7C�ٿ+]<�+�@��+�3@��Ϲ��!?��t�ʹ@��7C�ٿ+]<�+�@��+�3@��Ϲ��!?��t�ʹ@��7C�ٿ+]<�+�@��+�3@��Ϲ��!?��t�ʹ@p|����ٿ(���7�@��q��3@K�����!?���(��@p|����ٿ(���7�@��q��3@K�����!?���(��@p|����ٿ(���7�@��q��3@K�����!?���(��@^�ֱ �ٿ����O�@�
v,�3@�,��U�!?T+C2F<�@^�ֱ �ٿ����O�@�
v,�3@�,��U�!?T+C2F<�@^�ֱ �ٿ����O�@�
v,�3@�,��U�!?T+C2F<�@��s�͏ٿ��m�\��@`/�a��3@%�"�9�!?zt5��@��s�͏ٿ��m�\��@`/�a��3@%�"�9�!?zt5��@��$�H�ٿ�~���_�@��p��3@ii�ˇ�!?I�!�Qw�@��$�H�ٿ�~���_�@��p��3@ii�ˇ�!?I�!�Qw�@��$�H�ٿ�~���_�@��p��3@ii�ˇ�!?I�!�Qw�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@S��~�ٿY���@�@����3@l��G�!?��AN�S�@��h�G�ٿ��KDSs�@�+�H�3@�@4.��!?
9z"��@��h�G�ٿ��KDSs�@�+�H�3@�@4.��!?
9z"��@��h�G�ٿ��KDSs�@�+�H�3@�@4.��!?
9z"��@�`���ٿ�9\�_e�@G�9�{4@YF_�u�!?��52���@�`���ٿ�9\�_e�@G�9�{4@YF_�u�!?��52���@�`���ٿ�9\�_e�@G�9�{4@YF_�u�!?��52���@xDb#��ٿ�����ӿ@Fa4P�3@�����!?2a_ ��@xDb#��ٿ�����ӿ@Fa4P�3@�����!?2a_ ��@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@)N/"-�ٿK�}f'�@��H �3@k8��<�!?��򇵴@FO	c#�ٿ��%��@��� 4@\ZBv��!?��5�Ӿ�@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@Y3;�e�ٿɦS}���@i�F1�4@-��:o�!?�R5�{��@�o�1	�ٿ �����@8�!���3@V�j�l�!?Уv�@����_�ٿ Or���@P��k�4@Uq�I�!?��w���@ygl�7�ٿ�骒Fy�@M��h�3@:q�*�!?ke|i�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@�ס͜ٿ�'$��z�@�y]�3@ލ&�p�!?���H�G�@���݄�ٿi�����@��Q�8�3@h�3)�!?�~���@���݄�ٿi�����@��Q�8�3@h�3)�!?�~���@TgqΉ�ٿt]-��N�@*{��D4@�b^N�!?� `��@TgqΉ�ٿt]-��N�@*{��D4@�b^N�!?� `��@TgqΉ�ٿt]-��N�@*{��D4@�b^N�!?� `��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@�����ٿ��y4%�@X����3@��%ua�!?MBg��@K�dٖٿb��ˍ�@=5���3@���a�!?�(Cm��@�J�]�ٿr@甈��@���4�3@Z�93M�!?K���Ʈ�@L�t��ٿ�*�{cu�@�ʒo��3@h�t�d�!?��t�b��@L�t��ٿ�*�{cu�@�ʒo��3@h�t�d�!?��t�b��@L�t��ٿ�*�{cu�@�ʒo��3@h�t�d�!?��t�b��@L�t��ٿ�*�{cu�@�ʒo��3@h�t�d�!?��t�b��@L�t��ٿ�*�{cu�@�ʒo��3@h�t�d�!?��t�b��@��m�L�ٿ#ψ,���@�%*���3@c3��S�!?>����ε@��m�L�ٿ#ψ,���@�%*���3@c3��S�!?>����ε@��m�L�ٿ#ψ,���@�%*���3@c3��S�!?>����ε@��m�L�ٿ#ψ,���@�%*���3@c3��S�!?>����ε@��L��ٿzѳ���@��|&4@�0{�|�!?y>j,�ȴ@��L��ٿzѳ���@��|&4@�0{�|�!?y>j,�ȴ@��L��ٿzѳ���@��|&4@�0{�|�!?y>j,�ȴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@x��*�ٿ_�$)���@ �n�4@F�u�T�!?����ƴ@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�δh@�ٿ�H���@�S<h|�3@G���(�!?�nS���@�����ٿh��#���@�M+R��3@�x�H�!?�U8z��@�����ٿh��#���@�M+R��3@�x�H�!?�U8z��@�����ٿh��#���@�M+R��3@�x�H�!?�U8z��@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@Ђ�1�ٿ$Tu��O�@W�!<�4@��aM�!?�ٚE�%�@���'^�ٿ=p���1�@P��=4@���;�!?�������@���'^�ٿ=p���1�@P��=4@���;�!?�������@���'^�ٿ=p���1�@P��=4@���;�!?�������@��#g��ٿ��d�]�@���3@��\�s�!?���ʙY�@��#g��ٿ��d�]�@���3@��\�s�!?���ʙY�@\1�^�ٿ�Q�--~�@oJ4@�uc�V�!?f�m��9�@\1�^�ٿ�Q�--~�@oJ4@�uc�V�!?f�m��9�@\1�^�ٿ�Q�--~�@oJ4@�uc�V�!?f�m��9�@\1�^�ٿ�Q�--~�@oJ4@�uc�V�!?f�m��9�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@��/%�ٿ�������@�,����3@�]
 4�!?&�?�/�@�5Ii��ٿ�w����@�vl��3@�P�!"�!?R�!0#�@�5Ii��ٿ�w����@�vl��3@�P�!"�!?R�!0#�@6'�nȘٿ�n�N��@C�u�3@`uO�4�!?�:�頴@6'�nȘٿ�n�N��@C�u�3@`uO�4�!?�:�頴@�~}i^�ٿ�����@M���D�3@k���|�!?�����@�~}i^�ٿ�����@M���D�3@k���|�!?�����@�~}i^�ٿ�����@M���D�3@k���|�!?�����@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�T���ٿ̍;����@�-���3@p5��P�!?#�,���@�k�ٿ�v/Ҁ��@
��;�3@Et�?4�!?+��Gw��@�k�ٿ�v/Ҁ��@
��;�3@Et�?4�!?+��Gw��@�k�ٿ�v/Ҁ��@
��;�3@Et�?4�!?+��Gw��@�k�ٿ�v/Ҁ��@
��;�3@Et�?4�!?+��Gw��@��L�ٿ�<3�\�@�<�3@h�M2	�!?��IX�m�@��L�ٿ�<3�\�@�<�3@h�M2	�!?��IX�m�@��L�ٿ�<3�\�@�<�3@h�M2	�!?��IX�m�@��L�ٿ�<3�\�@�<�3@h�M2	�!?��IX�m�@��L�ٿ�<3�\�@�<�3@h�M2	�!?��IX�m�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�DO���ٿ�(��0`�@�"}�3@�ݰ�!?�j{d�@�0�ٿ�}}��@���/�3@}l�t.�!?}��4�a�@��
���ٿi�ۀj��@�@��3@��A�!?��g��@��
���ٿi�ۀj��@�@��3@��A�!?��g��@��
���ٿi�ۀj��@�@��3@��A�!?��g��@��
���ٿi�ۀj��@�@��3@��A�!?��g��@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@g�m��ٿ���&\�@�]q��3@+�D�T�!?��8z=�@Q�w�ٿ?����@���4@�}�(��!?$Ꙅ�@b�%O�ٿ�=¸���@h�!Ѵ4@˳\�!?>W|r��@b�%O�ٿ�=¸���@h�!Ѵ4@˳\�!?>W|r��@��n�&�ٿ3�m���@?b�Q]�3@�I�
�!?z�R��@��n�&�ٿ3�m���@?b�Q]�3@�I�
�!?z�R��@��n�&�ٿ3�m���@?b�Q]�3@�I�
�!?z�R��@��n�&�ٿ3�m���@?b�Q]�3@�I�
�!?z�R��@��n�&�ٿ3�m���@?b�Q]�3@�I�
�!?z�R��@7�ׁs�ٿ�X^���@˧�G�4@�mP$�!?�6RT���@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@j�Y��ٿ#I��u)�@'�{C:�3@�Y@��!?G������@�w�l�ٿDR�ro��@���4�3@#��!�!?��F]�@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@x+�䫗ٿ:�}g�@��kQp�3@JJh>�!?�V�6��@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@9p���ٿK{�)��@�q��3@]���!?_�H{ڋ�@�"P]��ٿ��,_�@F��k��3@O�~�!?S��ʭ�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@��2{G�ٿ����@o{�4C�3@D-�kΐ!?q<�/�%�@2�T (�ٿx�w�9�@�?��n4@��!?�V��e�@2�T (�ٿx�w�9�@�?��n4@��!?�V��e�@2�T (�ٿx�w�9�@�?��n4@��!?�V��e�@2�T (�ٿx�w�9�@�?��n4@��!?�V��e�@?ɖ�ٿ):�P/�@�����3@�uCP\�!?J�?Yx�@?ɖ�ٿ):�P/�@�����3@�uCP\�!?J�?Yx�@��˩��ٿ�C�#H�@�҉��3@u�f�!?J��W�@��˩��ٿ�C�#H�@�҉��3@u�f�!?J��W�@��˩��ٿ�C�#H�@�҉��3@u�f�!?J��W�@��˩��ٿ�C�#H�@�҉��3@u�f�!?J��W�@��˩��ٿ�C�#H�@�҉��3@u�f�!?J��W�@��0F�ٿհ ����@=�k���3@��!?��/�Ӵ@���}�ٿM �� �@�t.���3@�pC2�!?��12��@���}�ٿM �� �@�t.���3@�pC2�!?��12��@���}�ٿM �� �@�t.���3@�pC2�!?��12��@���}�ٿM �� �@�t.���3@�pC2�!?��12��@3�x�E�ٿ���u>�@��Bdx�3@��ku�!?�z>a�A�@3�x�E�ٿ���u>�@��Bdx�3@��ku�!?�z>a�A�@3�x�E�ٿ���u>�@��Bdx�3@��ku�!?�z>a�A�@3�x�E�ٿ���u>�@��Bdx�3@��ku�!?�z>a�A�@3�x�E�ٿ���u>�@��Bdx�3@��ku�!?�z>a�A�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@Z�O��ٿ/���y�@����3@r}�H��!??/s��~�@)y��ٿl�;�� �@L���3@��`��!?m���O�@)y��ٿl�;�� �@L���3@��`��!?m���O�@)y��ٿl�;�� �@L���3@��`��!?m���O�@)y��ٿl�;�� �@L���3@��`��!?m���O�@)y��ٿl�;�� �@L���3@��`��!?m���O�@)y��ٿl�;�� �@L���3@��`��!?m���O�@O�~��ٿُ���@U��p��3@B!fu�!?��L�?�@O�~��ٿُ���@U��p��3@B!fu�!?��L�?�@O�~��ٿُ���@U��p��3@B!fu�!?��L�?�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@2K_��ٿs!����@���5c�3@}j��!?����Z�@�n9�ٿ?��E��@.:�I�3@Q��KU�!?�{��/�@�n9�ٿ?��E��@.:�I�3@Q��KU�!?�{��/�@�n9�ٿ?��E��@.:�I�3@Q��KU�!?�{��/�@-ܸ�Y�ٿ&�qxL��@0��3t�3@�b=�=�!?§�pH�@-ܸ�Y�ٿ&�qxL��@0��3t�3@�b=�=�!?§�pH�@-ܸ�Y�ٿ&�qxL��@0��3t�3@�b=�=�!?§�pH�@-ܸ�Y�ٿ&�qxL��@0��3t�3@�b=�=�!?§�pH�@-ܸ�Y�ٿ&�qxL��@0��3t�3@�b=�=�!?§�pH�@��l��ٿg>�Ex�@'�H�*�3@_�9�u�!?L,�u��@��l��ٿg>�Ex�@'�H�*�3@_�9�u�!?L,�u��@g����ٿ��4c�'�@�; �o�3@A2L��!?��ꓺ�@g����ٿ��4c�'�@�; �o�3@A2L��!?��ꓺ�@���y��ٿHq���@W֐CE�3@R�,�i�!?�U0q�@���y��ٿHq���@W֐CE�3@R�,�i�!?�U0q�@7�]�ٿs�4v��@�w���3@k�p�U�!?����z�@7�]�ٿs�4v��@�w���3@k�p�U�!?����z�@FH����ٿw�����@��<Y��3@��rp~�!?7%Ѓ\��@|���֓ٿٮW���@�F)B�3@ބ0�/�!?�of����@|���֓ٿٮW���@�F)B�3@ބ0�/�!?�of����@|���֓ٿٮW���@�F)B�3@ބ0�/�!?�of����@|���֓ٿٮW���@�F)B�3@ބ0�/�!?�of����@|���֓ٿٮW���@�F)B�3@ބ0�/�!?�of����@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@�o��U�ٿ������@�d6��3@O�(U�!?�Ď��@V�b�ڒٿ��	���@L��!�3@�S�u�!?JW4�ڞ�@�
�H{�ٿ}�@���@-��x�3@|X� Ð!?0tǸ�O�@�
�H{�ٿ}�@���@-��x�3@|X� Ð!?0tǸ�O�@��d�ٿ��0/�@#��H�3@=�񒻐!?)�wi\�@��d�ٿ��0/�@#��H�3@=�񒻐!?)�wi\�@ö6�R�ٿEBkj��@�cӶ�3@��Y�H�!?x����y�@ö6�R�ٿEBkj��@�cӶ�3@��Y�H�!?x����y�@ö6�R�ٿEBkj��@�cӶ�3@��Y�H�!?x����y�@ö6�R�ٿEBkj��@�cӶ�3@��Y�H�!?x����y�@�-�e��ٿ�|�u��@vv@U��3@o��M�!?g��ߍ��@�_S�ٿbQ�yJ��@���Mf�3@E���>�!?��y4fp�@w���;�ٿ!�oC��@���3@�����!?t���s��@w���;�ٿ!�oC��@���3@�����!?t���s��@ߺj�}�ٿ��ҋo�@��w�4�3@�e^�!? ���I��@ߺj�}�ٿ��ҋo�@��w�4�3@�e^�!? ���I��@�Ǚ��ٿ}��4���@S4 .��3@s���!?����@A�Ugi�ٿ�J6�l��@�˾�H4@�_�
�!?�]���δ@A�Ugi�ٿ�J6�l��@�˾�H4@�_�
�!?�]���δ@A�Ugi�ٿ�J6�l��@�˾�H4@�_�
�!?�]���δ@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@���ٿ�<8���@Y�� $4@E�]pc�!?���ε@��8A^�ٿ�RB|C��@�Р+4@��gf(�!?�Y^�|�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@d�@�3�ٿ�U�l�2�@roU���3@9�o[:�!?��r�>�@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@��B�u�ٿ:�4e���@~�Gp��3@��:�!?�`B�)��@���N��ٿF_3ǚ��@��g��4@f����!?�P"��'�@��� 	�ٿ���!�@��ER4@����!?7��Ê�@��� 	�ٿ���!�@��ER4@����!?7��Ê�@��� 	�ٿ���!�@��ER4@����!?7��Ê�@��� 	�ٿ���!�@��ER4@����!?7��Ê�@��� 	�ٿ���!�@��ER4@����!?7��Ê�@x1J_�ٿs^��T�@˿s�S�3@L:���!?��?\� �@����ٿ�����@�$��3@����q�!?�bi�۵@��mi�ٿګ%�;��@�bR��3@Zza�M�!?�Z���@+��Y�ٿk+�H(��@4ϕ��3@��_d�!?)҄Q6�@+��Y�ٿk+�H(��@4ϕ��3@��_d�!?)҄Q6�@+��Y�ٿk+�H(��@4ϕ��3@��_d�!?)҄Q6�@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@����ٿ��eEO�@9R&��3@a%��Y�!?�(��n��@ÝM�+�ٿj�P���@�����3@^��_�!?��M��@ÝM�+�ٿj�P���@�����3@^��_�!?��M��@ÝM�+�ٿj�P���@�����3@^��_�!?��M��@ÝM�+�ٿj�P���@�����3@^��_�!?��M��@ÝM�+�ٿj�P���@�����3@^��_�!?��M��@�'I��ٿ�j�s��@nE�|P�3@��I�!?�tF,�@�'I��ٿ�j�s��@nE�|P�3@��I�!?�tF,�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@�՝�.�ٿ���N��@8�Z��3@q����!?��P�@b�� ��ٿ�DR���@Z��u�3@x��8a�!?�&�^�@b�� ��ٿ�DR���@Z��u�3@x��8a�!?�&�^�@b�� ��ٿ�DR���@Z��u�3@x��8a�!?�&�^�@�Wuw�ٿ��daR�@?�i!�3@��|�!?I�S1�@�Wuw�ٿ��daR�@?�i!�3@��|�!?I�S1�@�Wuw�ٿ��daR�@?�i!�3@��|�!?I�S1�@��8kߟٿ�K����@���q�3@�]<o�!?��77P�@��7.Q�ٿ2�7wnW�@��n��3@^��Z��!?�S���@��7.Q�ٿ2�7wnW�@��n��3@^��Z��!?�S���@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@[����ٿ?�fY��@��R��3@E(�#�!?���K g�@�]���ٿ���pG5�@�{_�8�3@m�C ��!?7��]�h�@�]���ٿ���pG5�@�{_�8�3@m�C ��!?7��]�h�@�]���ٿ���pG5�@�{_�8�3@m�C ��!?7��]�h�@�]���ٿ���pG5�@�{_�8�3@m�C ��!?7��]�h�@%�V�I�ٿj���W�@���>4�3@8ӤŲ�!?��w��o�@%�V�I�ٿj���W�@���>4�3@8ӤŲ�!?��w��o�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@���"�ٿ ���-��@�g��3@�+a��!?X�678K�@Q�F㯚ٿ�Y���@�W4��3@J�:q��!?�FY�ȵ@Q�F㯚ٿ�Y���@�W4��3@J�:q��!?�FY�ȵ@Q�F㯚ٿ�Y���@�W4��3@J�:q��!?�FY�ȵ@�MǐٿWR[:=U�@�C#c��3@��x͠�!?��(�!�@�MǐٿWR[:=U�@�C#c��3@��x͠�!?��(�!�@AK���ٿk�_���@V~���3@T��W�!?I��F�\�@AK���ٿk�_���@V~���3@T��W�!?I��F�\�@AK���ٿk�_���@V~���3@T��W�!?I��F�\�@AK���ٿk�_���@V~���3@T��W�!?I��F�\�@-�C�P�ٿl>S ���@T�����3@�D�a�!?�Ѯ��@-�C�P�ٿl>S ���@T�����3@�D�a�!?�Ѯ��@-�C�P�ٿl>S ���@T�����3@�D�a�!?�Ѯ��@-�C�P�ٿl>S ���@T�����3@�D�a�!?�Ѯ��@-�C�P�ٿl>S ���@T�����3@�D�a�!?�Ѯ��@,�C��ٿfG��x!�@/-���3@O���!?�����δ@�?�CӖٿL����@�U�x�3@Ѷ��!?<{=δ@;**Z�ٿ"���!��@�(�õ�3@p'\b��!?������@;**Z�ٿ"���!��@�(�õ�3@p'\b��!?������@;**Z�ٿ"���!��@�(�õ�3@p'\b��!?������@;**Z�ٿ"���!��@�(�õ�3@p'\b��!?������@;**Z�ٿ"���!��@�(�õ�3@p'\b��!?������@ۮ���ٿ$�r��@/��3@t���!?�L��Դ@ۮ���ٿ$�r��@/��3@t���!?�L��Դ@�C�H�ٿ�آ{��@q�d��3@=�����!?(@���״@�C�H�ٿ�آ{��@q�d��3@=�����!?(@���״@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@~Y*��ٿ:��Y��@�R��m4@o�ۅ�!?G'�^j�@^Ϣ+L�ٿÙ��'�@��e��3@~E���!?�����@^Ϣ+L�ٿÙ��'�@��e��3@~E���!?�����@^Ϣ+L�ٿÙ��'�@��e��3@~E���!?�����@^Ϣ+L�ٿÙ��'�@��e��3@~E���!?�����@^Ϣ+L�ٿÙ��'�@��e��3@~E���!?�����@�A���ٿ�|�n}h�@P��7��3@�9Wv�!?�B�클@�A���ٿ�|�n}h�@P��7��3@�9Wv�!?�B�클@�A���ٿ�|�n}h�@P��7��3@�9Wv�!?�B�클@�>.��ٿ�^ϡ�b�@���mf�3@1"�y�!?�Q$ hT�@�>.��ٿ�^ϡ�b�@���mf�3@1"�y�!?�Q$ hT�@׵t�~�ٿ���=/�@q�����3@��{H��!?�o��Z�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@w
턠ٿ���ι��@�s�X��3@צ0Fm�!?5%ǲ3!�@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@]�G�Ơٿ	�Usȳ�@@Ėt�3@<n,�2�!??����@&g��ٿ������@rƓC&�3@7?N�z�!?���O-�@&g��ٿ������@rƓC&�3@7?N�z�!?���O-�@&g��ٿ������@rƓC&�3@7?N�z�!?���O-�@&g��ٿ������@rƓC&�3@7?N�z�!?���O-�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@tץ� �ٿ�0>����@�%�Oo�3@��$*�!?�Z��;t�@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@�p�g�ٿJ����@��T���3@����g�!?�@eq��@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@TMxY��ٿ]�`���@�;�C�3@�b2�u�!?q����@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�`rg��ٿ֎�=/��@�8����3@�.�!?Ғ3N�U�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@�Ye'�ٿt@�X�@=xߍG�3@N���t�!?h+�J�@s�-�ٿ)���@X��T�3@�E�2�!?�=�cĴ@s�-�ٿ)���@X��T�3@�E�2�!?�=�cĴ@s�-�ٿ)���@X��T�3@�E�2�!?�=�cĴ@m_O��ٿ	��?��@:�����3@f��3�!?���a/�@m_O��ٿ	��?��@:�����3@f��3�!?���a/�@m_O��ٿ	��?��@:�����3@f��3�!?���a/�@m_O��ٿ	��?��@:�����3@f��3�!?���a/�@�6���ٿI"$��@��$�3@��J17�!?�(��'�@?��6
�ٿ "��@�����3@H�(E��!?�I���@sC��ٿ#Ǆ�.��@RT��3@퀽�l�!?��6h��@sC��ٿ#Ǆ�.��@RT��3@퀽�l�!?��6h��@6�
��ٿ*���@(�@�1���3@�=Q)�!?P�P�d��@6�
��ٿ*���@(�@�1���3@�=Q)�!?P�P�d��@6�
��ٿ*���@(�@�1���3@�=Q)�!?P�P�d��@6�
��ٿ*���@(�@�1���3@�=Q)�!?P�P�d��@{;g�I�ٿ�-�R��@�LJ6��3@��G|*�!?ii�Fs%�@{;g�I�ٿ�-�R��@�LJ6��3@��G|*�!?ii�Fs%�@{;g�I�ٿ�-�R��@�LJ6��3@��G|*�!?ii�Fs%�@�"/�S�ٿ��bI�u�@�3�!�3@b�ox�!?�^*R�@�"/�S�ٿ��bI�u�@�3�!�3@b�ox�!?�^*R�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@	�R$��ٿ#,"��o�@o��-��3@^�<�W�!?F��}�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@lRԚٿ�p=��H�@%V����3@nJh&�!?���'�@�hAO�ٿ�N*&�@p���6�3@��;b�!?K՜�x�@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@�+�G�ٿ��R����@l��3@�¥�9�!?�!~o��@T*��ٿع���@&)�>	�3@�~�%�!?0�K���@T*��ٿع���@&)�>	�3@�~�%�!?0�K���@dp{D�ٿP�r����@W���3@>Xt_�!?jUQ3V$�@dp{D�ٿP�r����@W���3@>Xt_�!?jUQ3V$�@dp{D�ٿP�r����@W���3@>Xt_�!?jUQ3V$�@dp{D�ٿP�r����@W���3@>Xt_�!?jUQ3V$�@dp{D�ٿP�r����@W���3@>Xt_�!?jUQ3V$�@		���ٿ�N��S�@�L=��3@\�;��!?��^m0�@		���ٿ�N��S�@�L=��3@\�;��!?��^m0�@		���ٿ�N��S�@�L=��3@\�;��!?��^m0�@B�W���ٿ#q�Q��@�����3@Ғ�0�!?����i�@B�W���ٿ#q�Q��@�����3@Ғ�0�!?����i�@B�W���ٿ#q�Q��@�����3@Ғ�0�!?����i�@B�W���ٿ#q�Q��@�����3@Ғ�0�!?����i�@ݢ\~j�ٿ�ս�J?�@���3@k�f�!?���ؚ�@��aB4�ٿJ*T���@����3@�Q���!?�6ڳ��@��aB4�ٿJ*T���@����3@�Q���!?�6ڳ��@��aB4�ٿJ*T���@����3@�Q���!?�6ڳ��@��aB4�ٿJ*T���@����3@�Q���!?�6ڳ��@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@�;���ٿ؊#?/�@�5�T;�3@R�1�E�!?�;_P�@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@��׷d�ٿFxL?z��@3?(���3@�U.p`�!?�+��1��@q��V�ٿ�t=�l�@�`��3@[=��L�!?�sH^�H�@q��V�ٿ�t=�l�@�`��3@[=��L�!?�sH^�H�@]w�/.�ٿ��,�R��@��P��3@i�Xt�!?���=�<�@q�).v�ٿ�=jM6�@��N�3@�K}}M�!?��񥩵@q�).v�ٿ�=jM6�@��N�3@�K}}M�!?��񥩵@�v����ٿXߦ�"�@����3@W���N�!?5�(����@�v����ٿXߦ�"�@����3@W���N�!?5�(����@z�7�ʘٿsMJ�;��@�����3@M�	���!?�a戺�@z�7�ʘٿsMJ�;��@�����3@M�	���!?�a戺�@z�7�ʘٿsMJ�;��@�����3@M�	���!?�a戺�@z�7�ʘٿsMJ�;��@�����3@M�	���!?�a戺�@z�7�ʘٿsMJ�;��@�����3@M�	���!?�a戺�@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@����ٿ��5�f�@_�p�3@�i!�j�!?mHϜ��@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@�#�L��ٿ������@n:�u��3@WB��q�!?�q⊖�@��ҋf�ٿ<���N�@*2)��3@R��⊐!?Ĩ�x�\�@��ҋf�ٿ<���N�@*2)��3@R��⊐!?Ĩ�x�\�@��ҋf�ٿ<���N�@*2)��3@R��⊐!?Ĩ�x�\�@��ҋf�ٿ<���N�@*2)��3@R��⊐!?Ĩ�x�\�@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@ 1�ٿ'+��W��@*�39�3@�>��b�!?��<��@�c�)�ٿ���E�@�x�d�3@-Ú$P�!?blL���@I"�<��ٿ��O���@������3@Zˢh�!?��4F�@I"�<��ٿ��O���@������3@Zˢh�!?��4F�@I"�<��ٿ��O���@������3@Zˢh�!?��4F�@I"�<��ٿ��O���@������3@Zˢh�!?��4F�@I"�<��ٿ��O���@������3@Zˢh�!?��4F�@�D�7&�ٿ�����N�@���& 4@�fNt�!?��?��1�@�D�7&�ٿ�����N�@���& 4@�fNt�!?��?��1�@�D�7&�ٿ�����N�@���& 4@�fNt�!?��?��1�@�D�7&�ٿ�����N�@���& 4@�fNt�!?��?��1�@�D�7&�ٿ�����N�@���& 4@�fNt�!?��?��1�@�Hb�y�ٿ�r���@Ċ|.�4@�WG��!?�f�޳��@�Hb�y�ٿ�r���@Ċ|.�4@�WG��!?�f�޳��@�Hb�y�ٿ�r���@Ċ|.�4@�WG��!?�f�޳��@�Hb�y�ٿ�r���@Ċ|.�4@�WG��!?�f�޳��@�љ8��ٿB��F��@��]u�3@��D/S�!?'��)���@x�$PГٿ����
��@)�VyA�3@��_�!?!�D8�)�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@ɝ�%��ٿl/兯�@���4@F�Kk=�!?�A\�k�@א?>��ٿ��%�>�@�+]T�3@@��!?��E���@X��іٿ����"��@<䏌��3@J��p�!?� #3<��@X��іٿ����"��@<䏌��3@J��p�!?� #3<��@X��іٿ����"��@<䏌��3@J��p�!?� #3<��@f��4Q�ٿnC&F�@!��e�3@<JQ�!?Onh��@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@�q�b�ٿkJ�W�C�@�����3@�-��!?=mT?�@���Օٿ-z8_��@
��2�3@���KS�!?3S8s��@���Օٿ-z8_��@
��2�3@���KS�!?3S8s��@� .���ٿ�e͑[�@=�4@�
�<�!?���l�@��T��ٿ���,$�@*@�L��3@���u�!?sDOP�@��T��ٿ���,$�@*@�L��3@���u�!?sDOP�@��/� �ٿ:�<-��@�ψ�0�3@��4�!?uS� �M�@��/� �ٿ:�<-��@�ψ�0�3@��4�!?uS� �M�@��/� �ٿ:�<-��@�ψ�0�3@��4�!?uS� �M�@��/� �ٿ:�<-��@�ψ�0�3@��4�!?uS� �M�@
��c��ٿ�zh���@��}F��3@��j�1�!?�Q��2�@
��c��ٿ�zh���@��}F��3@��j�1�!?�Q��2�@
��c��ٿ�zh���@��}F��3@��j�1�!?�Q��2�@
��c��ٿ�zh���@��}F��3@��j�1�!?�Q��2�@
��c��ٿ�zh���@��}F��3@��j�1�!?�Q��2�@˸6Ub�ٿ��Ȟ>�@N~[�3@��?M�!?��/У��@���<�ٿ��7gm�@��i/��3@F�&|�!?�gh�k�@���<�ٿ��7gm�@��i/��3@F�&|�!?�gh�k�@���<�ٿ��7gm�@��i/��3@F�&|�!?�gh�k�@	��s��ٿO���\��@@b�s��3@�;�?�!?s�c�-=�@cӈ�5�ٿ�0��_i�@-��ٖ�3@�SM6�!?�Q
;�9�@�!��ٿ�̧�m��@^6��3@��B�'�!?sWhx�@���ٿ��nO���@�@|34@�2(�!?X!d?x�@���ٿ��nO���@�@|34@�2(�!?X!d?x�@���ٿ��nO���@�@|34@�2(�!?X!d?x�@���ٿ��nO���@�@|34@�2(�!?X!d?x�@���ٿ��nO���@�@|34@�2(�!?X!d?x�@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@�<Q剘ٿɞ����@�:#f�3@��_��!?a�Da��@5�_���ٿ=�%<��@Q!׸@�3@��k'I�!?�9��'[�@֎b�B�ٿE���#��@䄒o�3@�>P�'�!?+Ʌ!�X�@֎b�B�ٿE���#��@䄒o�3@�>P�'�!?+Ʌ!�X�@ԯOT��ٿ����q��@a-U���3@� Um�!?��¥<�@ԯOT��ٿ����q��@a-U���3@� Um�!?��¥<�@ԯOT��ٿ����q��@a-U���3@� Um�!?��¥<�@ԯOT��ٿ����q��@a-U���3@� Um�!?��¥<�@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@;T��ٿ[�����@��� 4@i�.��!?��L��մ@�m>� �ٿ���)���@BU�`��3@A��^�!?f�M�>�@�m>� �ٿ���)���@BU�`��3@A��^�!?f�M�>�@�m>� �ٿ���)���@BU�`��3@A��^�!?f�M�>�@�m>� �ٿ���)���@BU�`��3@A��^�!?f�M�>�@�m>� �ٿ���)���@BU�`��3@A��^�!?f�M�>�@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@��%M	�ٿ���k��@C�����3@7,%�k�!?����@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�l:��ٿ�0xG�@�����3@�R]X�!?��x۲C�@�-���ٿ��1$~��@iD���3@���e�!?�玓��@��U<�ٿ��P �c�@�����3@D��i�!?w��\Տ�@��U<�ٿ��P �c�@�����3@D��i�!?w��\Տ�@��U<�ٿ��P �c�@�����3@D��i�!?w��\Տ�@�V-	�ٿ�97	��@i��4o�3@-��(�!?�v>ot��@��ҏٿ����`A�@ �3*Q�3@u~@�!?�B��1�@��ҏٿ����`A�@ �3*Q�3@u~@�!?�B��1�@uU�ϔٿ�P��V�@�A+Z�3@�r��!?�th%�1�@uU�ϔٿ�P��V�@�A+Z�3@�r��!?�th%�1�@uU�ϔٿ�P��V�@�A+Z�3@�r��!?�th%�1�@w����ٿT�����@Yˑ	��3@I3�j�!?����@w����ٿT�����@Yˑ	��3@I3�j�!?����@w����ٿT�����@Yˑ	��3@I3�j�!?����@w����ٿT�����@Yˑ	��3@I3�j�!?����@w����ٿT�����@Yˑ	��3@I3�j�!?����@w����ٿT�����@Yˑ	��3@I3�j�!?����@�-%�n�ٿY�#�8t�@�-N��3@	4!?Ot����@�-%�n�ٿY�#�8t�@�-N��3@	4!?Ot����@�-%�n�ٿY�#�8t�@�-N��3@	4!?Ot����@����՗ٿ���kء�@����3@�a�.��!?�r��m1�@����՗ٿ���kء�@����3@�a�.��!?�r��m1�@�L��ٿ�V��\��@`��3@��═!?�'��?N�@�L��ٿ�V��\��@`��3@��═!?�'��?N�@Ey���ٿ	ꢄ�Q�@�֩ј�3@*�C���!?d^1-��@Ey���ٿ	ꢄ�Q�@�֩ј�3@*�C���!?d^1-��@Ey���ٿ	ꢄ�Q�@�֩ј�3@*�C���!?d^1-��@Ey���ٿ	ꢄ�Q�@�֩ј�3@*�C���!?d^1-��@Ey���ٿ	ꢄ�Q�@�֩ј�3@*�C���!?d^1-��@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�Kx�ϑٿ$�l��.�@#W^�w�3@�-o�Y�!?����}�@�LK��ٿ߽=�/�@���U��3@�e�LM�!?טφ5��@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@�#����ٿ*ʠ�h�@kY�:V�3@��E�!?�\Jв�@��)QC�ٿyZX?��@1��3�3@�l�C�!?h�a7��@��)QC�ٿyZX?��@1��3�3@�l�C�!?h�a7��@��)QC�ٿyZX?��@1��3�3@�l�C�!?h�a7��@��7,4�ٿu-�b���@����3@��6��!?n�o����@�55�=�ٿ�;��L�@�[��L�3@�P��T�!?��\���@�55�=�ٿ�;��L�@�[��L�3@�P��T�!?��\���@  ��ٿ�)�6���@,D1�e�3@����e�!?��:��@2F�*�ٿ<J�`���@���C��3@Ŝ1l{�!?��V�3�@2F�*�ٿ<J�`���@���C��3@Ŝ1l{�!?��V�3�@2F�*�ٿ<J�`���@���C��3@Ŝ1l{�!?��V�3�@b0'�7�ٿ%�ԣ��@�(l��3@@��s7�!?�+/h	�@b0'�7�ٿ%�ԣ��@�(l��3@@��s7�!?�+/h	�@�����ٿ���˲5�@B���+�3@n��0�!?���N"�@�����ٿ���˲5�@B���+�3@n��0�!?���N"�@�����ٿ���˲5�@B���+�3@n��0�!?���N"�@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�FF��ٿC�&&}�@�*f��3@n�K
>�!?eb��@�}j�z�ٿ��ឨ%�@b�r-X�3@X��F`�!?��� l�@�}j�z�ٿ��ឨ%�@b�r-X�3@X��F`�!?��� l�@�}j�z�ٿ��ឨ%�@b�r-X�3@X��F`�!?��� l�@�}j�z�ٿ��ឨ%�@b�r-X�3@X��F`�!?��� l�@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@���f��ٿ1�rf<K�@�Ц���3@�3����!?T����@�qu�ٿ�u�"A��@OZ@��3@qi!?x^���@�qu�ٿ�u�"A��@OZ@��3@qi!?x^���@���*ϔٿ�Ԯa��@��g[��3@�zgê�!?R�wb��@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@V�d�ߕٿ>�X�W�@�`[>��3@Ø9oΐ!?o�����@����H�ٿfr�cW*�@���/�3@w�r��!?��M	��@����H�ٿfr�cW*�@���/�3@w�r��!?��M	��@�!m�i�ٿDǡ��{�@Ww&J4@B	��@�!?�rF��.�@�!m�i�ٿDǡ��{�@Ww&J4@B	��@�!?�rF��.�@�!m�i�ٿDǡ��{�@Ww&J4@B	��@�!?�rF��.�@�^e*�ٿ���g2�@s�3��4@��o�=�!?PLu�?�@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@��#NE�ٿ;���߮�@��k�4@ż�7/�!?���ƴ@�O1K��ٿy�N���@A�vߦ�3@��y��!?b���.B�@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@�N�˘ٿX��f���@�Y1T�3@{vu�d�!?Ec7��@��ŲO�ٿ��|���@B��QH�3@��&�!?:}�ZD�@��ŲO�ٿ��|���@B��QH�3@��&�!?:}�ZD�@��ŲO�ٿ��|���@B��QH�3@��&�!?:}�ZD�@��ŲO�ٿ��|���@B��QH�3@��&�!?:}�ZD�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@6*��5�ٿr0z�V��@J��3�3@t�8<9�!?փO�|s�@q�"ͽ�ٿP*��Z�@-�Y���3@�JZ+�!?uL8sȵ@q�"ͽ�ٿP*��Z�@-�Y���3@�JZ+�!?uL8sȵ@q�"ͽ�ٿP*��Z�@-�Y���3@�JZ+�!?uL8sȵ@q�"ͽ�ٿP*��Z�@-�Y���3@�JZ+�!?uL8sȵ@q�"ͽ�ٿP*��Z�@-�Y���3@�JZ+�!?uL8sȵ@�y2M��ٿj�o�3��@@�)BK�3@�i��:�!?T�Ҡ�@�y2M��ٿj�o�3��@@�)BK�3@�i��:�!?T�Ҡ�@=�+/�ٿ��DF8��@�ZQx�3@�rJgl�!?��<�=�@=�+/�ٿ��DF8��@�ZQx�3@�rJgl�!?��<�=�@����q�ٿ��+��@]G+�k�3@�o�A�!?���4`�@����q�ٿ��+��@]G+�k�3@�o�A�!?���4`�@����q�ٿ��+��@]G+�k�3@�o�A�!?���4`�@atg%j�ٿm����@���
�3@ׂ풒�!?J>ֱ��@���j�ٿ���}��@�I��3@�C�_�!?�'6$���@���j�ٿ���}��@�I��3@�C�_�!?�'6$���@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@��l�ٿ�=s���@��׫�3@�����!?w��,��@�X�VՐٿ���{���@�V�H��3@<P�x�!?ݢI�5�@�X�VՐٿ���{���@�V�H��3@<P�x�!?ݢI�5�@�X�VՐٿ���{���@�V�H��3@<P�x�!?ݢI�5�@�X�VՐٿ���{���@�V�H��3@<P�x�!?ݢI�5�@�X�VՐٿ���{���@�V�H��3@<P�x�!?ݢI�5�@y_�75�ٿp��|�0�@����v�3@�C�O�!?6���@ʈ)��ٿ?�X�[��@�ű��3@i'�FC�!?oq��@�@ʈ)��ٿ?�X�[��@�ű��3@i'�FC�!?oq��@�@�P�B�ٿz�%�{��@�^:M��3@�|� �!?���0�)�@����V�ٿ'�n��@�oij�3@����!?��X;#�@����V�ٿ'�n��@�oij�3@����!?��X;#�@����V�ٿ'�n��@�oij�3@����!?��X;#�@����V�ٿ'�n��@�oij�3@����!?��X;#�@����V�ٿ'�n��@�oij�3@����!?��X;#�@FgՄ�ٿ�8�-�3�@W�%om�3@�CЀ5�!?J9�'�޴@FgՄ�ٿ�8�-�3�@W�%om�3@�CЀ5�!?J9�'�޴@;�uy �ٿ�X�={�@R؍��3@`-��K�!?�D����@;�uy �ٿ�X�={�@R؍��3@`-��K�!?�D����@;�uy �ٿ�X�={�@R؍��3@`-��K�!?�D����@;�uy �ٿ�X�={�@R؍��3@`-��K�!?�D����@;�uy �ٿ�X�={�@R؍��3@`-��K�!?�D����@��!���ٿ/m�����@�.(��3@�\�t�!?R��9��@��!���ٿ/m�����@�.(��3@�\�t�!?R��9��@��!���ٿ/m�����@�.(��3@�\�t�!?R��9��@&!����ٿ�S����@�Э=�3@;�/n/�!?��f�1�@G
��#�ٿJ���=�@��R7Z�3@ACL��!?���/9��@G
��#�ٿJ���=�@��R7Z�3@ACL��!?���/9��@�X��ޒٿ��F�T�@��U���3@����T�!?�gs���@�X��ޒٿ��F�T�@��U���3@����T�!?�gs���@�X��ޒٿ��F�T�@��U���3@����T�!?�gs���@��;p͛ٿt�N�ɐ�@������3@�(� J�!?z�r�nQ�@��;p͛ٿt�N�ɐ�@������3@�(� J�!?z�r�nQ�@��;p͛ٿt�N�ɐ�@������3@�(� J�!?z�r�nQ�@��;p͛ٿt�N�ɐ�@������3@�(� J�!?z�r�nQ�@��;p͛ٿt�N�ɐ�@������3@�(� J�!?z�r�nQ�@�l�؟ٿ ���@,+y��3@4��$�!?��ӈ��@r~Q�8�ٿ���x1�@����3@�C���!?���\$��@r~Q�8�ٿ���x1�@����3@�C���!?���\$��@r~Q�8�ٿ���x1�@����3@�C���!?���\$��@r~Q�8�ٿ���x1�@����3@�C���!?���\$��@{����ٿQ�KM3U�@U�N���3@�X�B�!?��0㵵@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@�P�ٿO�"��@��]��3@���R�!?��K���@X�$3�ٿ��D�Ŵ�@b�r���3@ 0��U�!?8
��@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@s��/��ٿ `Ni�@񽗖H�3@��f�!?�Ϟ�2N�@0�0��ٿ�u�\m�@���=@�3@��7�R�!?��p��Z�@0�0��ٿ�u�\m�@���=@�3@��7�R�!?��p��Z�@0�0��ٿ�u�\m�@���=@�3@��7�R�!?��p��Z�@0�0��ٿ�u�\m�@���=@�3@��7�R�!?��p��Z�@d�	 %�ٿ���U�V�@w��c4@iu �!?�h��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@l��'�ٿ�V����@9֣=�3@� Eg�!?�x�3��@�k=�ٿ�j�+,+�@{��44@�hxv��!?�
S}%�@�k=�ٿ�j�+,+�@{��44@�hxv��!?�
S}%�@2"�e�ٿ%�z�SR�@�>�/4@r�� ��!?����͑�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@�v�p��ٿ@����@��L��3@�-���!?�,�8�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@���`B�ٿ������@GLS.�3@u����!?�t�B�@	wa)&�ٿ�կ��@x*�I�3@O_2�̐!?t���
�@}b�4�ٿ��W��@��#��3@e�G�T�!?"�Ռ.ڴ@o5/x�ٿ��P����@-c;���3@3	P9�!?��l���@�/6~l�ٿ�Nf�Nu�@"Nx�+�3@��۸�!?��L�|��@�"�Gԗٿ$%���8�@L�'���3@v9E{<�!?�S�(v�@�"�Gԗٿ$%���8�@L�'���3@v9E{<�!?�S�(v�@�"�Gԗٿ$%���8�@L�'���3@v9E{<�!?�S�(v�@@!���ٿ{���q��@���O�3@�yBP�!?�pW��@@!���ٿ{���q��@���O�3@�yBP�!?�pW��@�����ٿ�����@?�s�#�3@T�X0�!?��s�2�@�����ٿ�����@?�s�#�3@T�X0�!?��s�2�@�����ٿ�����@?�s�#�3@T�X0�!?��s�2�@�����ٿ�����@?�s�#�3@T�X0�!?��s�2�@�����ٿ�����@?�s�#�3@T�X0�!?��s�2�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@C�A6�ٿJ+z]t��@�6��%�3@={���!?@6�*�@��꾊ٿp�p��@@�9O�3@������!?����i�@�q�3��ٿ�������@Жت��3@��"�I�!?B�I�T�@�q�3��ٿ�������@Жت��3@��"�I�!?B�I�T�@�q�3��ٿ�������@Жت��3@��"�I�!?B�I�T�@�q�3��ٿ�������@Жت��3@��"�I�!?B�I�T�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@���O�ٿ5�VG��@�I�[4@�7��T�!?78��X8�@u���ƙٿ��s�s�@���f��3@"�G�<�!?�wE�V�@u���ƙٿ��s�s�@���f��3@"�G�<�!?�wE�V�@u���ƙٿ��s�s�@���f��3@"�G�<�!?�wE�V�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@���ėٿ��Ӫѱ�@��J&��3@�U���!?�����M�@�q���ٿ�"����@�11F��3@��"G\�!?{�'I�@0��oq�ٿr��r�@��s���3@�J�h�!?��7�̑�@0��oq�ٿr��r�@��s���3@�J�h�!?��7�̑�@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@1�T�ޑٿ�����j�@Go�3@����,�!?��n���@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@Vi�n�ٿ̲����@׀a�.�3@�âR�!?	��x�c�@�G�ҹ�ٿ��m��@ ��4@�~΂Y�!?W=�*]��@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@�-��(�ٿ$9V�@E����3@�cP)�!?���Ե@���k�ٿ����{�@/��%�3@����[�!?�5�~��@���k�ٿ����{�@/��%�3@����[�!?�5�~��@���k�ٿ����{�@/��%�3@����[�!?�5�~��@���k�ٿ����{�@/��%�3@����[�!?�5�~��@���k�ٿ����{�@/��%�3@����[�!?�5�~��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@+�I��ٿ=��B.��@nxB]��3@,�P�v�!?�b(��@	�#�5�ٿ38�]f��@�½:�3@q]t�!?#d�4t�@7v53�ٿ�Ym�ζ�@����3@o�uph�!?�����@7v53�ٿ�Ym�ζ�@����3@o�uph�!?�����@c�2�I�ٿ�p�6�s�@t����3@��ԻI�!?�S�X�@c�2�I�ٿ�p�6�s�@t����3@��ԻI�!?�S�X�@c�2�I�ٿ�p�6�s�@t����3@��ԻI�!?�S�X�@c�2�I�ٿ�p�6�s�@t����3@��ԻI�!?�S�X�@�|��Y�ٿ��S��a�@�P�C��3@T�o�G�!?���5���@�|��Y�ٿ��S��a�@�P�C��3@T�o�G�!?���5���@�|��Y�ٿ��S��a�@�P�C��3@T�o�G�!?���5���@�|��Y�ٿ��S��a�@�P�C��3@T�o�G�!?���5���@�|��Y�ٿ��S��a�@�P�C��3@T�o�G�!?���5���@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@�}��ٿ�2���&�@�j�Ä�3@�1��{�!?���|tS�@_@3-�ٿ"�{c��@�����3@k�j_J�!?¢��Zg�@_@3-�ٿ"�{c��@�����3@k�j_J�!?¢��Zg�@_@3-�ٿ"�{c��@�����3@k�j_J�!?¢��Zg�@_@3-�ٿ"�{c��@�����3@k�j_J�!?¢��Zg�@W�Jl}�ٿ�=��Z<�@���\��3@��<�)�!?�p'�24�@��_�,�ٿ�c�L2�@�
����3@�λ!�!?5�TGwR�@uF٥�ٿ�C�!K�@�R�S�3@�;�3�!?Մ�*{��@uF٥�ٿ�C�!K�@�R�S�3@�;�3�!?Մ�*{��@<1�J�ٿ�cT�o�@&~F��3@��=a�!?c�^q���@<1�J�ٿ�cT�o�@&~F��3@��=a�!?c�^q���@�̳>��ٿ�:�ț�@gu�NY�3@�Z�F�!?���`z�@�U�M�ٿj�-�]�@����3@4]���!?Ҧ��_޵@�O�YޘٿG\-��@�x��3@O��?i�!?4�4���@�O�YޘٿG\-��@�x��3@O��?i�!?4�4���@�O�YޘٿG\-��@�x��3@O��?i�!?4�4���@zM*i��ٿ�51��R�@$FA"�3@7���'�!?,���m�@zM*i��ٿ�51��R�@$FA"�3@7���'�!?,���m�@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@�}��ٿqI�H��@H.0��3@قل�!?KT�!��@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@��-�Жٿ���͏�@A��ƍ�3@�l�槐!?���'5�@����ٿ�&T4~��@�E�(��3@���gk�!?��}�@����ٿ�&T4~��@�E�(��3@���gk�!?��}�@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@�D����ٿ?y{ӥ�@�d.���3@4~]>��!?2��� �@R7���ٿ�)~��@���0��3@)��z��!?D�K��ŵ@R7���ٿ�)~��@���0��3@)��z��!?D�K��ŵ@̱C���ٿ�'>�o�@Ag���3@�_ln�!?��>~��@̱C���ٿ�'>�o�@Ag���3@�_ln�!?��>~��@̱C���ٿ�'>�o�@Ag���3@�_ln�!?��>~��@̱C���ٿ�'>�o�@Ag���3@�_ln�!?��>~��@̱C���ٿ�'>�o�@Ag���3@�_ln�!?��>~��@�%6D'�ٿ�&���@jJ�e4@.J s�!?���*IK�@�%6D'�ٿ�&���@jJ�e4@.J s�!?���*IK�@�%6D'�ٿ�&���@jJ�e4@.J s�!?���*IK�@��4�ٿl�� ��@�<�M�	4@�� ��!?mn1s���@��4�ٿl�� ��@�<�M�	4@�� ��!?mn1s���@kƠp��ٿ@&/����@��g�3@�1���!?R;*4�@kƠp��ٿ@&/����@��g�3@�1���!?R;*4�@kƠp��ٿ@&/����@��g�3@�1���!?R;*4�@LM���ٿ��̈́��@�y3;(�3@Ϝ�rd�!?�	Wv]״@LM���ٿ��̈́��@�y3;(�3@Ϝ�rd�!?�	Wv]״@LM���ٿ��̈́��@�y3;(�3@Ϝ�rd�!?�	Wv]״@LM���ٿ��̈́��@�y3;(�3@Ϝ�rd�!?�	Wv]״@LM���ٿ��̈́��@�y3;(�3@Ϝ�rd�!?�	Wv]״@Ka�ٿh�����@2�%K4@���;d�!?6����
�@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@W��4�ٿqA)jE��@�p��U4@�g�琐!?�����@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@��9��ٿF�A�H�@n���3@�_41��!?�kS_��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@ݠ����ٿ�2˥���@��8���3@G�Ɂ�!?����9��@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@�����ٿ?4`��@��d���3@�U��|�!?�+[����@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@ޛi�͗ٿ�?f���@�����3@�N �*�!?2����$�@lc2+�ٿ��e�Te�@�8�A��3@�MQ.�!?	3�c""�@lc2+�ٿ��e�Te�@�8�A��3@�MQ.�!?	3�c""�@� ��Ôٿr4�c8%�@>́Q��3@�j�
�!?a~|M��@� ��Ôٿr4�c8%�@>́Q��3@�j�
�!?a~|M��@� ��Ôٿr4�c8%�@>́Q��3@�j�
�!?a~|M��@� ��Ôٿr4�c8%�@>́Q��3@�j�
�!?a~|M��@� ��Ôٿr4�c8%�@>́Q��3@�j�
�!?a~|M��@P6Cӿ�ٿ�u@Ve�@��.U��3@�1�Q!�!?���6�@w����ٿT��Z�8�@t����3@�v�(�!?F���Z�@w����ٿT��Z�8�@t����3@�v�(�!?F���Z�@w����ٿT��Z�8�@t����3@�v�(�!?F���Z�@w����ٿT��Z�8�@t����3@�v�(�!?F���Z�@�{�b�ٿ,�(��'�@O���3@��y9�!?O&B��ش@��K	�ٿ�
|���@�h����3@��f�I�!?��[����@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@rz���ٿ��[��@��� 4@{�#�%�!?}qH{�@+�0��ٿ[�Q��@�E.�4@;l�}-�!? '-}�۴@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@*��Z�ٿ��`(��@'�5�.�3@�H��;�!?{q�q�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@ɓ�L��ٿֳ#%���@qS"�R�3@�L]�!?^�#�@n+�?�ٿ?��lL�@A��{��3@X&��Y�!?����I�@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@R��D�ٿU�d����@!���p�3@uz
�T�!?��8���@C
�C�ٿU��fQ�@��̻��3@��>�?�!?��2��@�&�ٿ"��Rs��@	��Z�3@�d���!?FZ-�\+�@�&�ٿ"��Rs��@	��Z�3@�d���!?FZ-�\+�@�&�ٿ"��Rs��@	��Z�3@�d���!?FZ-�\+�@¢�(��ٿz��{���@�����3@��⤐!?�q�	��@>z�T�ٿ��栙��@î2�G�3@">���!?j+~͵@>z�T�ٿ��栙��@î2�G�3@">���!?j+~͵@>z�T�ٿ��栙��@î2�G�3@">���!?j+~͵@Ŧ���ٿ�����@"u���3@�t��|�!?@l�1�@8"f���ٿ�6��p��@�r~L��3@j.��[�!?�).K���@��U�*�ٿ�ϲ�Y�@1��Q"�3@'9O���!?2�0�"�@��U�*�ٿ�ϲ�Y�@1��Q"�3@'9O���!?2�0�"�@�T��ٿ�]��&)�@u��3@
Cς�!?*��$��@�T��ٿ�]��&)�@u��3@
Cς�!?*��$��@�T��ٿ�]��&)�@u��3@
Cς�!?*��$��@�T��ٿ�]��&)�@u��3@
Cς�!?*��$��@�T��ٿ�]��&)�@u��3@
Cς�!?*��$��@ǆS��ٿ1�w���@����8�3@��0�!?8�1��@ǆS��ٿ1�w���@����8�3@��0�!?8�1��@ǆS��ٿ1�w���@����8�3@��0�!?8�1��@Y���ٿĜMP��@� ˰��3@q�A�L�!?}p����@Y���ٿĜMP��@� ˰��3@q�A�L�!?}p����@[R��G�ٿ�e�0�@ (����3@��}��!?,�u�Y�@[R��G�ٿ�e�0�@ (����3@��}��!?,�u�Y�@�."(�ٿjS �-��@?z��3@k1d澐!?�ۄ�)��@}�yd��ٿ�~xl��@�*}&�4@��5G�!?R"d��@}�yd��ٿ�~xl��@�*}&�4@��5G�!?R"d��@}�yd��ٿ�~xl��@�*}&�4@��5G�!?R"d��@| N���ٿ7OM:��@�*�:�3@�����!?����p�@xe&��ٿI=�Y�@�����3@����w�!?b�5��_�@xe&��ٿI=�Y�@�����3@����w�!?b�5��_�@xe&��ٿI=�Y�@�����3@����w�!?b�5��_�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@��ԙ��ٿ�#l����@/y���3@d�[�!?� ��:�@�\��[�ٿ?�lc���@�� ��3@e�}��!?�O��?�@�\��[�ٿ?�lc���@�� ��3@e�}��!?�O��?�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@:V{��ٿV�Pe�@"G�34@Y�f��!?2k�]�@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@�v����ٿ���ԕ��@v6�O�
4@rֈ��!?>����ܴ@(����ٿ�qG�&��@/�^��3@)�`���!?����@(����ٿ�qG�&��@/�^��3@)�`���!?����@(����ٿ�qG�&��@/�^��3@)�`���!?����@(����ٿ�qG�&��@/�^��3@)�`���!?����@(����ٿ�qG�&��@/�^��3@)�`���!?����@(����ٿ�qG�&��@/�^��3@)�`���!?����@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@�R�A��ٿ����	�@j�FtN�3@+�2o��!?�ǯ<��@N�e?�ٿbfϬ���@�:��4@�Ւ�!?��h�e״@N�e?�ٿbfϬ���@�:��4@�Ւ�!?��h�e״@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@H��ϐٿ���χ��@pL�4@tȁP�!?�r�$Qt�@l��}F�ٿ;� ����@��+�3@*�!?+Iȃnx�@l��}F�ٿ;� ����@��+�3@*�!?+Iȃnx�@l��}F�ٿ;� ����@��+�3@*�!?+Iȃnx�@Bۨ�t�ٿ[�k�^�@���?4@��}�׏!?���?���@Bۨ�t�ٿ[�k�^�@���?4@��}�׏!?���?���@��\��ٿ�Ԭ�1�@UU�� 4@�ܐ��!?k��NJ��@��\��ٿ�Ԭ�1�@UU�� 4@�ܐ��!?k��NJ��@��\��ٿ�Ԭ�1�@UU�� 4@�ܐ��!?k��NJ��@��\��ٿ�Ԭ�1�@UU�� 4@�ܐ��!?k��NJ��@rӝ�]�ٿ܃�u��@y�0_�3@-�p�F�!?���[F��@rӝ�]�ٿ܃�u��@y�0_�3@-�p�F�!?���[F��@rӝ�]�ٿ܃�u��@y�0_�3@-�p�F�!?���[F��@rӝ�]�ٿ܃�u��@y�0_�3@-�p�F�!?���[F��@rӝ�]�ٿ܃�u��@y�0_�3@-�p�F�!?���[F��@*���ٿ\'��P�@��Ng�3@�r?��!?��-^��@*���ٿ\'��P�@��Ng�3@�r?��!?��-^��@*���ٿ\'��P�@��Ng�3@�r?��!?��-^��@*���ٿ\'��P�@��Ng�3@�r?��!?��-^��@*���ٿ\'��P�@��Ng�3@�r?��!?��-^��@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@������ٿօN�#�@�&���3@��.7U�!?H�)�y+�@VrM��ٿoI2���@������3@Fa��$�!?�N�#��@VrM��ٿoI2���@������3@Fa��$�!?�N�#��@VrM��ٿoI2���@������3@Fa��$�!?�N�#��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@����ٿ�*��:��@�����3@�j܏!?H�$D3��@ҁ~�D�ٿ�%����@q����3@�N���!?�,&m{��@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�8ل;�ٿŁ�ႁ�@3d[�a�3@��=�!?�m���@�cf"<�ٿ��V���@	>T��3@uT39�!?4l���?�@�cf"<�ٿ��V���@	>T��3@uT39�!?4l���?�@�cf"<�ٿ��V���@	>T��3@uT39�!?4l���?�@�cf"<�ٿ��V���@	>T��3@uT39�!?4l���?�@�cf"<�ٿ��V���@	>T��3@uT39�!?4l���?�@���ٿ;��	�@JWԋ��3@Ͼ�v�!?!���R�@���ٿ;��	�@JWԋ��3@Ͼ�v�!?!���R�@���ٿ;��	�@JWԋ��3@Ͼ�v�!?!���R�@���ٿ;��	�@JWԋ��3@Ͼ�v�!?!���R�@���ٿ;��	�@JWԋ��3@Ͼ�v�!?!���R�@���/�ٿ(�sڠ�@	�?G��3@���x�!?���˰^�@���/�ٿ(�sڠ�@	�?G��3@���x�!?���˰^�@���/�ٿ(�sڠ�@	�?G��3@���x�!?���˰^�@���/�ٿ(�sڠ�@	�?G��3@���x�!?���˰^�@���/�ٿ(�sڠ�@	�?G��3@���x�!?���˰^�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@f2W�H�ٿI������@��p��3@�:�Q�!?�����f�@�̌¨�ٿ{�ϟ��@��Zc��3@FDBWb�!?RCC[�K�@u��L��ٿ1+����@(�� 4@J��!?�]�����@u��L��ٿ1+����@(�� 4@J��!?�]�����@����ٿ��i=�#�@>3�7�3@�w6���!?�ؠsGc�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@2;��"�ٿ:��r���@�����3@�p�b�!?uL��T�@U����ٿ��Ɇ�t�@ߓ� I�3@���T~�!?��})ڴ@U����ٿ��Ɇ�t�@ߓ� I�3@���T~�!?��})ڴ@U����ٿ��Ɇ�t�@ߓ� I�3@���T~�!?��})ڴ@U����ٿ��Ɇ�t�@ߓ� I�3@���T~�!?��})ڴ@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@Ec �N�ٿy������@�W�~�3@(�?�!?)TWàS�@I�g��ٿ������@ª���3@86+��!?׬O�6�@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@�za��ٿ`^�m8V�@I��C�3@n[>��!?G��s��@���d��ٿ����bV�@�L����3@�3M�)�!?�o�l��@ xy�ٿ�u�:Ta�@�-��3@QŊS�!?o��3�@ xy�ٿ�u�:Ta�@�-��3@QŊS�!?o��3�@ xy�ٿ�u�:Ta�@�-��3@QŊS�!?o��3�@ xy�ٿ�u�:Ta�@�-��3@QŊS�!?o��3�@�dR�ٿsB�����@�=��>�3@�Z
.�!?�v�J�@�dR�ٿsB�����@�=��>�3@�Z
.�!?�v�J�@�dR�ٿsB�����@�=��>�3@�Z
.�!?�v�J�@[��2�ٿ�|�l���@������3@��i�T�!?�A��}�@w9�ޔٿzj�K<�@,��[*�3@�U�싐!?��7D��@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@$���ٿ7��+=D�@��N� �3@*}���!?�r��[�@�a(��ٿk�LU]%�@u�.��3@q�#�~�!?-��3���@�a(��ٿk�LU]%�@u�.��3@q�#�~�!?-��3���@z[�n×ٿ;PD�,�@ܔc��3@^��+��!?�a.��q�@z[�n×ٿ;PD�,�@ܔc��3@^��+��!?�a.��q�@r���ٿ� u��@� 9a�3@Kˬ�w�!?@��m�@r���ٿ� u��@� 9a�3@Kˬ�w�!?@��m�@r���ٿ� u��@� 9a�3@Kˬ�w�!?@��m�@c���ٿ0(���2�@�Q���3@5ؙѡ�!?��BG�@c���ٿ0(���2�@�Q���3@5ؙѡ�!?��BG�@c���ٿ0(���2�@�Q���3@5ؙѡ�!?��BG�@c���ٿ0(���2�@�Q���3@5ؙѡ�!?��BG�@�k�.�ٿE���@�S����3@>o�kѐ!?4�z��1�@y70M��ٿ��X3��@�3-v��3@"����!?��st�	�@y70M��ٿ��X3��@�3-v��3@"����!?��st�	�@y70M��ٿ��X3��@�3-v��3@"����!?��st�	�@y70M��ٿ��X3��@�3-v��3@"����!?��st�	�@��d��ٿ
{t��K�@q!,&u4@E����!?<�p�7��@��d��ٿ
{t��K�@q!,&u4@E����!?<�p�7��@��d��ٿ
{t��K�@q!,&u4@E����!?<�p�7��@��d��ٿ
{t��K�@q!,&u4@E����!?<�p�7��@v���?�ٿ4�s�<�@}e�4@��`�!?���yIe�@v���?�ٿ4�s�<�@}e�4@��`�!?���yIe�@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@d�Y���ٿ�z���S�@�2Ώ$4@�Q��d�!?TXh��@l +؞ٿ����E�@��c]�	4@�
�:��!?Z/�=�8�@l +؞ٿ����E�@��c]�	4@�
�:��!?Z/�=�8�@I�/l�ٿ�y��G�@�A'�3@d/[���!?I�q�N�@I�/l�ٿ�y��G�@�A'�3@d/[���!?I�q�N�@I�/l�ٿ�y��G�@�A'�3@d/[���!?I�q�N�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@����ٿ��R���@[z����3@3��\.�!?�mE6>�@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@:"��.�ٿi��<��@S�_���3@q�*�!?ny(/,��@{���m�ٿ@jb����@8,�V�3@=�$��!?Wp���@{���m�ٿ@jb����@8,�V�3@=�$��!?Wp���@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@��}6��ٿ@�^M���@�G8R�3@�|���!?���x��@���ŗٿ�3�-���@���c��3@�?�Ꙑ!?*_���@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@�T�� �ٿ��i���@��_���3@o�*�!?A�ş��@ۨ�aӔٿ��E	��@ʊ�{4@�E�9�!?0�#b��@ۨ�aӔٿ��E	��@ʊ�{4@�E�9�!?0�#b��@ۨ�aӔٿ��E	��@ʊ�{4@�E�9�!?0�#b��@0/�s�ٿ8��~�@��N!'�3@"�!?ôe>���@0/�s�ٿ8��~�@��N!'�3@"�!?ôe>���@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@mݚ�\�ٿ �`)*��@Yʡ�'�3@��@c�!?L�wX�õ@_/��ٿ�b��(F�@5�$K�3@tu�8�!?�eS�"z�@pI6���ٿm۽(@��@�o<�3@���};�!?�/��;*�@pI6���ٿm۽(@��@�o<�3@���};�!?�/��;*�@pI6���ٿm۽(@��@�o<�3@���};�!?�/��;*�@pI6���ٿm۽(@��@�o<�3@���};�!?�/��;*�@pI6���ٿm۽(@��@�o<�3@���};�!?�/��;*�@*���<�ٿ��+�F��@�pv��3@�W�(�!?�U���ݵ@*���<�ٿ��+�F��@�pv��3@�W�(�!?�U���ݵ@�kU�b�ٿ���_�@�F��3@�f�?(�!?���(���@�kU�b�ٿ���_�@�F��3@�f�?(�!?���(���@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@���c�ٿݩ����@�󧙫�3@��X�!?��~��@{ �I�ٿ�
YM��@/^� �3@����=�!?�m���@{ �I�ٿ�
YM��@/^� �3@����=�!?�m���@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@n�/.��ٿD������@_�lA4@'��r?�!?��
�8ε@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@�_Fr�ٿæ(L[�@0Cʡ�3@t���\�!?b%p<��@���A�ٿU�;e�@��)��3@+"X���!?��u_��@���A�ٿU�;e�@��)��3@+"X���!?��u_��@Ё���ٿ�Ѷ��@d���3@&f>8r�!?�#�܇��@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�n��d�ٿ�������@���3��3@t�a�<�!?y[�٨�@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@�2�l��ٿ���0�y�@�צ�#�3@�hx�G�!?9# ���@lX���ٿ�%��@�gR���3@��/	r�!?�9ǃ���@lX���ٿ�%��@�gR���3@��/	r�!?�9ǃ���@lX���ٿ�%��@�gR���3@��/	r�!?�9ǃ���@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@��MBݔٿ.oCw��@b����3@�V��b�!?	G��!�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�M��h�ٿ�Éo���@̧���3@��t8�!?Z�ɞX�@�
8)�ٿ&F��?޿@k2���3@�%	�	�!?�'�*�@�
8)�ٿ&F��?޿@k2���3@�%	�	�!?�'�*�@�
8)�ٿ&F��?޿@k2���3@�%	�	�!?�'�*�@poC�ؕٿ_�ۏ<#�@��b�s4@���!?�G���@poC�ؕٿ_�ۏ<#�@��b�s4@���!?�G���@����ٿ�0\�@��E4@w��u�!?��@��@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�M&v�ٿ�S�����@��9�4@9�1��!?�S�Os)�@�ǳZ�ٿ"����x�@g���F�3@x Mdѐ!?Dg�j�@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@%�
�R�ٿF?�k�K�@�}+t4@ެ�83�!?�L�A��@M��0.�ٿ7�}���@*�En�4@mE�w�!?x?�ŵ@2bu��ٿ���u��@��|`p�3@��:>*�!?X�5ZRõ@2bu��ٿ���u��@��|`p�3@��:>*�!?X�5ZRõ@2bu��ٿ���u��@��|`p�3@��:>*�!?X�5ZRõ@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@�N�^��ٿ��x���@�柾"�3@l��!?UM��̴@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��襞ٿ�{Q�@��sy��3@0ܬ�J�!?�4/��.�@��Խ�ٿ��=��@rXe��4@)�s�(�!?hx?��Y�@��Խ�ٿ��=��@rXe��4@)�s�(�!?hx?��Y�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@�xOLّٿV4�c��@>����3@"��([�!?!���.�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@}X�:�ٿ���E[��@��	���3@߳�IM�!?��D�4�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@�${�z�ٿ�Om�6q�@x�E���3@ȅ�v�!?r�ݗf8�@)�x�ٿ>D+��@eY�9��3@�c	A��!?��+!l��@)�x�ٿ>D+��@eY�9��3@�c	A��!?��+!l��@)�x�ٿ>D+��@eY�9��3@�c	A��!?��+!l��@)�x�ٿ>D+��@eY�9��3@�c	A��!?��+!l��@)�x�ٿ>D+��@eY�9��3@�c	A��!?��+!l��@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@��	՗�ٿ.�"�X��@՜��h�3@�H\�!? �x2�ӵ@#7<�ٿW�a���@%��7�3@���yҐ!?ݖB�0�@#7<�ٿW�a���@%��7�3@���yҐ!?ݖB�0�@���)�ٿ^�*��@�

u4@Il��!?P�Ւ�a�@c��A��ٿ:Fh^�@�l����3@N&�~��!?���s܅�@c��A��ٿ:Fh^�@�l����3@N&�~��!?���s܅�@c��A��ٿ:Fh^�@�l����3@N&�~��!?���s܅�@��5~�ٿd�ɧ���@�r-�m�3@�E	��!?�
��z��@��Ȝq�ٿ-M�u��@�;���3@��(=y�!? 1f��@��Ȝq�ٿ-M�u��@�;���3@��(=y�!? 1f��@��Ȝq�ٿ-M�u��@�;���3@��(=y�!? 1f��@��Ȝq�ٿ-M�u��@�;���3@��(=y�!? 1f��@���O�ٿ�s�B�'�@uU���3@sL@�!?�j��h�@/VƔٿ�|�4��@���j�3@�X���!?y7����@/VƔٿ�|�4��@���j�3@�X���!?y7����@'�
��ٿ@����@�����3@Bb���!?���յ@&=�H&�ٿ��h�h#�@qa�Ȝ�3@p-�!?���@s�vٿb&��ݪ�@��Ȅ��3@Zu5�l�!?��,{�@s�vٿb&��ݪ�@��Ȅ��3@Zu5�l�!?��,{�@s�vٿb&��ݪ�@��Ȅ��3@Zu5�l�!?��,{�@�s�y�ٿ�7��z�@y��DG 4@��[�!?Ĩ9A|j�@�s�y�ٿ�7��z�@y��DG 4@��[�!?Ĩ9A|j�@OdsE�ٿm-*��@7[8�V4@�0�)U�!?�&�(��@OdsE�ٿm-*��@7[8�V4@�0�)U�!?�&�(��@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@�&�ۍ�ٿ%��b�:�@�RU��4@��?�G�!?��W�@��U霖ٿ�?.��L�@Xi&7�3@k�=���!?�Q��%��@�/���ٿ�	y�=�@��w�4@��W�S�!?t�Ɍ��@�/���ٿ�	y�=�@��w�4@��W�S�!?t�Ɍ��@�/���ٿ�	y�=�@��w�4@��W�S�!?t�Ɍ��@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@��]j�ٿ��<���@4�Qo�3@m��9�!?$L�J?�@?s��ٿ�UO��7�@�_.���3@����C�!?#�6��@?s��ٿ�UO��7�@�_.���3@����C�!?#�6��@"���D�ٿ�O�Q)P�@��F�3@WLk�%�!?�3�|��@"���D�ٿ�O�Q)P�@��F�3@WLk�%�!?�3�|��@�cO�ٿW�]֥�@P�gb�3@0��Q�!?��:�̴@pb^o�ٿ�Z ���@��њo�3@ԑ�ԏ!?���#�@pb^o�ٿ�Z ���@��њo�3@ԑ�ԏ!?���#�@R���ʐٿ�?|h�@���u�3@5�$�!?�\�]A�@2���s�ٿnHN���@T ����3@G�M�ߏ!?h���za�@2���s�ٿnHN���@T ����3@G�M�ߏ!?h���za�@��g-�ٿ����H�@�6K�x�3@��� �!?��uNQ	�@��g-�ٿ����H�@�6K�x�3@��� �!?��uNQ	�@��g-�ٿ����H�@�6K�x�3@��� �!?��uNQ	�@��g-�ٿ����H�@�6K�x�3@��� �!?��uNQ	�@��g-�ٿ����H�@�6K�x�3@��� �!?��uNQ	�@����ٿ���{;�@���0��3@�҈�!?%]����@��.�ٿ����z��@H���N�3@F�;�G�!?8��ə�@��.�ٿ����z��@H���N�3@F�;�G�!?8��ə�@��.�ٿ����z��@H���N�3@F�;�G�!?8��ə�@��.�ٿ����z��@H���N�3@F�;�G�!?8��ə�@��.�ٿ����z��@H���N�3@F�;�G�!?8��ə�@�)a�S�ٿ���䡿@^��4��3@��]8�!?<�1����@�NO�%�ٿCE����@�rb���3@Xz��ˏ!?r���@� �$��ٿyM��ڼ�@|C�4@��ُͤ!?��瞵@� �$��ٿyM��ڼ�@|C�4@��ُͤ!?��瞵@� �$��ٿyM��ڼ�@|C�4@��ُͤ!?��瞵@� �$��ٿyM��ڼ�@|C�4@��ُͤ!?��瞵@� �$��ٿyM��ڼ�@|C�4@��ُͤ!?��瞵@�sA��ٿM�����@>)�$��3@|��!?.�P�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@��R�ٿA��U�N�@��U�	4@� w��!?]����7�@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�3v��ٿ�I���p�@<�=���3@��}<M�!?5��@�)-2�ٿ�i���@y�F^t�3@;,���!?��U�s�@������ٿ�^�|��@����3@+{�ɏ!?��~ 0�@�*h��ٿ8��.u�@*�/�4@TBM��!?6�|�v�@�*h��ٿ8��.u�@*�/�4@TBM��!?6�|�v�@�*h��ٿ8��.u�@*�/�4@TBM��!?6�|�v�@�*h��ٿ8��.u�@*�/�4@TBM��!?6�|�v�@���^��ٿ5�(���@�|@h4@&��Q�!?6�ݸbM�@���^��ٿ5�(���@�|@h4@&��Q�!?6�ݸbM�@�.r�ٿtր�`��@"~�E?4@� �0V�!?��t��@�.r�ٿtր�`��@"~�E?4@� �0V�!?��t��@�.r�ٿtր�`��@"~�E?4@� �0V�!?��t��@�.r�ٿtր�`��@"~�E?4@� �0V�!?��t��@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@���`�ٿ3Ե�]��@�W|{�3@���(F�!?���O-�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@5g(�@�ٿm�g�|�@���mQ	4@A}
��!?��~K�W�@ö�_{�ٿ���:���@�H�w4@z�)�!?�Ӆ&�>�@ö�_{�ٿ���:���@�H�w4@z�)�!?�Ӆ&�>�@ö�_{�ٿ���:���@�H�w4@z�)�!?�Ӆ&�>�@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@j.2�I�ٿ$ɏ�k��@)��3@����!?�E����@pv|���ٿF��fRo�@���F�3@�ة?�!?3�@&߇�@pv|���ٿF��fRo�@���F�3@�ة?�!?3�@&߇�@pv|���ٿF��fRo�@���F�3@�ة?�!?3�@&߇�@pv|���ٿF��fRo�@���F�3@�ة?�!?3�@&߇�@pv|���ٿF��fRo�@���F�3@�ة?�!?3�@&߇�@�,�r�ٿ�,x�*�@��wM3�3@�� �R�!?S���=�@�,�r�ٿ�,x�*�@��wM3�3@�� �R�!?S���=�@�,�r�ٿ�,x�*�@��wM3�3@�� �R�!?S���=�@�,�r�ٿ�,x�*�@��wM3�3@�� �R�!?S���=�@�,�r�ٿ�,x�*�@��wM3�3@�� �R�!?S���=�@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@2�(�)�ٿ�s*�?�@�rZ�x�3@�{�Q�!?���!��@6��h�ٿλ�^O��@nF��3@%[�#�!?��k�{ô@6��h�ٿλ�^O��@nF��3@%[�#�!?��k�{ô@6��h�ٿλ�^O��@nF��3@%[�#�!?��k�{ô@6��h�ٿλ�^O��@nF��3@%[�#�!?��k�{ô@6��h�ٿλ�^O��@nF��3@%[�#�!?��k�{ô@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�5�דٿ���a�@b�|���3@�PW4�!?#H����@�s4e�ٿ���v���@cY��3@���=.�!?&�FZ?�@�s4e�ٿ���v���@cY��3@���=.�!?&�FZ?�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�w����ٿ�̤,�@��*�3@���j��!?�!k�P�@�Y����ٿ�/"D@��@J*���3@�;�	=�!?ͻ����@���+^�ٿ11�Zo�@����3@�"
O�!?�D�8�@���+^�ٿ11�Zo�@����3@�"
O�!?�D�8�@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@_�hА�ٿ,�#����@*m�X4@���䀐!?�]�?㬴@gF7)��ٿ.�N���@}y��3@�	�bB�!?e�
�0~�@gF7)��ٿ.�N���@}y��3@�	�bB�!?e�
�0~�@���#
�ٿO����@j$� ��3@y��=�!?2^#�20�@���#
�ٿO����@j$� ��3@y��=�!?2^#�20�@f�����ٿ�+��=�@�7}BY�3@� j�B�!?��ʐ�@��3��ٿY��R���@�����3@rb�^�!?�|�jh�@��3��ٿY��R���@�����3@rb�^�!?�|�jh�@��3��ٿY��R���@�����3@rb�^�!?�|�jh�@��3��ٿY��R���@�����3@rb�^�!?�|�jh�@-m��ٿy;X�R�@����u�3@D��^(�!?��#���@-m��ٿy;X�R�@����u�3@D��^(�!?��#���@-m��ٿy;X�R�@����u�3@D��^(�!?��#���@-m��ٿy;X�R�@����u�3@D��^(�!?��#���@-m��ٿy;X�R�@����u�3@D��^(�!?��#���@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@� ��Y�ٿqSl\�@��E3 �3@,m�SZ�!?�ޒc��@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@A?Xc#�ٿ�r���-�@@`9��3@Eǔ힐!?4�"?p�@YJ�"×ٿ3�򍑧�@s��5P�3@�t𜾐!?��ٓ�@YJ�"×ٿ3�򍑧�@s��5P�3@�t𜾐!?��ٓ�@V<�Y�ٿ+�f&C��@D���3@�'��|�!?l�6�mB�@����w�ٿ�ֱ�@\���3@�4|�0�!?���ը%�@����w�ٿ�ֱ�@\���3@�4|�0�!?���ը%�@����w�ٿ�ֱ�@\���3@�4|�0�!?���ը%�@����w�ٿ�ֱ�@\���3@�4|�0�!?���ը%�@����w�ٿ�ֱ�@\���3@�4|�0�!?���ը%�@���ٿVk�ig�@�x,+��3@�Ur�!?��~Ѵ@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@Q��/5�ٿ(�����@��Є=�3@�J���!?�Y�@�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�w��ٿ�Ye
�*�@��v;�3@ys�š�!?HU��G�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�ꈽT�ٿ������@��{�3@�YzI�!?lt�K�6�@�K��}�ٿp=�75��@[#-D�3@�1��|�!?��	�5ε@�K��}�ٿp=�75��@[#-D�3@�1��|�!?��	�5ε@�K��}�ٿp=�75��@[#-D�3@�1��|�!?��	�5ε@�K��}�ٿp=�75��@[#-D�3@�1��|�!?��	�5ε@�K��}�ٿp=�75��@[#-D�3@�1��|�!?��	�5ε@jwTF��ٿ����~6�@�0���3@œ��q�!?�{D���@jwTF��ٿ����~6�@�0���3@œ��q�!?�{D���@jwTF��ٿ����~6�@�0���3@œ��q�!?�{D���@��ʖٿ�v����@���F��3@a�"�!?�/�s�@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@_A���ٿ���I�@^7V��3@�$+)1�!?��J�*Դ@q��fw�ٿ�]^6�@�����3@��n��!?:��?BU�@�r���ٿ������@��u�3@Ѧ{RS�!?f9�E&�@�r���ٿ������@��u�3@Ѧ{RS�!?f9�E&�@�r���ٿ������@��u�3@Ѧ{RS�!?f9�E&�@�r���ٿ������@��u�3@Ѧ{RS�!?f9�E&�@Lx7��ٿ#n����@�՜Xi�3@[��CJ�!?�$�LH�@Lx7��ٿ#n����@�՜Xi�3@[��CJ�!?�$�LH�@Lx7��ٿ#n����@�՜Xi�3@[��CJ�!?�$�LH�@Lx7��ٿ#n����@�՜Xi�3@[��CJ�!?�$�LH�@���"C�ٿ8��u4�@@h٦r�3@Z�uh'�!?��$��@���"C�ٿ8��u4�@@h٦r�3@Z�uh'�!?��$��@���"C�ٿ8��u4�@@h٦r�3@Z�uh'�!?��$��@���"C�ٿ8��u4�@@h٦r�3@Z�uh'�!?��$��@>��ke�ٿ _j�*�@��c7�3@���v/�!?ҽ�M?�@>��ke�ٿ _j�*�@��c7�3@���v/�!?ҽ�M?�@>��ke�ٿ _j�*�@��c7�3@���v/�!?ҽ�M?�@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@9����ٿ�:˘�=�@��]��4@}��L�!?��Y*��@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@���"ښٿ���km|�@�� �3@�I��O�!?1?��\W�@r��᫘ٿ����@aN���3@)�[A�!?���q�o�@����ٿ��jR3e�@a�T�g4@�c�i�!?P`���@����ٿ��jR3e�@a�T�g4@�c�i�!?P`���@����ٿ��jR3e�@a�T�g4@�c�i�!?P`���@����ٿ��jR3e�@a�T�g4@�c�i�!?P`���@����ٿ��jR3e�@a�T�g4@�c�i�!?P`���@|6��+�ٿ0#�!=�@ѽV��4@���q�!?�9�@|6��+�ٿ0#�!=�@ѽV��4@���q�!?�9�@|6��+�ٿ0#�!=�@ѽV��4@���q�!?�9�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��h͕ٿ��l�c��@K,���4@%�
R|�!?���ı�@��܈�ٿIw���@�����3@��e�O�!?�r�_5�@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@a�7��ٿ�<%��@��}���3@���a$�!?ˈ�1ٴ@�jh�ٿEO���?�@�V�8 4@�'��@�!?����Fƴ@$��ǜٿ�T/����@:��3@CBLA�!?4I�@p�@$��ǜٿ�T/����@:��3@CBLA�!?4I�@p�@$��ǜٿ�T/����@:��3@CBLA�!?4I�@p�@$��ǜٿ�T/����@:��3@CBLA�!?4I�@p�@$��ǜٿ�T/����@:��3@CBLA�!?4I�@p�@)�f�ٿ������@�����3@�y�c�!?� @��@)�f�ٿ������@�����3@�y�c�!?� @��@)�f�ٿ������@�����3@�y�c�!?� @��@�����ٿ���nO�@�/���3@Kr;�!?�ʸ�П�@�����ٿ���nO�@�/���3@Kr;�!?�ʸ�П�@�����ٿ���nO�@�/���3@Kr;�!?�ʸ�П�@ls��ٿ���Ū��@��/�3@m���!?�?��@ls��ٿ���Ū��@��/�3@m���!?�?��@ls��ٿ���Ū��@��/�3@m���!?�?��@ls��ٿ���Ū��@��/�3@m���!?�?��@ls��ٿ���Ū��@��/�3@m���!?�?��@u?����ٿ�JHMk��@?�|yd�3@��j2!�!?Mh�}��@c����ٿ�{=ֹ�@����N�3@�/�g�!?O��`�6�@���əٿӪ�#��@#�W��3@��:�!?Q�l�@r��(y�ٿ2릁Ɉ�@��8I��3@1�B�Y�!?�/?� �@r��(y�ٿ2릁Ɉ�@��8I��3@1�B�Y�!?�/?� �@r��(y�ٿ2릁Ɉ�@��8I��3@1�B�Y�!?�/?� �@r��(y�ٿ2릁Ɉ�@��8I��3@1�B�Y�!?�/?� �@$O��ٿ!�4qn�@,T�aC�3@��ee�!?���u(�@M��E��ٿ!V"��q�@*�����3@����w�!?TG���˴@M��E��ٿ!V"��q�@*�����3@����w�!?TG���˴@M��E��ٿ!V"��q�@*�����3@����w�!?TG���˴@M��E��ٿ!V"��q�@*�����3@����w�!?TG���˴@A����ٿ�rD�5�@�%�7�3@�aѳj�!?n�f�k�@f�}��ٿ��a����@
Vی�3@d����!?N�����@f�}��ٿ��a����@
Vی�3@d����!?N�����@f�}��ٿ��a����@
Vی�3@d����!?N�����@5E�Y�ٿ���L��@�v~�3@O,��7�!?�:�ĵ@5E�Y�ٿ���L��@�v~�3@O,��7�!?�:�ĵ@5E�Y�ٿ���L��@�v~�3@O,��7�!?�:�ĵ@5E�Y�ٿ���L��@�v~�3@O,��7�!?�:�ĵ@��p���ٿuqe�q&�@�rw�3@N>���!?�D�܅��@�a2��ٿ��W���@�k����3@��tJ�!?�eg��@�a2��ٿ��W���@�k����3@��tJ�!?�eg��@�����ٿW�a]u��@Ooނ��3@�E�� �!? �V�Ȓ�@�����ٿW�a]u��@Ooނ��3@�E�� �!? �V�Ȓ�@���|�ٿym�rd�@����7�3@���q�!?`��GɎ�@���|�ٿym�rd�@����7�3@���q�!?`��GɎ�@���|�ٿym�rd�@����7�3@���q�!?`��GɎ�@���|�ٿym�rd�@����7�3@���q�!?`��GɎ�@ Y=�x�ٿn�(�_�@����3@�w���!?d����@ Y=�x�ٿn�(�_�@����3@�w���!?d����@ Y=�x�ٿn�(�_�@����3@�w���!?d����@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@�e�Ҙٿ�0����@�A�(�3@
{J
�!?�T�ɳ�@2A�Z�ٿ* Z�(�@<�X�Q�3@�6r��!?k������@2A�Z�ٿ* Z�(�@<�X�Q�3@�6r��!?k������@Y��ߕٿ��aN;�@92�Zt�3@�vȲ �!?+p�D�@Y��ߕٿ��aN;�@92�Zt�3@�vȲ �!?+p�D�@Y��ߕٿ��aN;�@92�Zt�3@�vȲ �!?+p�D�@�WM��ٿȤ��k�@+o���3@N7w���!?��C��@�WM��ٿȤ��k�@+o���3@N7w���!?��C��@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���"�ٿ����j�@�N���3@�/��:�!?!U~���@���×ٿ�C6<�@h.��3@2[�n�!?��A״@���×ٿ�C6<�@h.��3@2[�n�!?��A״@P\Ƭ$�ٿ��Z7�@�y���3@�V��j�!?�ջp���@P\Ƭ$�ٿ��Z7�@�y���3@�V��j�!?�ջp���@�f�T9�ٿ��|,H��@7ۏQ�3@Yn���!?q�W����@�f�T9�ٿ��|,H��@7ۏQ�3@Yn���!?q�W����@�3�ٿJ&��oM�@Ƅ0]�3@A(�O�!?z�o���@�Q��W�ٿ����tP�@�'��3@U�#��!?ˬ�K�-�@��;��ٿU��^�@��5��3@����!?�Q�
^x�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@�A����ٿ�د�$��@��ܜ#�3@�C�!?k���R�@<�mٕٿ�O�>��@�u����3@��}�!?�ڰz0�@<�mٕٿ�O�>��@�u����3@��}�!?�ڰz0�@1�wn�ٿ%����@��S���3@��k�!?Y��*�@1�wn�ٿ%����@��S���3@��k�!?Y��*�@�\���ٿ!35:
^�@�{]v=�3@��R�`�!?=6ױ1��@�\���ٿ!35:
^�@�{]v=�3@��R�`�!?=6ױ1��@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@ }(��ٿ�:�F�k�@�ʈw�3@sb��A�!?����@S�l�}�ٿ7�!�Ͳ�@e5"�&�3@0� wX�!?��u�е@>�����ٿD���@M�6*�3@��ܱ0�!?�)��-��@>�����ٿD���@M�6*�3@��ܱ0�!?�)��-��@`���ٿ�,�#��@鏢�`�3@Mm���!?�.���s�@`���ٿ�,�#��@鏢�`�3@Mm���!?�.���s�@`���ٿ�,�#��@鏢�`�3@Mm���!?�.���s�@MZ��ٿ��6�E�@^g���3@(?ū�!?�S<'~��@~N��ٿ�(�m'��@��,%b�3@`��1\�!?W"�A}�@������ٿ<G��C,�@�/I��3@D/��a�!?�Xf�z�@������ٿ<G��C,�@�/I��3@D/��a�!?�Xf�z�@������ٿ<G��C,�@�/I��3@D/��a�!?�Xf�z�@������ٿ<G��C,�@�/I��3@D/��a�!?�Xf�z�@������ٿ<G��C,�@�/I��3@D/��a�!?�Xf�z�@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@�%�↔ٿ�8�����@		�g��3@�jW�h�!?��V���@��
�~�ٿg�8sC�@P����3@w�O�!?�D� >�@��
�~�ٿg�8sC�@P����3@w�O�!?�D� >�@ `N��ٿ��H�{��@yE\ ��3@(}>d9�!?������@ `N��ٿ��H�{��@yE\ ��3@(}>d9�!?������@ `N��ٿ��H�{��@yE\ ��3@(}>d9�!?������@ `N��ٿ��H�{��@yE\ ��3@(}>d9�!?������@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@�C�^h�ٿd;�ط/�@�����3@�H���!?:k�O�@3���ɚٿ#͌Ŵ��@~�v�W�3@� ���!?*!�Nڳ�@3���ɚٿ#͌Ŵ��@~�v�W�3@� ���!?*!�Nڳ�@3���ɚٿ#͌Ŵ��@~�v�W�3@� ���!?*!�Nڳ�@��<�P�ٿ��S*$��@��"U�3@�)`k��!?B�;1���@��<�P�ٿ��S*$��@��"U�3@�)`k��!?B�;1���@��<�P�ٿ��S*$��@��"U�3@�)`k��!?B�;1���@��}��ٿ�={5m�@����3@�{��^�!?lKưp�@��}��ٿ�={5m�@����3@�{��^�!?lKưp�@��}��ٿ�={5m�@����3@�{��^�!?lKưp�@5�B)�ٿ`g����@�j�#�3@ܖe��!?����2�@I�h��ٿ`��C�n�@Ӝ� �3@��ֹ&�!?�/�"LT�@��!g��ٿ4��/d_�@ �)�3@��|��!?"ɼ�73�@��!g��ٿ4��/d_�@ �)�3@��|��!?"ɼ�73�@��!g��ٿ4��/d_�@ �)�3@��|��!?"ɼ�73�@��!g��ٿ4��/d_�@ �)�3@��|��!?"ɼ�73�@5B�p�ٿU�jh��@��K�g�3@�v\�8�!?�B-�2��@5B�p�ٿU�jh��@��K�g�3@�v\�8�!?�B-�2��@T@���ٿt�QU��@�O��P4@ՠ��Տ!?��S�^P�@T@���ٿt�QU��@�O��P4@ՠ��Տ!?��S�^P�@T@���ٿt�QU��@�O��P4@ՠ��Տ!?��S�^P�@T@���ٿt�QU��@�O��P4@ՠ��Տ!?��S�^P�@�v�e�ٿ�u�.2��@��L��3@8����!?K��i���@2����ٿ$�v�q�@�Y����3@F><���!?R�z�H�@2����ٿ$�v�q�@�Y����3@F><���!?R�z�H�@���ږٿ�ߘ���@�*��3@o����!?�D��Q��@:ő��ٿ�Д���@�����3@T� ��!?���@	Ѵ@:ő��ٿ�Д���@�����3@T� ��!?���@	Ѵ@:ő��ٿ�Д���@�����3@T� ��!?���@	Ѵ@:ő��ٿ�Д���@�����3@T� ��!?���@	Ѵ@��ߎ
�ٿ��X���@��-��3@���J�!?\�W���@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@ �{7��ٿi��G�f�@8�1i�3@�IY*�!?,�ϖ/��@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@�Wp���ٿ8��\V��@��I D�3@��)�!?�׾� �@���ٿ�����@y�]<�3@b|qr?�!?�x�&ܴ@���ٿ�����@y�]<�3@b|qr?�!?�x�&ܴ@��lH��ٿ���`8�@��I4@����*�!?�Re3I��@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@+N�~�ٿ�S}��@�*��@4@��'a�!?�c�Ur�@���k�ٿ�T�v��@�[T1E�3@
�_�!?~���>Ǵ@���k�ٿ�T�v��@�[T1E�3@
�_�!?~���>Ǵ@���k�ٿ�T�v��@�[T1E�3@
�_�!?~���>Ǵ@2+U>)�ٿ_�1� ��@� sU��3@�/o܈�!?}��Z��@2+U>)�ٿ_�1� ��@� sU��3@�/o܈�!?}��Z��@2+U>)�ٿ_�1� ��@� sU��3@�/o܈�!?}��Z��@����ٿ)x�yD�@D��~��3@R�E�T�!?�2''ش@����ٿ)x�yD�@D��~��3@R�E�T�!?�2''ش@����ٿ)x�yD�@D��~��3@R�E�T�!?�2''ش@����ٿ)x�yD�@D��~��3@R�E�T�!?�2''ش@����ٿ)x�yD�@D��~��3@R�E�T�!?�2''ش@����ٿ�y����@��� @�3@��]�!?�����@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��k��ٿV�tK�c�@�����3@���za�!?�]$`x��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@��ݓٿ��*�(��@d���e�3@�M̯C�!?��d*��@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@�j8�ٿ��0�B;�@��3@�6�*Y�!?�h�ဵ@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@[���͗ٿYE��Q��@&��3@=���h�!?	�^��@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@64�ٿH�S���@wl?x��3@G�YE_�!?w�I�@U�G�ٿ �e,18�@+����3@�$Gw�!?٦�kش@U�G�ٿ �e,18�@+����3@�$Gw�!?٦�kش@�����ٿ��|����@��ӥ��3@�N%ao�!?��N�M�@�����ٿ��|����@��ӥ��3@�N%ao�!?��N�M�@�����ٿ��|����@��ӥ��3@�N%ao�!?��N�M�@u�����ٿ3�e�f�@#��>`�3@o��"'�!?%��Nj�@u�����ٿ3�e�f�@#��>`�3@o��"'�!?%��Nj�@�����ٿdx�tH��@Å�G�3@�&��3�!?sx��-�@�����ٿdx�tH��@Å�G�3@�&��3�!?sx��-�@�,U�ٿ)�H�/��@t�&���3@�M�I��!?����g�@{@2֊�ٿ���|0�@#��Ԃ�3@��6~�!?2VaE斴@{@2֊�ٿ���|0�@#��Ԃ�3@��6~�!?2VaE斴@)��7ٿ_�L*���@�'c�1�3@gum1�!?ۺY	���@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@7\XV��ٿHcl�M|�@A�O�/�3@��0�5�!?��Ї��@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@6ƹ0��ٿ{�jD��@��
�L�3@�9Q�5�!?�0SYȴ@�D�b�ٿ����*�@�����3@��6�!?Q�}$�Ӵ@�D�b�ٿ����*�@�����3@��6�!?Q�}$�Ӵ@�S|ۢ�ٿ��c�@%߫x*�3@2q�o@�!?�ې`�@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@�h�s�ٿ`�,r���@Vԣھ�3@J�*�!?�<U���@���A�ٿ1���;��@@��k�3@�'�2�!?�h��@���A�ٿ1���;��@@��k�3@�'�2�!?�h��@���A�ٿ1���;��@@��k�3@�'�2�!?�h��@���A�ٿ1���;��@@��k�3@�'�2�!?�h��@-��=�ٿ-�i�1X�@���a�3@Ŗ��!?�V�⎵@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@`L4$��ٿ<U�p��@�����3@ˆx�[�!?��q~2 �@&�󡮚ٿE�&Q9�@����3@}4$+F�!?�ŜV�@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�l�.>�ٿ�9����@`O|�3@$I�?Y�!?�ُ���@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@�ɗ��ٿU<K����@�Hxw�4@���9�!?�.֞��@'�+��ٿ�s�7�u�@����;�3@�z��!?z:����@'�+��ٿ�s�7�u�@����;�3@�z��!?z:����@�>�ǘٿ��,��@<0p|E�3@}h���!?��ZZ�@�>�ǘٿ��,��@<0p|E�3@}h���!?��ZZ�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@��c�}�ٿ�.���@�{���3@�$��!?�`v4t�@�g�ٿw�=����@ab�V��3@���=7�!?�X q9��@�g�ٿw�=����@ab�V��3@���=7�!?�X q9��@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@�'���ٿ������@&��ZC�3@1"\�,�!?$���j�@���!ݙٿ�t�'s��@pR�P��3@�o��ߏ!?^q�,�@�:��ޒٿs7;nC��@�'��3@)����!?(�DMo�@+<#�ٿx$&���@��U�	�3@����!?U�媕ص@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@�@�^�ٿp�P�R�@7:���3@l�D �!?�s��X��@.�Zߑٿ*h�A�Z�@��9�5�3@~B/yǏ!?_�#��w�@.�Zߑٿ*h�A�Z�@��9�5�3@~B/yǏ!?_�#��w�@�x���ٿZQ ���@l�?�3@+��ɏ!??�Z�Rش@�ab��ٿ�ZT���@ڶ�7�3@��_E�!?i��j	��@�ab��ٿ�ZT���@ڶ�7�3@��_E�!?i��j	��@�ab��ٿ�ZT���@ڶ�7�3@��_E�!?i��j	��@�ab��ٿ�ZT���@ڶ�7�3@��_E�!?i��j	��@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@F,��ٿ�S�&�@�4�Z��3@N�l�!?��Pp���@�3�&Ùٿ�aП�]�@؁"v�3@}@����!?[��EG�@�3�&Ùٿ�aП�]�@؁"v�3@}@����!?[��EG�@�3�&Ùٿ�aП�]�@؁"v�3@}@����!?[��EG�@�3�&Ùٿ�aП�]�@؁"v�3@}@����!?[��EG�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@�QW��ٿ�I}���@�q^�3@��va�!?���#�@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@T>��p�ٿ����b�@�e ���3@��,b]�!?dt=����@h/��ٿl���:�@	�g�3@�cyo�!?Yʜ��@��{�ٿ]��W�I�@s�i��3@�o�;�!?elޮ��@�|N�ٿ�O
�@q����3@*��O�!?=���<�@�|N�ٿ�O
�@q����3@*��O�!?=���<�@Lc�jF�ٿ��c�Y@�@y���3@�z�	�!?e7by�@Lc�jF�ٿ��c�Y@�@y���3@�z�	�!?e7by�@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@-{���ٿdmWE"��@�,Xe�3@Y�U�!?����"��@�7��ٿ��j�P��@>j8b��3@�ր.M�!?�&����@�7��ٿ��j�P��@>j8b��3@�ր.M�!?�&����@�7��ٿ��j�P��@>j8b��3@�ր.M�!?�&����@�1ǆ��ٿr2Hn�2�@���3@/��$y�!?i2t4!�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@���ȳ�ٿ�
ۅi��@�d��� 4@�x/j��!?��`L"�@��f��ٿp�*[��@b���l�3@ {0汐!?a�(\��@��f��ٿp�*[��@b���l�3@ {0汐!?a�(\��@��f��ٿp�*[��@b���l�3@ {0汐!?a�(\��@��f��ٿp�*[��@b���l�3@ {0汐!?a�(\��@��f��ٿp�*[��@b���l�3@ {0汐!?a�(\��@`7=p��ٿ�)�{�@ӱ��1�3@�W��O�!?�����&�@`7=p��ٿ�)�{�@ӱ��1�3@�W��O�!?�����&�@`7=p��ٿ�)�{�@ӱ��1�3@�W��O�!?�����&�@`7=p��ٿ�)�{�@ӱ��1�3@�W��O�!?�����&�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@)�#��ٿﷴF�@���vy�3@;ԯI�!?���Cn,�@�V�ᢎٿ�y�J��@�����3@06�U�!?����PP�@�k�/��ٿ���`���@�ee���3@?��W��!?�$�+�@�k�/��ٿ���`���@�ee���3@?��W��!?�$�+�@�k�/��ٿ���`���@�ee���3@?��W��!?�$�+�@�k�/��ٿ���`���@�ee���3@?��W��!?�$�+�@s(V:�ٿ���T���@��%:>�3@3��;��!?TӅ_��@s(V:�ٿ���T���@��%:>�3@3��;��!?TӅ_��@Bw��ȖٿIwF�J��@��vl�3@Z����!?2O�@Bw��ȖٿIwF�J��@��vl�3@Z����!?2O�@Bw��ȖٿIwF�J��@��vl�3@Z����!?2O�@Bw��ȖٿIwF�J��@��vl�3@Z����!?2O�@Bw��ȖٿIwF�J��@��vl�3@Z����!?2O�@�/����ٿ:���@�r��3@��&��!?�e���@�Qd�/�ٿs�s��B�@�%��3@��g�Ɛ!?[�����@K��;�ٿ/<ˋ\,�@�z��3@K�\c��!?����Ѵ@K��;�ٿ/<ˋ\,�@�z��3@K�\c��!?����Ѵ@K��;�ٿ/<ˋ\,�@�z��3@K�\c��!?����Ѵ@Z����ٿ��$��@�S���3@Nw��N�!?�?a�b��@DP�W*�ٿ����6n�@�L����3@�n�L�!?�Gw�/�@DP�W*�ٿ����6n�@�L����3@�n�L�!?�Gw�/�@DP�W*�ٿ����6n�@�L����3@�n�L�!?�Gw�/�@6�+Rƚٿ:bZ��@����3@QKi��!?��U�-��@����ٿKD!� ��@`�$�3@qλ�!�!?�hIE�׵@����ٿKD!� ��@`�$�3@qλ�!�!?�hIE�׵@����ٿKD!� ��@`�$�3@qλ�!�!?�hIE�׵@����ٿKD!� ��@`�$�3@qλ�!�!?�hIE�׵@����ٿKD!� ��@`�$�3@qλ�!�!?�hIE�׵@͐�$�ٿ����IZ�@;�,��3@ڦ�=�!?��U�u��@͐�$�ٿ����IZ�@;�,��3@ڦ�=�!?��U�u��@3-��'�ٿD*jA���@{���3@���9@�!?�eB�;��@3-��'�ٿD*jA���@{���3@���9@�!?�eB�;��@3-��'�ٿD*jA���@{���3@���9@�!?�eB�;��@3-��'�ٿD*jA���@{���3@���9@�!?�eB�;��@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@�V%C��ٿ�dex�@z(�KQ�3@r����!?[# �ڴ@��d�ٿi��q�@��Ν��3@|�y�j�!?�!��r�@��d�ٿi��q�@��Ν��3@|�y�j�!?�!��r�@���Zۑٿ<8��
��@9ڻ>~�3@�_�^K�!?������@���Zۑٿ<8��
��@9ڻ>~�3@�_�^K�!?������@���Zۑٿ<8��
��@9ڻ>~�3@�_�^K�!?������@���Zۑٿ<8��
��@9ڻ>~�3@�_�^K�!?������@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�澹˛ٿ���q���@{�R��3@{��׆�!?��E�Zش@�Z)۝ٿm�V�}�@�4H��3@�o��(�!?{��}��@�Z)۝ٿm�V�}�@�4H��3@�o��(�!?{��}��@�Z)۝ٿm�V�}�@�4H��3@�o��(�!?{��}��@/P�k@�ٿ
� ��/�@@rd	�3@�aS���!?L�.@�@/P�k@�ٿ
� ��/�@@rd	�3@�aS���!?L�.@�@/P�k@�ٿ
� ��/�@@rd	�3@�aS���!?L�.@�@/P�k@�ٿ
� ��/�@@rd	�3@�aS���!?L�.@�@/P�k@�ٿ
� ��/�@@rd	�3@�aS���!?L�.@�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@{ԧ�ٿ��xT��@q��(�3@c+�Ő!?��nj�(�@H@��4�ٿ���h:<�@2$g��3@��b�M�!?H�J���@H@��4�ٿ���h:<�@2$g��3@��b�M�!?H�J���@H@��4�ٿ���h:<�@2$g��3@��b�M�!?H�J���@H@��4�ٿ���h:<�@2$g��3@��b�M�!?H�J���@R~ǐ��ٿ{��4��@ע}Dj�3@�+V/�!?ץ�)��@R~ǐ��ٿ{��4��@ע}Dj�3@�+V/�!?ץ�)��@R~ǐ��ٿ{��4��@ע}Dj�3@�+V/�!?ץ�)��@R~ǐ��ٿ{��4��@ע}Dj�3@�+V/�!?ץ�)��@nQ�x�ٿ��A���@�Ѯ�3@ٝ��Y�!?�.Y�`�@nQ�x�ٿ��A���@�Ѯ�3@ٝ��Y�!?�.Y�`�@�Q��<�ٿ-�0Rj�@r�1�3@#�US>�!?S0�y���@I.�ٿ�"#�Ӽ�@�P� ��3@_�Ԇ�!?�Pf*Ǵ@I.�ٿ�"#�Ӽ�@�P� ��3@_�Ԇ�!?�Pf*Ǵ@I.�ٿ�"#�Ӽ�@�P� ��3@_�Ԇ�!?�Pf*Ǵ@m^�=�ٿ������@Ї�n0�3@�@{]�!?/���׸�@m^�=�ٿ������@Ї�n0�3@�@{]�!?/���׸�@m^�=�ٿ������@Ї�n0�3@�@{]�!?/���׸�@m^�=�ٿ������@Ї�n0�3@�@{]�!?/���׸�@m^�=�ٿ������@Ї�n0�3@�@{]�!?/���׸�@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@)��Ѡ�ٿ;"y�'�@��V�3@�9�{P�!?e�v'���@�G�	�ٿ�?2H	��@ ���3@纫��!? 7%h�@�G�	�ٿ�?2H	��@ ���3@纫��!? 7%h�@��d:�ٿF�Xl�@�ʬ��3@a-e�!?��E$���@��d:�ٿF�Xl�@�ʬ��3@a-e�!?��E$���@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@��n��ٿ�&���l�@I�'��3@cQ�q�!?��-��@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@O���ٿ��؁���@�`�ާ�3@Y�Âr�!?�
 ���@6�3X}�ٿ_�#)���@���c�3@�o����!?���I�@6�3X}�ٿ_�#)���@���c�3@�o����!?���I�@6�3X}�ٿ_�#)���@���c�3@�o����!?���I�@6�3X}�ٿ_�#)���@���c�3@�o����!?���I�@6�3X}�ٿ_�#)���@���c�3@�o����!?���I�@���D��ٿ�3�Ϥ�@�])���3@��>��!?�@m�~ƴ@���D��ٿ�3�Ϥ�@�])���3@��>��!?�@m�~ƴ@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�y5���ٿ�*�����@xwC�#�3@�$�<�!?�cϴQ��@�V���ٿ{P8��@��7)�3@r�[6��!?�||7Kϴ@�V���ٿ{P8��@��7)�3@r�[6��!?�||7Kϴ@�V���ٿ{P8��@��7)�3@r�[6��!?�||7Kϴ@��{χ�ٿl^�B��@��"M�3@��҉�!?���R�T�@m��z�ٿ(��E���@aѷ�o�3@LP;a��!?B*�׵δ@6����ٿ��V�@D�~��3@�.;�!?B�A�ִ@���f�ٿ0�0qU�@�7��3@��U@�!?�`kw�@���f�ٿ0�0qU�@�7��3@��U@�!?�`kw�@���f�ٿ0�0qU�@�7��3@��U@�!?�`kw�@>_(V�ٿ_M%$�k�@i�5��3@䋧��!?.����A�@>_(V�ٿ_M%$�k�@i�5��3@䋧��!?.����A�@�m�Q�ٿ�v��s�@.k��3@��ꄪ�!?P
U.��@�m�Q�ٿ�v��s�@.k��3@��ꄪ�!?P
U.��@�m�Q�ٿ�v��s�@.k��3@��ꄪ�!?P
U.��@�m�Q�ٿ�v��s�@.k��3@��ꄪ�!?P
U.��@V���ٿ�}�lu�@����3@ ��ؐ!?�&��@V���ٿ�}�lu�@����3@ ��ؐ!?�&��@V���ٿ�}�lu�@����3@ ��ؐ!?�&��@V���ٿ�}�lu�@����3@ ��ؐ!?�&��@V���ٿ�}�lu�@����3@ ��ؐ!?�&��@��.�/�ٿJ���@�Z��4@~���!?��!�@��.�/�ٿJ���@�Z��4@~���!?��!�@��.�/�ٿJ���@�Z��4@~���!?��!�@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@�UЍ��ٿ�+�8p��@���
4@_���s�!?���w��@ǝ7P�ٿ�������@t���3@T��ૐ!?zcҖ�o�@ǝ7P�ٿ�������@t���3@T��ૐ!?zcҖ�o�@��1�`�ٿR#�j/r�@ � ��3@u>�?�!?�fIc�a�@��1�`�ٿR#�j/r�@ � ��3@u>�?�!?�fIc�a�@�R0��ٿ���!���@�^�?)�3@9aW\�!?����	��@�R0��ٿ���!���@�^�?)�3@9aW\�!?����	��@�R0��ٿ���!���@�^�?)�3@9aW\�!?����	��@_6���ٿ��j���@�W*�3@k�,z<�!?�����@_6���ٿ��j���@�W*�3@k�,z<�!?�����@_6���ٿ��j���@�W*�3@k�,z<�!?�����@#�+R)�ٿ���&Da�@e����3@�a�$�!?ݙ+c�t�@�����ٿ�j����@��*k�3@e��$1�!?�!����@�����ٿ�j����@��*k�3@e��$1�!?�!����@�����ٿ�j����@��*k�3@e��$1�!?�!����@�����ٿ�j����@��*k�3@e��$1�!?�!����@�����ٿ�j����@��*k�3@e��$1�!?�!����@a��l^�ٿ��?Y�g�@ms�z�3@��k��!?��d25Ŵ@a��l^�ٿ��?Y�g�@ms�z�3@��k��!?��d25Ŵ@a��l^�ٿ��?Y�g�@ms�z�3@��k��!?��d25Ŵ@a��l^�ٿ��?Y�g�@ms�z�3@��k��!?��d25Ŵ@a��l^�ٿ��?Y�g�@ms�z�3@��k��!?��d25Ŵ@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@6�E�ʚٿ�&f�k�@PDs���3@,w���!?d��R3}�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@������ٿ     ��@      4@�t><K�!?�<��4A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@���ٿ��m ��@���? 4@��	�J�!?���H5A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�q��ٿ�4]) ��@��A 4@�V�Z�!?�15A�@�֣|�ٿ�.�# ��@>��9 4@bgY�!?o�@	5A�@�֣|�ٿ�.�# ��@>��9 4@bgY�!?o�@	5A�@�֣|�ٿ�.�# ��@>��9 4@bgY�!?o�@	5A�@�x��יٿl� ��@(�� 4@`�芐!?���4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��Y�ٿOd6 ��@��i� 4@c��� �!?n��4A�@��w���ٿ��$ ��@�<E 4@�ُ!?.��4A�@��w���ٿ��$ ��@�<E 4@�ُ!?.��4A�@��(8��ٿ��� ��@�2�� 4@H�jɀ�!?Yb��4A�@��(8��ٿ��� ��@�2�� 4@H�jɀ�!?Yb��4A�@�﹮�ٿp� ��@�{�� 4@�����!?�C�5A�@Q�HݙٿC�� ��@q�p 4@Q6C[�!?�T5A�@��֙ٿ� ��@~�		 4@�R���!?��O 5A�@��֙ٿ� ��@~�		 4@�R���!?��O 5A�@��֙ٿ� ��@~�		 4@�R���!?��O 5A�@��֙ٿ� ��@~�		 4@�R���!?��O 5A�@�ݥٙٿ1�= ��@��X 4@��r��!?Y���4A�@�)֙ٿF}f ��@A��� 4@�'���!?��E5A�@����ٿ�8�����@)��� 4@�_!�!?;}�5A�@����ٿ�8�����@)��� 4@�_!�!?;}�5A�@����ٿ�8�����@)��� 4@�_!�!?;}�5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@t��ߙٿ��?����@�W!	 4@���i>�!?�O)5A�@pL�!��ٿ9�s����@��s�	 4@y~���!?�/5A�@pL�!��ٿ9�s����@��s�	 4@y~���!?�/5A�@pL�!��ٿ9�s����@��s�	 4@y~���!?�/5A�@���@ߙٿn������@<�
 4@��SB��!?���I5A�@���@ߙٿn������@<�
 4@��SB��!?���I5A�@�	��ۙٿ��8����@X��
 4@����(�!?�.K5A�@��3Sۙٿ� i����@�9
 4@����{�!?���>5A�@��3Sۙٿ� i����@�9
 4@����{�!?���>5A�@��3Sۙٿ� i����@�9
 4@����{�!?���>5A�@��3Sۙٿ� i����@�9
 4@����{�!?���>5A�@��3Sۙٿ� i����@�9
 4@����{�!?���>5A�@8r~ՙٿ6$�����@+��_ 4@�:G�!?}�n85A�@8r~ՙٿ6$�����@+��_ 4@�:G�!?}�n85A�@Ւa�ܙٿ�f����@�5�� 4@�I[懐!?�v�95A�@Ւa�ܙٿ�f����@�5�� 4@�I[懐!?�v�95A�@�q��ٿ�r�����@z�� 4@L_P�!?G��E5A�@�$���ٿӭ�����@+� 4@:�@��!?�z�T5A�@�$���ٿӭ�����@+� 4@:�@��!?�z�T5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@'�ŷ��ٿ�y����@A^pA 4@'�i*�!?���[5A�@ ~��ٿ������@��I 4@�����!?p�\5A�@ ~��ٿ������@��I 4@�����!?p�\5A�@ ~��ٿ������@��I 4@�����!?p�\5A�@z_Mݙٿ�t�����@9��C 4@���/a�!?xs�K5A�@z_Mݙٿ�t�����@9��C 4@���/a�!?xs�K5A�@�Rmߙٿ+�����@���" 4@�e�s�!?ҊZ5A�@�Rmߙٿ+�����@���" 4@�e�s�!?ҊZ5A�@p s��ٿ3?u����@ƍ�  4@@ �Lq�!?P=P5A�@��Q��ٿ��O����@N�p 4@4�c��!?>�hN5A�@��Q��ٿ��O����@N�p 4@4�c��!?>�hN5A�@��L��ٿ������@F�} 4@�k
k�!?9x|M5A�@��L��ٿ������@F�} 4@�k
k�!?9x|M5A�@��L��ٿ������@F�} 4@�k
k�!?9x|M5A�@z)>i�ٿA������@��U� 4@lb%�!?�^D5A�@�����ٿV.[����@��� 4@K��E�!?	��E5A�@�����ٿV.[����@��� 4@K��E�!?	��E5A�@�����ٿV.[����@��� 4@K��E�!?	��E5A�@�����ٿV.[����@��� 4@K��E�!?	��E5A�@B�ܙٿ2������@b�6 4@l�?�J�!?n��P5A�@+\oAڙٿ�'�����@L�7� 4@���c�!?���F5A�@�`a"ۙٿ�ö����@e�%J 4@䕼���!?���R5A�@��ؙٿ�J�����@���o 4@���U�!?XU�S5A�@��ؙٿ�J�����@���o 4@���U�!?XU�S5A�@���kؙٿ�������@�j�X 4@��=틐!?�2�V5A�@��Oԙٿ0�9����@ Ni� 4@���|��!?:��R5A�@�=ڙٿn�j����@"u 4@�`t�!?��FL5A�@O?}�ٙٿ*�<����@{P� 4@����~�!?��H5A�@+�>ՙٿg�� ��@�\J� 4@%�:E�!?���M5A�@+�>ՙٿg�� ��@�\J� 4@%�:E�!?���M5A�@+�>ՙٿg�� ��@�\J� 4@%�:E�!?���M5A�@^=��ҙٿ� ��@�.�* 4@�`-�8�!?��H5A�@^=��ҙٿ� ��@�.�* 4@�`-�8�!?��H5A�@�02	әٿ]ɻ ��@�MV
 4@����!?P�=5A�@�02	әٿ]ɻ ��@�MV
 4@����!?P�=5A�@�02	әٿ]ɻ ��@�MV
 4@����!?P�=5A�@x+��ՙٿ�N�! ��@2��	 4@��:�l�!?
�E65A�@x+��ՙٿ�N�! ��@2��	 4@��:�l�!?
�E65A�@_ɩԙٿ=$ ��@
�8	 4@M�>�M�!?��45A�@_ɩԙٿ=$ ��@
�8	 4@M�>�M�!?��45A�@��P|әٿ��) ��@-��� 4@/0�!?��*5A�@u,?.ԙٿ/ E. ��@���� 4@�m"Y�!?�~	&5A�@���ٙٿ�<�, ��@Q�p� 4@�6��d�!?�ml5A�@�\�Eՙٿ��&& ��@٩~� 4@�:>}�!?4�5A�@'}̿ՙٿWL�# ��@��2� 4@��e���!?�Q5A�@�-љٿ�6 ��@I  4@����!?E'5A�@��Qҙٿ��f ��@p� 4@ѣ� �!?�KK5A�@�}7̙ٿ��& ��@x?�� 4@���M�!?��
5A�@��{�əٿ*r�, ��@�� 4@
!��!?���5A�@��{�əٿ*r�, ��@�� 4@
!��!?���5A�@��Gƙٿ���8 ��@QV�* 4@�0�;�!?�L��4A�@Xa�ƙٿ��? ��@0"dR 4@ݣAMZ�!?�Nv�4A�@��g�Ǚٿp�vJ ��@�� 4@�ڙ�$�!?5��4A�@��g�Ǚٿp�vJ ��@�� 4@�ڙ�$�!?5��4A�@˵Q�řٿXrJ ��@�w�� 4@����2�!?$ �4A�@/2��ęٿaۙS ��@`�  4@D��1�!?�B��4A�@�l���ٿ��Z ��@P�,  4@ڬ2(d�!?%���4A�@��k��ٿj,^t ��@myx��3@ݺ��z�!?�|U�4A�@�@ϻ�ٿ�&�w ��@������3@b�؀5�!?��ø4A�@@OaK��ٿ�\} ��@��Q��3@�+��!?)��4A�@���Ùٿ���� ��@QL��3@֝���!?҂��4A�@���Ùٿ���� ��@QL��3@֝���!?҂��4A�@���Ùٿ���� ��@QL��3@֝���!?҂��4A�@ཊ���ٿu�� ��@�S���3@��i�a�!?6�ԡ4A�@Fk5쿙ٿ�$�� ��@0���3@���`�!?Xl��4A�@6�j�ęٿ��$r ��@��S|��3@��d=5�!?)0q�4A�@8d�ƙٿ�V3x ��@�T����3@3\@�!?v5�4A�@�o.�řٿt�o� ��@2�mE��3@��'x�!?i>�4A�@�o.�řٿt�o� ��@2�mE��3@��'x�!?i>�4A�@���ƙٿU*� ��@[�t ��3@�a+y��!?�LF�4A�@��0yʙٿAR>� ��@;k���3@7^ ���!?ۖ��4A�@��0yʙٿAR>� ��@;k���3@7^ ���!?ۖ��4A�@×̙ٿ�E~ ��@��p��3@�/���!?��4A�@×̙ٿ�E~ ��@��p��3@�/���!?��4A�@�i��͙ٿ�`-z ��@z�} 4@b����!?�-�4A�@;�sϙٿ0��~ ��@�%I�  4@�W1���!?���4A�@;�sϙٿ0��~ ��@�%I�  4@�W1���!?���4A�@;�sϙٿ0��~ ��@�%I�  4@�W1���!?���4A�@��i�əٿ�.'� ��@�W7���3@��2���!?J[��4A�@��i�əٿ�.'� ��@�W7���3@��2���!?J[��4A�@��i�əٿ�.'� ��@�W7���3@��2���!?J[��4A�@l��Ǚٿ0�{ ��@��[  4@o Lȯ�!?�<g�4A�@l��Ǚٿ0�{ ��@��[  4@o Lȯ�!?�<g�4A�@l��Ǚٿ0�{ ��@��[  4@o Lȯ�!?�<g�4A�@l��Ǚٿ0�{ ��@��[  4@o Lȯ�!?�<g�4A�@��,ęٿ��� ��@���!��3@�E���!?���4A�@��,ęٿ��� ��@���!��3@�E���!?���4A�@oUI�˙ٿ��to ��@�j�� 4@d��(ɐ!?�H�4A�@=�Ev̙ٿSwDx ��@]U_s 4@NR�n!?|@�4A�@��_�ϙٿ�B�] ��@3͠� 4@ݱ��]�!?�y6�4A�@݈��љٿu(�^ ��@�NB 4@���_�!?�%K�4A�@D�y�әٿmVCW ��@a�� 4@$��U�!?@ͥ�4A�@Ɛ��Йٿ���M ��@�F�; 4@�
/4�!?���4A�@����ԙٿxZ> ��@8�. 4@�l��!?��5A�@�#�9֙ٿ!�E ��@j� 4@��=S�!?�R*�4A�@�#�9֙ٿ!�E ��@j� 4@��=S�!?�R*�4A�@����˙ٿ��y ��@7L��  4@�>�`��!?��v�4A�@�lI֙ٿ-��O ��@�3� 4@4�I`�!?u���4A�@Ż}�ؙٿO��a ��@�{2 4@�I��~�!?�d�4A�@ݫ Aڙٿ{5]b ��@6Js	 4@5w���!?[w|�4A�@��;ۙٿ�B�o ��@�^� 4@��{2�!?Ո|�4A�@�/Bٙٿ��X ��@X��e 4@���7�!?֗�5A�@I��(ٙٿ���^ ��@j�  4@�_S�)�!?;r��4A�@ys?ٙٿ�7�} ��@�sf 4@g�Q�(�!?�R��4A�@ys?ٙٿ�7�} ��@�sf 4@g�Q�(�!?�R��4A�@�l�!ڙٿ�FOd ��@Ee$E 4@\�@pt�!?�I��4A�@Y�W�ڙٿ��y ��@Q�~� 4@5�1��!?u���4A�@�Qvڙٿ�	�o ��@�MG 4@�9�ꃐ!?�p�5A�@�Qvڙٿ�	�o ��@�MG 4@�9�ꃐ!?�p�5A�@S���ڙٿ� _ ��@QK�� 4@ڠ,�a�!?���5A�@r_�Sؙٿ���` ��@YԿS 4@�4@~=�!?��5A�@p|0�ҙٿ/��l ��@R��� 4@�A�A�!?J���4A�@cA�Ιٿ�� ��@���-  4@�;DX1�!?��t�4A�@cA�Ιٿ�� ��@���-  4@�;DX1�!?��t�4A�@�.z�љٿ���o ��@�ѡ9 4@�0�!?����4A�@���љٿي:z ��@`�?�  4@=V�)�!?NZ��4A�@���љٿي:z ��@`�?�  4@=V�)�!?NZ��4A�@�K��Ιٿ$A3g ��@�̮� 4@�s�$�!?�O.�4A�@W��tҙٿ��[ ��@�6 4@8��@�!?�zK5A�@�N:ۙٿ���@ ��@'rLo 4@),��!?�$5A�@�N:ۙٿ���@ ��@'rLo 4@),��!?�$5A�@�N:ۙٿ���@ ��@'rLo 4@),��!?�$5A�@�,}�ԙٿ��wX ��@[b� 4@OYP�t�!?x1X5A�@t�>�֙ٿ��%Y ��@(P�� 4@A'��a�!?�=r5A�@t�>�֙ٿ��%Y ��@(P�� 4@A'��a�!?�=r5A�@t�>�֙ٿ��%Y ��@(P�� 4@A'��a�!?�=r5A�@t�>�֙ٿ��%Y ��@(P�� 4@A'��a�!?�=r5A�@t�>�֙ٿ��%Y ��@(P�� 4@A'��a�!?�=r5A�@<T�X֙ٿ�B�[ ��@�e�� 4@��ԥr�!?���5A�@S�p�ҙٿVx�G ��@�yfP 4@"�{u�!?���$5A�@Y���әٿ��R ��@�a!� 4@ʧ���!?���5A�@���ՙٿ!R\ ��@옯� 4@Wc�!?'à5A�@@7�әٿK�T ��@�"�7 4@lS�.�!?�;/5A�@����Ǚٿ���9 ��@�oʹ 4@�F�a�!?oHz5A�@��{Ιٿ��	9 ��@��2 4@�EJ!�!?{�75A�@s�W;͙ٿZ��< ��@��t� 4@��(5�!?�|$5A�@�a�3יٿO��0 ��@r!${ 4@���f�!?x؆;5A�@�>Mۙٿ;w* ��@1�X
 4@8"r�o�!?���R5A�@3D@8�ٿ"{ ��@�_= 4@EI�!?��m5A�@3D@8�ٿ"{ ��@�_= 4@EI�!?��m5A�@3D@8�ٿ"{ ��@�_= 4@EI�!?��m5A�@3D@8�ٿ"{ ��@�_= 4@EI�!?��m5A�@3D@8�ٿ"{ ��@�_= 4@EI�!?��m5A�@�F�יٿO�#, ��@�� 4@ֿL�Z�!?G�<5A�@l9��ՙٿ�x�- ��@�u�� 4@�uhd�!?�4Z$5A�@qm;
ݙٿzT ��@���! 4@��yX�!?fA�R5A�@���ٙٿ*� ��@M�^
 4@��bh�!?W�M5A�@���ٙٿ*� ��@M�^
 4@��bh�!?W�M5A�@�P�Kҙٿ��� ��@�Ҹ� 4@�u��
�!?�W@5A�@����יٿ�݂ ��@�z� 4@�t~�Q�!?��m5A�@S0�ٿ/�����@��=l 4@`O�'A�!?����5A�@Gn��ٿo&�����@֗nq 4@�ҕ��!?ϓU�5A�@O�m��ٿT����@+��� 4@�k���!?�9~�5A�@�g�ٿD������@�]� 4@�r��\�!?T�4�5A�@�bR��ٿ�R�����@nMA 4@��s�!?��n�5A�@��PI�ٿ��	 ��@�dx� 4@�T�A�!?���5A�@��PI�ٿ��	 ��@�dx� 4@�T�A�!?���5A�@(o����ٿp<< ��@o�TM 4@�19?�!?�LH�5A�@d�RH�ٿ7ߑ7 ��@���� 4@W�Kz�!?�L�`5A�@���y�ٿi�%T ��@��
 4@+�eG�!?5�P@5A�@+���ٿ'_) ��@
x� 4@����]�!?2���5A�@=8ȋ��ٿ��� ��@��� 4@\C�V�!?xύ5A�@n�h��ٿ��� ��@�q� 4@û�Na�!?\�o5A�@2j���ٿ8k����@f�hu 4@]Af�!?Hp��5A�@ �����ٿ�� ��@�{1� 4@�(:�o�!?�T�5A�@�<���ٿ�0� ��@Ζ� 4@A��i�!?-P�Y5A�@���ٿ밙' ��@ x�y 4@ ,�)��!?���L5A�@5G�tޙٿE$J ��@w�h" 4@�Icȍ�!?� �5A�@5G�tޙٿE$J ��@w�h" 4@�Icȍ�!?� �5A�@@;s�ܙٿ�G�S ��@P� 4@5��S��!?k69	5A�@��Nϙٿ�jک ��@�r���3@����U�!?R�4A�@O���֙ٿ�ƒ ��@�v���3@�fiLH�!?����4A�@��Ɵęٿ�� ��@gG���3@̀d,A�!?�?Z<4A�@��J��ٿrͰ� ��@�
Z5��3@�;�+R�!?�^64A�@�3Yߙٿ]�@� ��@7\'� 4@tؼWQ�!?�k��4A�@���i��ٿ�|h ��@�Ȉ�
 4@",���!?�H�*5A�@�{�Eٙٿ;=�[ ��@�k:� 4@$\�!?�fo5A�@��~ϙٿ���j ��@�zȪ  4@��'C�!?��6�4A�@8
gϙٿ��>� ��@)�0w��3@f���!?���4A�@	 �۹�ٿa� ��@P!>���3@	�09�!?4W4�4A�@D�ؙٿ�~�N ��@�ު� 4@�:�!?��5A�@D�ؙٿ�~�N ��@�ު� 4@�:�!?��5A�@~�Y�ٿpZ{ ��@u��� 4@d�i�!?�͸_5A�@�#���ٿ?�| ��@�Y�� 4@+��[я!?����4A�@�#���ٿ?�| ��@�Y�� 4@+��[я!?����4A�@�%����ٿ��� ��@��� 4@gi� �!?CO�5A�@�%����ٿ��� ��@��� 4@gi� �!?CO�5A�@�%����ٿ��� ��@��� 4@gi� �!?CO�5A�@�%����ٿ��� ��@��� 4@gi� �!?CO�5A�@����ٿ	|P����@q� 4@��-�!?k�B6A�@Q�NZ"�ٿW	�C���@����- 4@�y1)7�!?&r�6A�@Q�NZ"�ٿW	�C���@����- 4@�y1)7�!?&r�6A�@�l(��ٿ�f�����@C�R�" 4@U�?;P�!?om�g6A�@Ny$��ٿ�+W���@F�t* 4@v�R�!?�%��6A�@Ny$��ٿ�+W���@F�t* 4@v�R�!?�%��6A�@�q���ٿ+@v���@Q�˫% 4@���$�!?*v;�6A�@�q���ٿ+@v���@Q�˫% 4@���$�!?*v;�6A�@����ٿ9��4���@U�- 4@�VM�$�!?"��6A�@$�� �ٿ�K)���@@���0 4@��RV=�!?��7A�@te�ٿ =����@D��O6 4@3��S�!?�J\7A�@-�ƚ�ٿ-�Zo���@0�S� 4@���_�!?�BF6A�@����ٿ�����@l��� 4@%�s��!?�$D�5A�@<zc�ٿ�v�o���@��;O 4@�XQ��!?�n�6A�@@�9��ٿ�;�����@�4- 4@�(C'}�!?@�6A�@@�9��ٿ�;�����@�4- 4@�(C'}�!?@�6A�@�tct��ٿġ����@®C 4@���
H�!?E�"�5A�@Q����ٿ�U����@9�H�. 4@��1�:�!?&U�6A�@K�N�B�ٿ������@^���M 4@p[��K�!?Xh58A�@�	��4�ٿ������@���-Q 4@��>�d�!?�]�b8A�@�	��4�ٿ������@���-Q 4@��>�d�!?�]�b8A�@��A��ٿ�#�����@��â2 4@�O�c�!?�E�6A�@��A��ٿ�#�����@��â2 4@�O�c�!?�E�6A�@�AS15�ٿ]�D���@u�7K 4@��X�!?��N8A�@����4�ٿ-�R���@��_G 4@m��3%�!?��b�7A�@�	�ٿ��E����@����1 4@�(�C�!?���6A�@�	�ٿ��E����@����1 4@�(�C�!?���6A�@��K��ٿH�J����@��
8 4@�����!?���=7A�@���1��ٿ��e����@���/ 4@Ê
gm�!?���6A�@���1��ٿ��e����@���/ 4@Ê
gm�!?���6A�@���1��ٿ��e����@���/ 4@Ê
gm�!?���6A�@=���ٿ�3�����@�^�( 4@�P�9z�!?�bD6A�@?J�k��ٿ׸� ��@f!��3@9z+dF�!?џ:�4A�@?J�k��ٿ׸� ��@f!��3@9z+dF�!?џ:�4A�@?J�k��ٿ׸� ��@f!��3@9z+dF�!?џ:�4A�@�����ٿf��`��@(F*���3@'M�&T�!?4��3A�@_8#��ٿ��= ��@���j��3@�C=�K�!?�e��4A�@uPB���ٿ\3��@��}(��3@���!?S\��3A�@r�ncg�ٿ	L���@8����3@�����!?I��F2A�@��!��ٿ�	fD��@ ?x��3@����b�!?���73A�@%�Q>�ٿ��/��@ B�ٶ�3@ ND�J�!?֕g�1A�@%�Q>�ٿ��/��@ B�ٶ�3@ ND�J�!?֕g�1A�@�oK���ٿ��q���@ζ[� 4@���F�!?���G5A�@V3~�ݙٿa�����@Kr�4 4@�'�s3�!?2�Q�5A�@x�c��ٿ�3����@��޶ 4@�u<�!?#��6A�@���y+�ٿ��r����@�� ; 4@\	
�p�!?V�q`7A�@s��e�ٿ~�����@ݮS�] 4@ȓk̅�!? �c�8A�@��)��ٿ�7[����@r��b 4@��Վ�!?��&9A�@Ȝms��ٿ�c
/���@���]� 4@1_�TS�!?�
l�<A�@Ȝms��ٿ�c
/���@���]� 4@1_�TS�!?�
l�<A�@m\?�ٛٿ�F����@�!��34@-ц�N�!?��bBA�@��y(�ٿ�:
���@��hg4@�rP�4�!?���cDA�@�O:!�ٿ�0����@GYs� 4@��S��!?��=A�@��7J�ٿ[H�^���@&PM�� 4@6B�*�!?^>�T?A�@3~�}��ٿ�\V���@�M>�� 4@`y�1�!?�4A><A�@�@�UV�ٿ�����@�B�4@�E�^�!?��AA�@Q��ٿ�ݤ����@�a�!� 4@��d�!?F��>A�@bV�7�ٿ��(���@	�4@�^
u�!?����HA�@bV�7�ٿ��(���@	�4@�^
u�!?����HA�@羇�8�ٿ$�)~��@��o�4@K�	�f�!?u��bQA�@羇�8�ٿ$�)~��@��o�4@K�	�f�!?u��bQA�@��+�ٿG�����@�22��4@@�钐!?���IA�@��W42�ٿ�1�,���@����� 4@����'�!?��|�:A�@�l�i4�ٿ=`����@*p�4@�+nm�!?�te�KA�@�l�i4�ٿ=`����@*p�4@�+nm�!?�te�KA�@�ЪO��ٿ=?�x��@}ɐHv4@l_�|�!?�>?/PA�@�ЪO��ٿ=?�x��@}ɐHv4@l_�|�!?�>?/PA�@�ЪO��ٿ=?�x��@}ɐHv4@l_�|�!?�>?/PA�@�]n̾�ٿ�����@k/� 4@O��1�!?OJ3d?A�@�]n̾�ٿ�����@k/� 4@O��1�!?OJ3d?A�@J%毛ٿ麒,��@JZ��4@�?�{�!?s��FA�@J%毛ٿ麒,��@JZ��4@�?�{�!?s��FA�@�v�ٿ�������@;p!i 4@��Ń}�!?xe�6A�@�v�ٿ�������@;p!i 4@��Ń}�!?xe�6A�@���f�ٿ��d���@��˥�4@Шe�@�!?�ƍ�UA�@ĿZ>ۜٿ�֦��@����4@̸�Ė�!?<5UA�@��d�ٿ�i��@��4@��쒛�!?�K�DWA�@��d�ٿ�i��@��4@��쒛�!?�K�DWA�@&p^�Ӟٿ
�VH҇�@=��
4@�A{6Z�!?/ �nA�@&p^�Ӟٿ
�VH҇�@=��
4@�A{6Z�!?/ �nA�@ Qm,�ٿb�ڄԇ�@xsl�4@��[�>�!?פ��jA�@ Qm,�ٿb�ڄԇ�@xsl�4@��[�>�!?פ��jA�@�ElU��ٿ(1��݇�@�1��4@��'�\�!?�^��`A�@�ElU��ٿ(1��݇�@�1��4@��'�\�!?�^��`A�@$	����ٿ�4f�؇�@t( �G4@��� V�!?����eA�@'xA�V�ٿ����Ї�@�BbQ4@�~5V�!?�,YQqA�@��2�ٿ����@	�̶�4@3���t�!?ױ��HA�@��2�ٿ����@	�̶�4@3���t�!?ױ��HA�@��2�ٿ����@	�̶�4@3���t�!?ױ��HA�@�Cs(o�ٿ=��N���@�#� �4@�#��|�!?�0�EA�@�DuT�ٿ��8B��@��?b��3@q�cِ!?����A�@�DuT�ٿ��8B��@��?b��3@q�cِ!?����A�@�DuT�ٿ��8B��@��?b��3@q�cِ!?����A�@�t1ږٿ��"!��@8�[ӆ�3@Q?�!?�G�~A�@�t1ږٿ��"!��@8�[ӆ�3@Q?�!?�G�~A�@��A��ٿ�.O-��@Q��B�3@�*!{�!?��z�@�@֟;��ٿ}��!��@�u7Mc�3@I5�zB�!?��yVA�@֟;��ٿ}��!��@�u7Mc�3@I5�zB�!?��yVA�@e,�3x�ٿ��]F��@Gh��C�3@h��U�!?��x A�@���d�ٿ�0�!1��@$��K��3@̠>�U�!?G�'�@�@?'Бӕٿ����)��@�d�1��3@�*�3܏!?�ZF"A�@?'Бӕٿ����)��@�d�1��3@�*�3܏!?�ZF"A�@�+��<�ٿn<��B��@74����3@<gW��!?-��L�@�@�٭UΛٿ����@@��v4@/�?w��!?��JCA�@�٭UΛٿ����@@��v4@/�?w��!?��JCA�@�٭UΛٿ����@@��v4@/�?w��!?��JCA�@�٭UΛٿ����@@��v4@/�?w��!?��JCA�@��3�ٿy,xP��@�B`d4@H�P6Ő!?�:�LA�@�
��e�ٿ��ތ��@��.z��3@��	ː!?#אq+A�@.[��ٿ��K
��@������3@��-j�!?"�7�'A�@Lb�)�ٿoF��@,�\� 4@����!?�o�M5A�@Lb�)�ٿoF��@,�\� 4@����!?�o�M5A�@Lb�)�ٿoF��@,�\� 4@����!?�o�M5A�@�f�E�ٿ9��ۇ�@96�@g4@����]�!?"��7hA�@�f�E�ٿ9��ۇ�@96�@g4@����]�!?"��7hA�@�f�E�ٿ9��ۇ�@96�@g4@����]�!?"��7hA�@�f�E�ٿ9��ۇ�@96�@g4@����]�!?"��7hA�@�f�E�ٿ9��ۇ�@96�@g4@����]�!?"��7hA�@�O���ٿd�I�߇�@]_YW4@�,y̜�!?ټneA�@�O���ٿd�I�߇�@]_YW4@�,y̜�!?ټneA�@'8|���ٿQ����@��~� 4@�m�א!?�Ϧ�;A�@'8|���ٿQ����@��~� 4@�m�א!?�Ϧ�;A�@'8|���ٿQ����@��~� 4@�m�א!?�Ϧ�;A�@'8|���ٿQ����@��~� 4@�m�א!?�Ϧ�;A�@�L��l�ٿ�{��0��@z�Ys>�3@=��'��!?�V ��@�@�L��l�ٿ�{��0��@z�Ys>�3@=��'��!?�V ��@�@�-G7��ٿ���0��@��&!�3@�<`��!?+����@�@�-G7��ٿ���0��@��&!�3@�<`��!?+����@�@����G�ٿ����@���ӌ4@�S�a�!?�)TA�@����G�ٿ����@���ӌ4@�S�a�!?�)TA�@v�?A�ٿ�й��@�w��) 4@�N��'�!?Q��w7A�@v�?A�ٿ�й��@�w��) 4@�N��'�!?Q��w7A�@v�?A�ٿ�й��@�w��) 4@�N��'�!?Q��w7A�@�+��	�ٿ\��ʄ��@
�u6�3@�T�� �!?wg�@�@���!2�ٿ��q���@9�dd��3@���`�!?�9>�}@�@`R���ٿ(
�|��@�*���3@{�A`u�!? :�@�@`R���ٿ(
�|��@�*���3@{�A`u�!? :�@�@d1��g�ٿE�/QЈ�@�����3@�7f[Z�!?�H%Om@�@���H�ٿ���ֈ�@��	hr�3@�?Lܮ�!?GR�$i@�@gC�ٿ ,6=W��@%�'?�3@q��G�!?�;���?�@.�ς�ٿ'�d�e��@uY��3@�I]�!�!?dF���?�@��;�2�ٿ9z��@�;@��3@��w��!?]l�9@�@��;�2�ٿ9z��@�;@��3@��w��!?]l�9@�@��;�2�ٿ9z��@�;@��3@��w��!?]l�9@�@�N��3�ٿ��m��@�gmd�3@zֲ�'�!?.B��S@�@�N��3�ٿ��m��@�gmd�3@zֲ�'�!?.B��S@�@�N��3�ٿ��m��@�gmd�3@zֲ�'�!?.B��S@�@����*�ٿ�\�و�@.���j�3@M�`q)�!?�h�O@�@�n�*��ٿ�)���@}�"$�3@괋E�!?�G�A�@�n�*��ٿ�)���@}�"$�3@괋E�!?�G�A�@�n�*��ٿ�)���@}�"$�3@괋E�!?�G�A�@�n�*��ٿ�)���@}�"$�3@괋E�!?�G�A�@�n�*��ٿ�)���@}�"$�3@괋E�!?�G�A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@�!at|�ٿ7)Q
ʇ�@`ak\4@]z�Qh�!?��`�]A�@}ͬ�ٿ��l(���@�'m�Q4@iY=K��!?��l]�A�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�g���ٿ 9�(��@l�}й�3@��2zd�!?P����@�@�Ѯ���ٿ��V�Q��@�Pq���3@�PL
�!?���@�@�Ѯ���ٿ��V�Q��@�Pq���3@�PL
�!?���@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�NR+�ٿt(�_:��@;s�3@����!?�h�N�@�@�!��ٿ�i�a��@��L-��3@����!?Q�"C�@�@�@�ٿ�&����@����`�3@�l@�-�!?j���@�@�@�ٿ�&����@����`�3@�l@�-�!?j���@�@�@�ٿ�&����@����`�3@�l@�-�!?j���@�@�@�ٿ�&����@����`�3@�l@�-�!?j���@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@���Փٿ(�<l^��@������3@֔ǈ4�!?I'[��@�@�3��s�ٿਬ��@Q�=�3@<��	�!?�𾙟@�@�3��s�ٿਬ��@Q�=�3@<��	�!?�𾙟@�@�3��s�ٿਬ��@Q�=�3@<��	�!?�𾙟@�@��Lڙٿ"�T���@�E�:�3@���L8�!?���Q�@�@��Lڙٿ"�T���@�E�:�3@���L8�!?���Q�@�@��Lڙٿ"�T���@�E�:�3@���L8�!?���Q�@�@��Lڙٿ"�T���@�E�:�3@���L8�!?���Q�@�@&��l�ٿr��	͇�@ �7�84@;OF%'�!?B���tA�@&��l�ٿr��	͇�@ �7�84@;OF%'�!?B���tA�@��{�i�ٿ2�b53��@�=I�3@��!?�/��A�@~V��͑ٿ���i��@2��|4@4o��!?�h_�A�@~V��͑ٿ���i��@2��|4@4o��!?�h_�A�@~V��͑ٿ���i��@2��|4@4o��!?�h_�A�@Ί�]�ٿj�4|��@��w$B�3@�4�TF�!?b��@�@�����ٿ�E����@�ʆ*f4@��Đ!?���m@A�@&���4�ٿER����@B��k^�3@"p�K.�!? ���5A�@&���4�ٿER����@B��k^�3@"p�K.�!? ���5A�@&���4�ٿER����@B��k^�3@"p�K.�!? ���5A�@&���4�ٿER����@B��k^�3@"p�K.�!? ���5A�@&���4�ٿER����@B��k^�3@"p�K.�!? ���5A�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@���ܝٿ���r��@�����3@�]u2Y�!?����@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@��L��ٿ�s?��@٢�a�3@; .�!?��[��@�@wO���ٿ���詇�@��&X�4@V��!�!?*o��A�@�Zɪ�ٿ��$�5��@���8�3@Lan��!?�l-�A�@�Zɪ�ٿ��$�5��@���8�3@Lan��!?�l-�A�@�Zɪ�ٿ��$�5��@���8�3@Lan��!?�l-�A�@*G9��ٿj'����@2a�A�3@��89 �!?j�m>$A�@*G9��ٿj'����@2a�A�3@��89 �!?j�m>$A�@*G9��ٿj'����@2a�A�3@��89 �!?j�m>$A�@*G9��ٿj'����@2a�A�3@��89 �!?j�m>$A�@��S�ٙٿu8�R��@��W���3@mɤ�,�!?Z�b��@�@��S�ٙٿu8�R��@��W���3@mɤ�,�!?Z�b��@�@��S�ٙٿu8�R��@��W���3@mɤ�,�!?Z�b��@�@ӭ�>�ٿ{u�&��@ �#)��3@�B�!?��|A�@ӭ�>�ٿ{u�&��@ �#)��3@�B�!?��|A�@ӭ�>�ٿ{u�&��@ �#)��3@�B�!?��|A�@ӭ�>�ٿ{u�&��@ �#)��3@�B�!?��|A�@Eu��&�ٿ�	��@cz�C 4@�m�-�!?	ni�A�@�����ٿ��Y���@�}�M� 4@+v<3�!?&RA�@�����ٿ��Y���@�}�M� 4@+v<3�!?&RA�@�����ٿ��Y���@�}�M� 4@+v<3�!?&RA�@�����ٿ��Y���@�}�M� 4@+v<3�!?&RA�@�2F��ٿK�wc���@%"4��4@��|#�!?;0HAA�@�2F��ٿK�wc���@%"4��4@��|#�!?;0HAA�@�2F��ٿK�wc���@%"4��4@��|#�!?;0HAA�@�2F��ٿK�wc���@%"4��4@��|#�!?;0HAA�@��ރ˕ٿ������@hƴ~^
4@�F���!?J�i�A�@��ރ˕ٿ������@hƴ~^
4@�F���!?J�i�A�@�[ʱ�ٿ%��=��@�yS7b�3@�Jۤ��!?�����@�@�[ʱ�ٿ%��=��@�yS7b�3@�Jۤ��!?�����@�@�[ʱ�ٿ%��=��@�yS7b�3@�Jۤ��!?�����@�@.�`)��ٿ�왽���@W�244@u��A��!?�� �A�@.�`)��ٿ�왽���@W�244@u��A��!?�� �A�@.�`)��ٿ�왽���@W�244@u��A��!?�� �A�@.�`)��ٿ�왽���@W�244@u��A��!?�� �A�@.�`)��ٿ�왽���@W�244@u��A��!?�� �A�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@�l���ٿ�$ ?���@N�R�3@~(�/��!?�����@�@N&]��ٿ�վ7��@S]����3@��@t�!?TE�*@�@N&]��ٿ�վ7��@S]����3@��@t�!?TE�*@�@N&]��ٿ�վ7��@S]����3@��@t�!?TE�*@�@��J�o�ٿ�!Έa��@��}E�3@�g�!?��5��@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@ 5����ٿ�j<�׈�@U�� �3@�I�U�!?��M@�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@]�4ʒٿ�����@�o�Q 4@u�#=v�!?����PA�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@�Ņ�5�ٿ�dCe��@����^�3@�
�j�!?�xJ�@�@%���5�ٿ�i���@�@�4��3@�u?h�!?@/Qm
A�@N�km�ٿ$��§��@����4@��x�8�!?J���xA�@N�km�ٿ$��§��@����4@��x�8�!?J���xA�@��F�ٿ��?�Ԉ�@<����3@>=m�)�!?���y@�@��F�ٿ��?�Ԉ�@<����3@>=m�)�!?���y@�@��F�ٿ��?�Ԉ�@<����3@>=m�)�!?���y@�@SW2I�ٿj��RB��@[eٻ�3@����!?�k�T�@�@SW2I�ٿj��RB��@[eٻ�3@����!?�k�T�@�@SW2I�ٿj��RB��@[eٻ�3@����!?�k�T�@�@ [e�1�ٿ�a��
��@�^q��3@�2����!?x��&A�@ [e�1�ٿ�a��
��@�^q��3@�2����!?x��&A�@ [e�1�ٿ�a��
��@�^q��3@�2����!?x��&A�@ [e�1�ٿ�a��
��@�^q��3@�2����!?x��&A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@���PS�ٿ��j_��@~)�M �3@��\���!?����A�@� A��ٿyǂ����@;zz�4@R}���!?�<x�A�@� A��ٿyǂ����@;zz�4@R}���!?�<x�A�@.���L�ٿW�bˈ�@{�m��3@��!?~3�,A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@sִ>��ٿg�����@�,T�)�3@�D̺�!?��gW�A�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@��H�E�ٿW1趹��@��� ��3@|y���!?[���qA�@RG�:��ٿ����@нqc�3@�>Y�!?% c�A�@RG�:��ٿ����@нqc�3@�>Y�!?% c�A�@RG�:��ٿ����@нqc�3@�>Y�!?% c�A�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@�f��g�ٿHŲY��@1|X9t�3@Z��V�!?�z�Z7@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@e�m��ٿ}�iUm��@32�_H4@ӥ^��!?r�Hv<@�@�{�l�ٿ�!d� ��@y��3@��_e�!?��ШA�@�{�l�ٿ�!d� ��@y��3@��_e�!?��ШA�@�{�l�ٿ�!d� ��@y��3@��_e�!?��ШA�@�{�l�ٿ�!d� ��@y��3@��_e�!?��ШA�@!H�)�ٿG�����@^����3@$��/�!?�k�,B�@!H�)�ٿG�����@^����3@$��/�!?�k�,B�@!H�)�ٿG�����@^����3@$��/�!?�k�,B�@�8Ğ�ٿe�6	���@
��i��3@O�y�!?%�	c�B�@�8Ğ�ٿe�6	���@
��i��3@O�y�!?%�	c�B�@�8Ğ�ٿe�6	���@
��i��3@O�y�!?%�	c�B�@H�d��ٿ���5��@M��3@pQT��!?P��A�@N����ٿ�kìY��@@-ܸ��3@3��}�!?EXMA�@N����ٿ�kìY��@@-ܸ��3@3��}�!?EXMA�@N����ٿ�kìY��@@-ܸ��3@3��}�!?EXMA�@N����ٿ�kìY��@@-ܸ��3@3��}�!?EXMA�@]"F��ٿ��̿��@�%G��3@%�; �!?O����A�@]"F��ٿ��̿��@�%G��3@%�; �!?O����A�@]"F��ٿ��̿��@�%G��3@%�; �!?O����A�@��`:�ٿ^%����@ N���3@W�`$�!?�5�2A�@��`:�ٿ^%����@ N���3@W�`$�!?�5�2A�@��`:�ٿ^%����@ N���3@W�`$�!?�5�2A�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@�g�+�ٿ3dԔ��@,/�Ÿ�3@�Mkݏ!?1~|T�@�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@����ٿ�d g@��@��m���3@Č�2��!?Ә˕"A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@mB�Si�ٿχ,�k��@B�q���3@W'�U�!?ӻ��A�@�3�ٿ��8���@AΧ�4@/�x?�!?�O߿A�@�3�ٿ��8���@AΧ�4@/�x?�!?�O߿A�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@R�֑��ٿ�.6�܇�@nt���3@����!?[-�ڂ@�@�/��ٿ���v��@��:*��3@?Mn�!?�fCA�@�/��ٿ���v��@��:*��3@?Mn�!?�fCA�@�/��ٿ���v��@��:*��3@?Mn�!?�fCA�@im*�R�ٿK����@*.Q� 4@��	�f�!?��N'@�@im*�R�ٿK����@*.Q� 4@��	�f�!?��N'@�@�*I���ٿ��<G0��@?�j	4@�s�
�!?��:��>�@�g(gߞٿoI ����@�m�4@K����!?,�/�?�@�qT��ٿ��7����@�����4@a�)c�!?w�ʯl?�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@ʝ�|��ٿZ�M�{��@�F �x�3@;wc�!?$V �fA�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@���|�ٿ�=�X��@�"�D�3@��݅�!?�mK&�@�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@�s�5�ٿ]�5���@�W�ч�3@�J��!?O;i��?�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@���6��ٿl:��@燰���3@�Z<�!?�A��N@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@��ʓ�ٿ��*�W��@�fG��3@F�dP�!?с�d@�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@="�^�ٿ-��Q��@�����3@��p��!?<U;A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@5�����ٿ}p��n��@���W�3@<�j�!?���~(A�@�og�љٿ!4>���@�Y����3@�κ4�!?� ���@�@�og�љٿ!4>���@�Y����3@�κ4�!?� ���@�@�og�љٿ!4>���@�Y����3@�κ4�!?� ���@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@�� ��ٿ�}�=��@psO�|�3@��A�!?�=~hM@�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@mgM��ٿ���&��@���z�3@1�j�n�!?��)A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@�0��K�ٿ�+�z|��@d����3@#pZ��!?�[��7A�@��ZN:�ٿC���s��@*�'�X�3@эbcW�!?�u��S@�@[\��y�ٿ�x�2��@�����3@�oq�!?زՉ�?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@܅凌�ٿ^�dy��@h�)�-�3@��6(�!?���K?�@DaM]��ٿ�Lli���@F���5�3@'���a�!?>��u�?�@-Ԥe^�ٿ�$ U��@�Z��3@g��6P�!?zK4�>�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@�댚�ٿ˗�/���@K��_��3@�bR'�!?~?�@�@,m��f�ٿ_��[���@�����4@�\H]��!?��Z@�@r3%��ٿ1w� ��@�BH���3@���q/�!?6e��%@�@r3%��ٿ1w� ��@�BH���3@���q/�!?6e��%@�@r3%��ٿ1w� ��@�BH���3@���q/�!?6e��%@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@B����ٿ��#��@+8ql�3@��R�!?���@�@d:���ٿ�`I�#��@+�ߴ\�3@�~�^\�!?	��'A�@d:���ٿ�`I�#��@+�ߴ\�3@�~�^\�!?	��'A�@c�a�ٿH���\��@��,4h�3@����!?�ʘ1@�@c�a�ٿH���\��@��,4h�3@����!?�ʘ1@�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@[�2V1�ٿ�C��4��@�Q@��3@�4�WI�!?��C�A�@�-�A��ٿr�	����@�*@4@�a��}�!?�B�'A�@�-�A��ٿr�	����@�*@4@�a��}�!?�B�'A�@�0@��ٿϔYl��@1դ��4@�d"\�!?�;x�}A�@�{���ٿm��<��@J�:���3@�_�b�!?W,��A�@�Ѧ���ٿ흰�)��@�&���3@��q���!?�1��2A�@#�S��ٿ���a���@=�3_s�3@�W�q�!?\����?�@�*�`��ٿ6�+I��@��.J�3@�u>a�!?�X��?�@,��6A�ٿ$�E<��@H�V9��3@Lf��F�!?��V�.?�@,��6A�ٿ$�E<��@H�V9��3@Lf��F�!?��V�.?�@,��6A�ٿ$�E<��@H�V9��3@Lf��F�!?��V�.?�@,��6A�ٿ$�E<��@H�V9��3@Lf��F�!?��V�.?�@3�ND�ٿ`0����@�ԧ���3@s鰸H�!?e�i\>�@3�ND�ٿ`0����@�ԧ���3@s鰸H�!?e�i\>�@3�ND�ٿ`0����@�ԧ���3@s鰸H�!?e�i\>�@\��l��ٿ��L 4��@0�9ڼ�3@��8[�!?��`B�=�@\��l��ٿ��L 4��@0�9ڼ�3@��8[�!?��`B�=�@^��Ғٿ�f�8
��@�:Q7�3@h��.�!?CD�">>�@^��Ғٿ�f�8
��@�:Q7�3@h��.�!?CD�">>�@^��Ғٿ�f�8
��@�:Q7�3@h��.�!?CD�">>�@�;���ٿ�b��@_&�B��3@�--�!?�b�<�@c4�Ꚑٿ+@$�(��@)0�W4@j��8�!?��]�;�@c4�Ꚑٿ+@$�(��@)0�W4@j��8�!?��]�;�@s-���ٿwcH����@7���V�3@^4�:B�!?��A:�@�R�q�ٿ�Ma���@F+(��3@j��j�!?�v�9�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ��A���@$A�͜ 4@���
�!?��yS5�@����ٿ�5u��@�� o��3@XBN �!?3Q[6<�@����ٿ�5u��@�� o��3@XBN �!?3Q[6<�@����ٿ�5u��@�� o��3@XBN �!?3Q[6<�@\K��ٿӧ����@'����3@�4<F�!?yc9K;�@\K��ٿӧ����@'����3@�4<F�!?yc9K;�@\K��ٿӧ����@'����3@�4<F�!?yc9K;�@\K��ٿӧ����@'����3@�4<F�!?yc9K;�@\K��ٿӧ����@'����3@�4<F�!?yc9K;�@�ޤ�`�ٿ��j<��@�1�P��3@�2�S�!?/��=4�@�ޤ�`�ٿ��j<��@�1�P��3@�2�S�!?/��=4�@�ޤ�`�ٿ��j<��@�1�P��3@�2�S�!?/��=4�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@؟��i�ٿTB���@t'}oK4@��d��!?��� �<�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���!;�ٿ�6�,P��@��U͓4@ �_(�!? Uoz:�@���ik�ٿ�c�n��@��\��3@�H�N?�!?�wA��;�@���ik�ٿ�c�n��@��\��3@�H�N?�!?�wA��;�@���	[�ٿ��u;��@�f�9^4@nD4IA�!?H
f=�@���	[�ٿ��u;��@�f�9^4@nD4IA�!?H
f=�@\�����ٿJ����@`�[-�3@���Xr�!?'bV�,�@\�����ٿJ����@`�[-�3@���Xr�!?'bV�,�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@)�'��ٿ���`��@�{<[��3@�
L�J�!?3�w'�@��E��ٿ��Լz��@�HL�3@�о^U�!?H��U��@n4(���ٿPig���@�vD*��3@�?W��!?zSg�@n4(���ٿPig���@�vD*��3@�?W��!?zSg�@�h�N�ٿW�&΂�@Oq��K4@�h=l��!?$�;t��@�h�N�ٿW�&΂�@Oq��K4@�h=l��!?$�;t��@�h�N�ٿW�&΂�@Oq��K4@�h=l��!?$�;t��@�h�N�ٿW�&΂�@Oq��K4@�h=l��!?$�;t��@>�%��ٿ��ؼ��@1�{� 4@4��f�!?#�b�i8�@>�%��ٿ��ؼ��@1�{� 4@4��f�!?#�b�i8�@����&�ٿ��sB��@�&
y�3@0+%V3�!?*	�=2�@����&�ٿ��sB��@�&
y�3@0+%V3�!?*	�=2�@����&�ٿ��sB��@�&
y�3@0+%V3�!?*	�=2�@����&�ٿ��sB��@�&
y�3@0+%V3�!?*	�=2�@����&�ٿ��sB��@�&
y�3@0+%V3�!?*	�=2�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@Z{��ƛٿ�j���@ �G�4@ �\�s�!?���p-�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@����b�ٿ�02C]��@�Q��y�3@���5P�!?`���f:�@dq�~^�ٿ=Awc8��@c~U$�3@���,�!?|6�9�@dq�~^�ٿ=Awc8��@c~U$�3@���,�!?|6�9�@��1�ٿ�r����@~�*�4@�.��2�!?;~b��"�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@��r�4�ٿ�㋁�|�@�AI��4@H�bJJ�!?D�lER�@�A���ٿ���a"��@
l|?��3@֬�$�!?n��9�@�A���ٿ���a"��@
l|?��3@֬�$�!?n��9�@�A���ٿ���a"��@
l|?��3@֬�$�!?n��9�@�@u?�ٿH��~7}�@Z�˴4@P;�5Ϗ!?8�(ǥ�@W2r�ٿm�H�|�@����4@,AU�!?�݊S�۶@W2r�ٿm�H�|�@����4@,AU�!?�݊S�۶@W2r�ٿm�H�|�@����4@,AU�!?�݊S�۶@��ꨟٿ'���Gr�@2����4@��ߜ�!?�"����@KՊ��ٿ%�E+l�@^t��!4@�T)��!?ak�AQ�@�t��ٿT�Sq�@e�-�4@ ��]��!?2�B8}�@�t��ٿT�Sq�@e�-�4@ ��]��!?2�B8}�@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@սG釚ٿ2�Nf�@��*�v4@s�P���!?�����@Y�&�S�ٿ.V�q�@'���4@�WŤ�!?)s"
{�@Y�&�S�ٿ.V�q�@'���4@�WŤ�!?)s"
{�@Y�&�S�ٿ.V�q�@'���4@�WŤ�!?)s"
{�@8��E��ٿ� �ubv�@����� 4@Y��Z�!?gB�v���@8��E��ٿ� �ubv�@����� 4@Y��Z�!?gB�v���@8��E��ٿ� �ubv�@����� 4@Y��Z�!?gB�v���@8��E��ٿ� �ubv�@����� 4@Y��Z�!?gB�v���@�WJ��ٿ\�>�n�@�Ί���3@��{���!?Iۭ�da�@�WJ��ٿ\�>�n�@�Ί���3@��{���!?Iۭ�da�@z�J�ٿ��h6T�@�
8;�4@.?S0o�!?r��z�@z�J�ٿ��h6T�@�
8;�4@.?S0o�!?r��z�@z�J�ٿ��h6T�@�
8;�4@.?S0o�!?r��z�@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@OfHl�ٿ��-�lW�@J!0�3@��tU"�!?"�1����@�lLR�ٿ����Y�@�_4��3@���b�!?�VE`��@�lLR�ٿ����Y�@�_4��3@���b�!?�VE`��@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@����%�ٿ>��X�@��Z���3@i �Xb�!?��뜵@8(�	��ٿ��5�R�@�5'>�4@����!?�jo^i�@8(�	��ٿ��5�R�@�5'>�4@����!?�jo^i�@8(�	��ٿ��5�R�@�5'>�4@����!?�jo^i�@8(�	��ٿ��5�R�@�5'>�4@����!?�jo^i�@�)��F�ٿ�(���2�@���VU�3@����%�!?�"wO�@�)��F�ٿ�(���2�@���VU�3@����%�!?�"wO�@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@�{�93�ٿ��]z<�@�g54&�3@w�%�!?��;���@s�F�d�ٿ���H8�@+q6��3@Hc��!?乺���@s�F�d�ٿ���H8�@+q6��3@Hc��!?乺���@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@k�����ٿZ�\}L�@��rO;�3@��(�x�!?W�ʲ�0�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@F`��ٿ���UKL�@Fn��E�3@q���!?�T�3�@��)�ėٿI&��H�@@Ͱ��3@0��5�!?��,�@��)�ėٿI&��H�@@Ͱ��3@0��5�!?��,�@��+k�ٿ���S�@Z��5N4@M��!�!?�$WY�v�@����E�ٿ+a�?�@f?���3@&��V&�!?�.��WĴ@NSÿK�ٿi]qVE�@���4@�t����!?=�5���@NSÿK�ٿi]qVE�@���4@�t����!?=�5���@NSÿK�ٿi]qVE�@���4@�t����!?=�5���@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@�&���ٿ}�M��N�@J�R�4@g4��!?ɟh�qF�@���oQ�ٿ騱�S2�@~>��� 4@?���7�!?z'��Q�@���oQ�ٿ騱�S2�@~>��� 4@?���7�!?z'��Q�@���oQ�ٿ騱�S2�@~>��� 4@?���7�!?z'��Q�@���oQ�ٿ騱�S2�@~>��� 4@?���7�!?z'��Q�@68��I�ٿ��&f	-�@:�0��3@�Č���!?��(2l�@68��I�ٿ��&f	-�@:�0��3@�Č���!?��(2l�@�O�˖ٿf��2�@?4�\��3@r��_�!?t��h�L�@�O�˖ٿf��2�@?4�\��3@r��_�!?t��h�L�@�O�˖ٿf��2�@?4�\��3@r��_�!?t��h�L�@�O�˖ٿf��2�@?4�\��3@r��_�!?t��h�L�@�(G��ٿYщ�S�@'ã� 4@fۇ��!?.�闊w�@
��3Řٿ��7U�4�@@�����3@r�*[��!?��G�t^�@
��3Řٿ��7U�4�@@�����3@r�*[��!?��G�t^�@
��3Řٿ��7U�4�@@�����3@r�*[��!?��G�t^�@
��3Řٿ��7U�4�@@�����3@r�*[��!?��G�t^�@�z�K�ٿol�|�h�@2w��3@n�Ã9�!? �4/]'�@�z�K�ٿol�|�h�@2w��3@n�Ã9�!? �4/]'�@�z�K�ٿol�|�h�@2w��3@n�Ã9�!? �4/]'�@�z�K�ٿol�|�h�@2w��3@n�Ã9�!? �4/]'�@|s��K�ٿ��K�@Cc���3@��6��!?.*�-�!�@|s��K�ٿ��K�@Cc���3@��6��!?.*�-�!�@|s��K�ٿ��K�@Cc���3@��6��!?.*�-�!�@|s��K�ٿ��K�@Cc���3@��6��!?.*�-�!�@|s��K�ٿ��K�@Cc���3@��6��!?.*�-�!�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@��-���ٿW�M}�O�@$���3@q�m���!?��{bM�@^����ٿ����S=�@w�� ��3@,�����!?��/P���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@�G��<�ٿ�*�a�@ST)\�3@Z��!?9���@��V�
�ٿ��=HN�@-�E�
�3@sB���!?{�л`;�@��V�
�ٿ��=HN�@-�E�
�3@sB���!?{�л`;�@��V�
�ٿ��=HN�@-�E�
�3@sB���!?{�л`;�@�}�-�ٿ����p4�@S���4@=k���!?�UY'�[�@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@��ֿ�ٿ�M��;�@|8R�4@�g}(�!?�}(Ћ��@I�*9��ٿ��j�V�@7��j3�3@_;b���!?mb�w��@I�*9��ٿ��j�V�@7��j3�3@_;b���!?mb�w��@I�*9��ٿ��j�V�@7��j3�3@_;b���!?mb�w��@I�*9��ٿ��j�V�@7��j3�3@_;b���!?mb�w��@xc�q4�ٿ�_�]�P�@��e��3@.�&�|�!?I�>��O�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@�b�ٿ>k^�A�@��3��3@BGR��!?�bGҼ�@��h�ٿ���aR�@�k4P�4@���s�!?�=�"{c�@��h�ٿ���aR�@�k4P�4@���s�!?�=�"{c�@��h�ٿ���aR�@�k4P�4@���s�!?�=�"{c�@��h�ٿ���aR�@�k4P�4@���s�!?�=�"{c�@��h�ٿ���aR�@�k4P�4@���s�!?�=�"{c�@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@��R��ٿq�HX�@��Aĩ�3@=P!\�!?��W��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@2�)� �ٿp@��dJ�@�{�$��3@�J�F$�!?�	Y��@uS4 Q�ٿ��J2�T�@+3�|��3@����0�!?�ab�l�@uS4 Q�ٿ��J2�T�@+3�|��3@����0�!?�ab�l�@uS4 Q�ٿ��J2�T�@+3�|��3@����0�!?�ab�l�@uS4 Q�ٿ��J2�T�@+3�|��3@����0�!?�ab�l�@uS4 Q�ٿ��J2�T�@+3�|��3@����0�!?�ab�l�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@�=�Țٿ��O�@'��hF�3@���]^�!?�I��G�@ȶ��>�ٿ��'A�@?��	4@�~8�!?M'�a�˴@ȶ��>�ٿ��'A�@?��	4@�~8�!?M'�a�˴@ȶ��>�ٿ��'A�@?��	4@�~8�!?M'�a�˴@ȶ��>�ٿ��'A�@?��	4@�~8�!?M'�a�˴@4��ѕٿ�w-��9�@��Df4@~�,�!?0FU����@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���['�ٿ	$s�|J�@���3@TS,3�!?S?v��@���u^�ٿ'�H�@������3@Z�q�!?����d�@���u^�ٿ'�H�@������3@Z�q�!?����d�@���u^�ٿ'�H�@������3@Z�q�!?����d�@#�]�ٿ �l�E�@���S��3@�O0u�!?]���@H�Yt�ٿ����Q�@��z��4@���s��!?]C4m\�@C�1�I�ٿ=�S�rS�@�#�3@U]�N*�!?4��K�m�@C�1�I�ٿ=�S�rS�@�#�3@U]�N*�!?4��K�m�@C�1�I�ٿ=�S�rS�@�#�3@U]�N*�!?4��K�m�@C�1�I�ٿ=�S�rS�@�#�3@U]�N*�!?4��K�m�@C�1�I�ٿ=�S�rS�@�#�3@U]�N*�!?4��K�m�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@�5ڤ�ٿ��lu�K�@y?��3@rp(;�!?5���B*�@��I��ٿ��c>�@
����4@�S�.ŏ!?��9'��@��I��ٿ��c>�@
����4@�S�.ŏ!?��9'��@��I��ٿ��c>�@
����4@�S�.ŏ!?��9'��@�|�]^�ٿQB]]�Q�@��#,�4@}?�Q�!?����T�@�|�]^�ٿQB]]�Q�@��#,�4@}?�Q�!?����T�@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@R%���ٿ�ktJ�@�æ�4@4+x5�!?9���@��L�яٿn�t�kI�@?�,s�3@�̌�!?�t��ߴ@��L�яٿn�t�kI�@?�,s�3@�̌�!?�t��ߴ@�eA��ٿ��N5�@�҃!.�3@��ؓ;�!?K$F�F5�@�eA��ٿ��N5�@�҃!.�3@��ؓ;�!?K$F�F5�@�eA��ٿ��N5�@�҃!.�3@��ؓ;�!?K$F�F5�@�#���ٿ��)�=�@��o�3@�u���!?�p�E��@�#���ٿ��)�=�@��o�3@�u���!?�p�E��@�#���ٿ��)�=�@��o�3@�u���!?�p�E��@�#���ٿ��)�=�@��o�3@�u���!?�p�E��@�#���ٿ��)�=�@��o�3@�u���!?�p�E��@����ٿD�ǿ,E�@F&�U��3@���L�!?�k9w��@��+Cl�ٿ��
P�@z��?�3@���zۏ!??,�;�$�@��+Cl�ٿ��
P�@z��?�3@���zۏ!??,�;�$�@��+Cl�ٿ��
P�@z��?�3@���zۏ!??,�;�$�@��+Cl�ٿ��
P�@z��?�3@���zۏ!??,�;�$�@���ٿ����M�@��ܮD	4@���!?y6/�0�@�ݽJ�ٿ�����C�@�����3@�0K��!?�/���@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@
�6�'�ٿ}5M��e�@��.F
4@�d7�!?��U>f�@�q?b�ٿSGrc�b�@��aN��3@�:���!?O�^D�@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@�JЖГٿ�p__�@�^d�3@3�#b{�!?oT��@Ib��ٿ��'��O�@!��3@T$6P�!?ُ��d�@Ib��ٿ��'��O�@!��3@T$6P�!?ُ��d�@Ib��ٿ��'��O�@!��3@T$6P�!?ُ��d�@Ib��ٿ��'��O�@!��3@T$6P�!?ُ��d�@zЮ�R�ٿ��gW�@̉�!�3@ii��_�!?�g�uޖ�@zЮ�R�ٿ��gW�@̉�!�3@ii��_�!?�g�uޖ�@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@0��[��ٿ�a��CH�@�:r�4@�=$�5�!?�%?��@�:2�Κٿ�ߏJ�@x��p�4@eM��C�!?�Z���@�:2�Κٿ�ߏJ�@x��p�4@eM��C�!?�Z���@�:2�Κٿ�ߏJ�@x��p�4@eM��C�!?�Z���@�:2�Κٿ�ߏJ�@x��p�4@eM��C�!?�Z���@��+ɖٿ/B�x�J�@��A�:	4@�#��!?�v�� �@��+ɖٿ/B�x�J�@��A�:	4@�#��!?�v�� �@��+ɖٿ/B�x�J�@��A�:	4@�#��!?�v�� �@ŵ)���ٿ�L�{uU�@-�����3@��-~�!?X>��B�@ŵ)���ٿ�L�{uU�@-�����3@��-~�!?X>��B�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@R2�~��ٿ����SX�@ƨ��3@�T$;Q�!?�h!;�Y�@�����ٿ��g=�@L����3@% �!?�
J��(�@�����ٿ��g=�@L����3@% �!?�
J��(�@�����ٿ��g=�@L����3@% �!?�
J��(�@�����ٿ��g=�@L����3@% �!?�
J��(�@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@���QҗٿN����B�@�l}$��3@��m��!?>��'���@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@�V���ٿ��G,�O�@�7ͥ4@pz(<я!?l�i�0�@`�]�@�ٿ,\ʹ@R�@�8 4@):�!?���wM�@`�]�@�ٿ,\ʹ@R�@�8 4@):�!?���wM�@`�]�@�ٿ,\ʹ@R�@�8 4@):�!?���wM�@`�]�@�ٿ,\ʹ@R�@�8 4@):�!?���wM�@`�]�@�ٿ,\ʹ@R�@�8 4@):�!?���wM�@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@6�>�(�ٿޓ%�G�@��h��3@���~�!?��<I!Ǵ@l�3�O�ٿ��fI�@J���3@4D�	�!?@�F���@l�3�O�ٿ��fI�@J���3@4D�	�!?@�F���@l�3�O�ٿ��fI�@J���3@4D�	�!?@�F���@�!�ʓٿ6z��_�@�p��3@���=�!?����@��@�!�ʓٿ6z��_�@�p��3@���=�!?����@��@�=9���ٿ��|}TO�@�kI�3@*��p%�!?��4��@k��߹�ٿ`�/�K�@~�n@��3@��!?�ܼGV´@k��߹�ٿ`�/�K�@~�n@��3@��!?�ܼGV´@y���ӘٿF��mO�@L|3��3@攔]K�!?\�~���@y���ӘٿF��mO�@L|3��3@攔]K�!?\�~���@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@־Aз�ٿ6�e�Q�@��
�q4@���z�!?��V�2!�@R����ٿZ��ozN�@�
��4@���%��!?�y�����@�Z��ٿ��+�N�@�2�T�3@*�$5�!?j�Q�_-�@�Z��ٿ��+�N�@�2�T�3@*�$5�!?j�Q�_-�@����ٿ�4�z�J�@��#�3@t�ֵr�!?��;��@����ٿ�4�z�J�@��#�3@t�ֵr�!?��;��@����ٿ�4�z�J�@��#�3@t�ֵr�!?��;��@�g��Ǔٿ���لj�@�����3@�pO���!?l�x5�@8F���ٿ��=��h�@q�z�!�3@t���S�!?�e2���@8F���ٿ��=��h�@q�z�!�3@t���S�!?�e2���@8F���ٿ��=��h�@q�z�!�3@t���S�!?�e2���@;��9:�ٿP�<�X�@؏ʾY�3@x/AU�!?w<M�i�@;��9:�ٿP�<�X�@؏ʾY�3@x/AU�!?w<M�i�@;��9:�ٿP�<�X�@؏ʾY�3@x/AU�!?w<M�i�@;��9:�ٿP�<�X�@؏ʾY�3@x/AU�!?w<M�i�@6��Lh�ٿm�]�@t0�2��3@��l�!?��09+i�@6��Lh�ٿm�]�@t0�2��3@��l�!?��09+i�@6��Lh�ٿm�]�@t0�2��3@��l�!?��09+i�@6��Lh�ٿm�]�@t0�2��3@��l�!?��09+i�@AW^�ٿ�4��|c�@L�7��3@�6q��!?�*x���@AW^�ٿ�4��|c�@L�7��3@�6q��!?�*x���@n�x.��ٿY=��O[�@���0�3@V?0�*�!?�Z���7�@n�x.��ٿY=��O[�@���0�3@V?0�*�!?�Z���7�@n�x.��ٿY=��O[�@���0�3@V?0�*�!?�Z���7�@=kSj�ٿ)�'U�b�@-"���3@v �-l�!?#Xu��H�@=kSj�ٿ)�'U�b�@-"���3@v �-l�!?#Xu��H�@=kSj�ٿ)�'U�b�@-"���3@v �-l�!?#Xu��H�@=kSj�ٿ)�'U�b�@-"���3@v �-l�!?#Xu��H�@=kSj�ٿ)�'U�b�@-"���3@v �-l�!?#Xu��H�@���i6�ٿ�c3��_�@����4@)�j$]�!?�Ǒg�@���i6�ٿ�c3��_�@����4@)�j$]�!?�Ǒg�@���i6�ٿ�c3��_�@����4@)�j$]�!?�Ǒg�@���i6�ٿ�c3��_�@����4@)�j$]�!?�Ǒg�@���i6�ٿ�c3��_�@����4@)�j$]�!?�Ǒg�@�2���ٿbп�Z\�@����Y�3@��!�!?剭U䚵@�2���ٿbп�Z\�@����Y�3@��!�!?剭U䚵@�2���ٿbп�Z\�@����Y�3@��!�!?剭U䚵@�2���ٿbп�Z\�@����Y�3@��!�!?剭U䚵@�2���ٿbп�Z\�@����Y�3@��!�!?剭U䚵@�mzd��ٿOP>,�]�@`�bv�	4@b��k�!?���se�@�mzd��ٿOP>,�]�@`�bv�	4@b��k�!?���se�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@Rn(]�ٿ���V�@�qS���3@z
�*�!?Yw��yK�@�G�oB�ٿ����{C�@�6� W�3@iB-�&�!?gљ�w��@�G�oB�ٿ����{C�@�6� W�3@iB-�&�!?gљ�w��@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@���^ԛٿ��V7H�@)��='�3@򺓛�!?1�	T^޴@�G ˟ٿ2�$�O�@���K�3@*�!�!?�/L�5��@?�g�ћٿQ���G�@ok%��3@���L�!?�	hO���@?�g�ћٿQ���G�@ok%��3@���L�!?�	hO���@7λTB�ٿ扮�RC�@9��@H�3@��W�!?��"'!�@CcAR@�ٿ1dS�O�@-��E��3@;Ř`!�!?p�r�٫�@W,��H�ٿo�Q|�7�@�Sb>��3@��3�w�!?.e�J_�@W,��H�ٿo�Q|�7�@�Sb>��3@��3�w�!?.e�J_�@W,��H�ٿo�Q|�7�@�Sb>��3@��3�w�!?.e�J_�@W,��H�ٿo�Q|�7�@�Sb>��3@��3�w�!?.e�J_�@W,��H�ٿo�Q|�7�@�Sb>��3@��3�w�!?.e�J_�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@Y_���ٿGb�i�*�@��#�]4@F�	j��!?��Ҳ�@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@�L�p��ٿm7�%,�@���s�3@q??��!?�=� ��@ٓ��s�ٿ/Z��,�@���c��3@�$"��!?A�d��@ٓ��s�ٿ/Z��,�@���c��3@�$"��!?A�d��@ٓ��s�ٿ/Z��,�@���c��3@�$"��!?A�d��@ٓ��s�ٿ/Z��,�@���c��3@�$"��!?A�d��@��Ǎ�ٿ��a6FE�@ըЂ��3@�a����!?�x���@��Ǎ�ٿ��a6FE�@ըЂ��3@�a����!?�x���@��Ǎ�ٿ��a6FE�@ըЂ��3@�a����!?�x���@����a�ٿ͕��=�@���F�3@cp'$��!?ܵ��K�@����a�ٿ͕��=�@���F�3@cp'$��!?ܵ��K�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@�����ٿ���G�C�@�����4@L����!?󪊄�@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@ʹ��Րٿ9f��C�@�����3@ꉄ�b�!?�z/µ@��z�ٿ��r	�P�@w0	� 4@�Ӽ�!?@�Y74�@��z�ٿ��r	�P�@w0	� 4@�Ӽ�!?@�Y74�@��z�ٿ��r	�P�@w0	� 4@�Ӽ�!?@�Y74�@��z�ٿ��r	�P�@w0	� 4@�Ӽ�!?@�Y74�@��z�ٿ��r	�P�@w0	� 4@�Ӽ�!?@�Y74�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@%��_f�ٿ�(6�E�@�c�3@�<��!?b�xjT-�@��)���ٿi�ޟM�@��Ip4@C#|V�!?�`C��.�@�ߣ*�ٿ]���D�@Y|B�
4@բ���!?�SN5���@�ߣ*�ٿ]���D�@Y|B�
4@բ���!?�SN5���@輝�}�ٿ^��W�@�腲4@͔$!?�~�є�@輝�}�ٿ^��W�@�腲4@͔$!?�~�є�@��r��ٿ�N��i�@8!���3@'JԾ?�!?ǹ��C�@��r��ٿ�N��i�@8!���3@'JԾ?�!?ǹ��C�@��r��ٿ�N��i�@8!���3@'JԾ?�!?ǹ��C�@��r��ٿ�N��i�@8!���3@'JԾ?�!?ǹ��C�@��r��ٿ�N��i�@8!���3@'JԾ?�!?ǹ��C�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@�4�M�ٿ�ⷞO^�@@�V2�3@O�x	��!?)�L�0�@5��]��ٿ�� �F�@Y��Y�3@HP��Ȑ!?�o`���@5��]��ٿ�� �F�@Y��Y�3@HP��Ȑ!?�o`���@��,�ٿ���4  �@N{����3@�#�ؐ!?�FE�>��@��,�ٿ���4  �@N{����3@�#�ؐ!?�FE�>��@Rgvw��ٿ����
�@N��c��3@��v�n�!?~�� ���@�8o�̔ٿc���^�@�ؿ��3@zj]��!?m1t��d�@�8o�̔ٿc���^�@�ؿ��3@zj]��!?m1t��d�@�8o�̔ٿc���^�@�ؿ��3@zj]��!?m1t��d�@ #J��ٿтw�?�@FV3�3@��]@+�!?��-�U��@ #J��ٿтw�?�@FV3�3@��]@+�!?��-�U��@ #J��ٿтw�?�@FV3�3@��]@+�!?��-�U��@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@�3��;�ٿ�&�"W�@�SWk*�3@T�r�4�!?����ǵ@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@Ʒ��ٿ�vT�@λk��3@����K�!?7����@y���ٿ�_��>�@@(����3@�N��+�!?�'���Ӵ@y���ٿ�_��>�@@(����3@�N��+�!?�'���Ӵ@y���ٿ�_��>�@@(����3@�N��+�!?�'���Ӵ@y���ٿ�_��>�@@(����3@�N��+�!?�'���Ӵ@y���ٿ�_��>�@@(����3@�N��+�!?�'���Ӵ@c�a���ٿ�L~K�8�@��ы:4@D�c<J�!?�>*�)��@c�a���ٿ�L~K�8�@��ы:4@D�c<J�!?�>*�)��@c�a���ٿ�L~K�8�@��ы:4@D�c<J�!?�>*�)��@c�a���ٿ�L~K�8�@��ы:4@D�c<J�!?�>*�)��@c�a���ٿ�L~K�8�@��ы:4@D�c<J�!?�>*�)��@g����ٿA7��fV�@\�i��3@�C=�.�!?���ʯ�@g����ٿA7��fV�@\�i��3@�C=�.�!?���ʯ�@g����ٿA7��fV�@\�i��3@�C=�.�!?���ʯ�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@n:5��ٿ�]�F!K�@��<��4@Җ�,��!?��^E1�@�t�AK�ٿ�x�$Jo�@�m����3@�y���!?y��_�@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@��63�ٿ�ME>�Z�@�Y9
��3@ⷞ��!?���۵@L�Y���ٿGCX��K�@���%�3@�1��!?���2�V�@L�Y���ٿGCX��K�@���%�3@�1��!?���2�V�@L�Y���ٿGCX��K�@���%�3@�1��!?���2�V�@L�Y���ٿGCX��K�@���%�3@�1��!?���2�V�@w�����ٿ�^X�@�@NM�4@��34�!?�&�{�@w�����ٿ�^X�@�@NM�4@��34�!?�&�{�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@�P��ٿ��\,�@	���3@ry}�!?y����;�@���w��ٿ
���;�@�HC7N4@�+��&�!?�װ?]�@���w��ٿ
���;�@�HC7N4@�+��&�!?�װ?]�@���w��ٿ
���;�@�HC7N4@�+��&�!?�װ?]�@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@���ۙٿ�_��ME�@��/7p4@�)�G�!?��^C��@.�kߒٿ8��;�q�@C�	�3@�@�L�!?ME=!�D�@.�kߒٿ8��;�q�@C�	�3@�@�L�!?ME=!�D�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@=1
B��ٿ?�R��g�@0���3@kژ�7�!?[��7�&�@z����ٿ�~�"��@�CF��3@���2��!?���\�Ӵ@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@ŧ�.��ٿ�# 卯�@�S�3f�3@%���!?h��e��@�-E��ٿůX����@MG�^�3@E:�J�!?��uCδ@��oQ��ٿ�����@*.��3@�2.A�!?��VU�۴@��oQ��ٿ�����@*.��3@�2.A�!?��VU�۴@��oQ��ٿ�����@*.��3@�2.A�!?��VU�۴@B�۠ܗٿk�%��M�@`ȅ���3@��1L�!?5\��.��@B�۠ܗٿk�%��M�@`ȅ���3@��1L�!?5\��.��@B�۠ܗٿk�%��M�@`ȅ���3@��1L�!?5\��.��@B�۠ܗٿk�%��M�@`ȅ���3@��1L�!?5\��.��@B�۠ܗٿk�%��M�@`ȅ���3@��1L�!?5\��.��@b�%���ٿD�x��B�@ �22�3@��C�6�!?��i�@b�%���ٿD�x��B�@ �22�3@��C�6�!?��i�@ c�%�ٿy$�2ZN�@���TA�3@0�x�!?�O��͵@V=�r �ٿ��vX�H�@(�]��3@��ʥ��!?-�.1���@V=�r �ٿ��vX�H�@(�]��3@��ʥ��!?-�.1���@V=�r �ٿ��vX�H�@(�]��3@��ʥ��!?-�.1���@V=�r �ٿ��vX�H�@(�]��3@��ʥ��!?-�.1���@����ٿA���6�@��E�N�3@�F���!?0d��@�@����ٿA���6�@��E�N�3@�F���!?0d��@�@����ٿA���6�@��E�N�3@�F���!?0d��@�@����ٿA���6�@��E�N�3@�F���!?0d��@�@����ٿA���6�@��E�N�3@�F���!?0d��@�@�\+���ٿ�[&��@���=�3@3�b|�!?������@�\+���ٿ�[&��@���=�3@3�b|�!?������@�\+���ٿ�[&��@���=�3@3�b|�!?������@a/#�h�ٿ]PA0��@@�;D�3@�����!?� �a��@a/#�h�ٿ]PA0��@@�;D�3@�����!?� �a��@��:�V�ٿ�]�����@�N�#4@(4��?�!?��텵@��:�V�ٿ�]�����@�N�#4@(4��?�!?��텵@��:�V�ٿ�]�����@�N�#4@(4��?�!?��텵@��:�V�ٿ�]�����@�N�#4@(4��?�!?��텵@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@']F�ٿKtY���@���J}�3@8a����!?ʝ�t�#�@���Ғٿ�󧚸`�@Ʈ��|�3@��E�!?�c�

��@���Ғٿ�󧚸`�@Ʈ��|�3@��E�!?�c�

��@2	ݔٿ��l�:�@yI��4@���u�!?�Jpz�)�@2	ݔٿ��l�:�@yI��4@���u�!?�Jpz�)�@2	ݔٿ��l�:�@yI��4@���u�!?�Jpz�)�@::cX�ٿY1@�N��@{��>�3@�����!?��w �@::cX�ٿY1@�N��@{��>�3@�����!?��w �@::cX�ٿY1@�N��@{��>�3@�����!?��w �@::cX�ٿY1@�N��@{��>�3@�����!?��w �@j⼑ٿ��,�]��@+�W�3@K��U�!?�;��@j⼑ٿ��,�]��@+�W�3@K��U�!?�;��@j⼑ٿ��,�]��@+�W�3@K��U�!?�;��@j⼑ٿ��,�]��@+�W�3@K��U�!?�;��@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@=���ٿ#�܍��@z�~/f�3@�[7�q�!?�l��I�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@��V��ٿ���Ư�@Z�
� �3@�`�A�!?F�rb�F�@#��눖ٿ�t;P�@��e�3@"�j�!?�[��@$�@#��눖ٿ�t;P�@��e�3@"�j�!?�[��@$�@#��눖ٿ�t;P�@��e�3@"�j�!?�[��@$�@#��눖ٿ�t;P�@��e�3@"�j�!?�[��@$�@#��눖ٿ�t;P�@��e�3@"�j�!?�[��@$�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@	0�2�ٿ�� )Ж�@'����3@=C���!?���a�k�@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@%�Y5]�ٿLw��[��@�ym%�3@3Pt&h�!?����Y��@r8���ٿ�4�L��@�?&��3@~
^���!?����,��@r8���ٿ�4�L��@�?&��3@~
^���!?����,��@r8���ٿ�4�L��@�?&��3@~
^���!?����,��@r8���ٿ�4�L��@�?&��3@~
^���!?����,��@r8���ٿ�4�L��@�?&��3@~
^���!?����,��@k�C���ٿHT��s�@LAS��3@Dg%�j�!?�;����@k�C���ٿHT��s�@LAS��3@Dg%�j�!?�;����@k�C���ٿHT��s�@LAS��3@Dg%�j�!?�;����@k�C���ٿHT��s�@LAS��3@Dg%�j�!?�;����@^*�x�ٿ�%R����@j�ws�3@�B�|S�!?7.Ɩ9ϴ@^*�x�ٿ�%R����@j�ws�3@�B�|S�!?7.Ɩ9ϴ@zb�F�ٿ�$h&��@oVf���3@U�z�!?,�@�V��@zb�F�ٿ�$h&��@oVf���3@U�z�!?,�@�V��@zb�F�ٿ�$h&��@oVf���3@U�z�!?,�@�V��@zb�F�ٿ�$h&��@oVf���3@U�z�!?,�@�V��@����ٿ�8} ���@A���h 4@�'�k
�!?��ͤ/��@	^(ٕٿ_��=��@;w��N�3@����U�!?ɕ0��@1�d[�ٿ�ɣ�>�@N���l4@'%A��!?C�-�S�@g��Ŕٿ=�H�*L�@���H24@Ѭ\�7�!??&HŴ@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@H��t�ٿŊ��a�@>�'��4@^F�6�!?�g�J��@�0UT�ٿ�m5���@���%�4@����`�!?P8�+gv�@�0UT�ٿ�m5���@���%�4@����`�!?P8�+gv�@�0UT�ٿ�m5���@���%�4@����`�!?P8�+gv�@�0UT�ٿ�m5���@���%�4@����`�!?P8�+gv�@�0UT�ٿ�m5���@���%�4@����`�!?P8�+gv�@����d�ٿx�Λ���@�D�[]4@oS�-t�!?������@�6�Y	�ٿ�N�0�-�@���%��3@��nV��!?]� �>E�@����ٿn1{'��@"O�n��3@��>��!?�7��@k�����ٿ�ru���@2�c��3@iC܄�!?M�$�]��@k�����ٿ�ru���@2�c��3@iC܄�!?M�$�]��@k�����ٿ�ru���@2�c��3@iC܄�!?M�$�]��@k�����ٿ�ru���@2�c��3@iC܄�!?M�$�]��@���께ٿ6��H9��@������3@��9$��!?v�I�]>�@���께ٿ6��H9��@������3@��9$��!?v�I�]>�@���께ٿ6��H9��@������3@��9$��!?v�I�]>�@���i�ٿ�ܡ��@�}�|��3@�m�٫�!?L!gi��@���i�ٿ�ܡ��@�}�|��3@�m�٫�!?L!gi��@���i�ٿ�ܡ��@�}�|��3@�m�٫�!?L!gi��@���i�ٿ�ܡ��@�}�|��3@�m�٫�!?L!gi��@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�Y?���ٿTń���@�}m4@�y�
%�!?%�X=�@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@�����ٿk `�,�@Y��i�4@�����!?=O����@���G�ٿ,-���@1-1�3@2�	��!?��q&g��@���G�ٿ,-���@1-1�3@2�	��!?��q&g��@���G�ٿ,-���@1-1�3@2�	��!?��q&g��@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@�'�8Ôٿ� ����@�	�Kh�3@��' ��!?��3����@U<|Ԗٿ_�����@���-�3@Հ�ﻐ!?�DI0�3�@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@��.�ٿ���%��@+^���3@�;m~�!?1��Bϵ@�y�Bz�ٿ8�!�@0���&�3@7����!?R/�Vٵ@�y�Bz�ٿ8�!�@0���&�3@7����!?R/�Vٵ@�y�Bz�ٿ8�!�@0���&�3@7����!?R/�Vٵ@�y�Bz�ٿ8�!�@0���&�3@7����!?R/�Vٵ@�y�Bz�ٿ8�!�@0���&�3@7����!?R/�Vٵ@Q�����ٿ-��({M�@��1��3@2�!?������@Q�����ٿ-��({M�@��1��3@2�!?������@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@r�4�˒ٿs��<��@���3@X���!?���p,�@!��o�ٿ]ֳo��@? 	���3@���@��!?�] ,>�@!��o�ٿ]ֳo��@? 	���3@���@��!?�] ,>�@!��o�ٿ]ֳo��@? 	���3@���@��!?�] ,>�@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@N>�ٿ�H`2�b�@�쯥��3@�p`�!?����@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@6vl�$�ٿ�*eu��@�����3@g�`6�!?�5��4�@�qt1n�ٿb��#�@�B*=0�3@7җVL�!?4��nX��@�qt1n�ٿb��#�@�B*=0�3@7җVL�!?4��nX��@�qt1n�ٿb��#�@�B*=0�3@7җVL�!?4��nX��@�qt1n�ٿb��#�@�B*=0�3@7җVL�!?4��nX��@���,�ٿ��r���@��O��3@�}ǫ�!?[Kl��ٴ@���,�ٿ��r���@��O��3@�}ǫ�!?[Kl��ٴ@���,�ٿ��r���@��O��3@�}ǫ�!?[Kl��ٴ@�����ٿ�"�|V9�@�|�1m�3@�I��8�!?&^��Z��@���J�ٿ��CҘ�@#Aˋ�3@5�0�!?|��L�ӵ@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@ڀh��ٿ�)[t�,�@<��n)�3@�2�%�!?IN�s��@o���z�ٿ�v6��@R�L<-�3@8Bs͏!?_v��@�@o���z�ٿ�v6��@R�L<-�3@8Bs͏!?_v��@�@�����ٿ� +mZE�@�`�]��3@z�kK�!?�����@�����ٿ� +mZE�@�`�]��3@z�kK�!?�����@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@&���_�ٿ[����@�O��g�3@IoĴ�!?������@5�􊪑ٿR�Ϣf�@�\L �3@m���!?8���@5�􊪑ٿR�Ϣf�@�\L �3@m���!?8���@5�􊪑ٿR�Ϣf�@�\L �3@m���!?8���@5�􊪑ٿR�Ϣf�@�\L �3@m���!?8���@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�����ٿ(��^���@j�2
"�3@C�+�!?��2Q��@�B���ٿ��5rU��@���x��3@6��E�!?<�aa�~�@�B���ٿ��5rU��@���x��3@6��E�!?<�aa�~�@�B���ٿ��5rU��@���x��3@6��E�!?<�aa�~�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@Ղ�2�ٿ98-hn��@j5��3@�_��J�!?`v+e�%�@ℵ���ٿ��WےD�@r���3@�M����!?��BY;8�@�1|.�ٿhb!�f��@:m�}� 4@V�	W�!?�$?qb̴@�1|.�ٿhb!�f��@:m�}� 4@V�	W�!?�$?qb̴@�1|.�ٿhb!�f��@:m�}� 4@V�	W�!?�$?qb̴@�И�^�ٿ���-��@�Զ_��3@Y -�l�!?O8_�ct�@�И�^�ٿ���-��@�Զ_��3@Y -�l�!?O8_�ct�@�И�^�ٿ���-��@�Զ_��3@Y -�l�!?O8_�ct�@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@��,a�ٿ �z�N�@JjB�f�3@���?�!?��Er��@�ά���ٿ�Ɍr(h�@
br9�3@,]|�~�!?������@�ά���ٿ�Ɍr(h�@
br9�3@,]|�~�!?������@+s7��ٿ@�&�4�@�;���3@����z�!?�@����@l��BŘٿFgm�W��@+�E��4@�|��d�!?��F�xA�@l��BŘٿFgm�W��@+�E��4@�|��d�!?��F�xA�@l��BŘٿFgm�W��@+�E��4@�|��d�!?��F�xA�@�j��z�ٿ#��i�@���4@�Ïw�!?���f�ٵ@m�q��ٿ+��w.��@DB7��3@��B�X�!?��a�u�@t~H��ٿε��H�@fV��3@�2�͆�!?�}��w�@t~H��ٿε��H�@fV��3@�2�͆�!?�}��w�@t~H��ٿε��H�@fV��3@�2�͆�!?�}��w�@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@-��ѷ�ٿ�Тu�"�@7��D�3@ �h<2�!?Q��ө��@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@��utM�ٿ1��JC��@WB|o�3@�l:9�!?�zdkVߴ@?�fĖٿ��" �"�@�W�{�3@��b�T�!?K�X����@|iD��ٿk<ni��@��q���3@^�cz�!?��J�۴@|iD��ٿk<ni��@��q���3@^�cz�!?��J�۴@��z�+�ٿ����@���O�3@���k�!?L-����@IOMj��ٿ�����@ ����3@X%��~�!?�@P�Fܴ@IOMj��ٿ�����@ ����3@X%��~�!?�@P�Fܴ@IOMj��ٿ�����@ ����3@X%��~�!?�@P�Fܴ@Yc��e�ٿ�{�O6�@dC���3@
��FB�!?�OŴ@Yc��e�ٿ�{�O6�@dC���3@
��FB�!?�OŴ@k�ّ`�ٿf��eS�@�0+d��3@��:�!?���<1;�@f���,�ٿn\��AJ�@P
����3@Y���!?���K�@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@ǫ��ٿ �U3T�@�)�1��3@�d��S�!?Љ8Jdڴ@�/i�#�ٿ��90���@�;�3!�3@���!?PDZ���@�/i�#�ٿ��90���@�;�3!�3@���!?PDZ���@�/i�#�ٿ��90���@�;�3!�3@���!?PDZ���@m�[�ٿEZ�E=��@~So}34@�V!�\�!?e�t���@m�[�ٿEZ�E=��@~So}34@�V!�\�!?e�t���@b��I�ٿ��G�h	�@���m��3@6����!?g(h�H(�@·���ٿ�l+�4��@r>���3@W~T���!?�`�C6�@�hԜ�ٿ��^B��@�n��3@&d�N�!?�F;5�,�@�hԜ�ٿ��^B��@�n��3@&d�N�!?�F;5�,�@�hԜ�ٿ��^B��@�n��3@&d�N�!?�F;5�,�@�hԜ�ٿ��^B��@�n��3@&d�N�!?�F;5�,�@�hԜ�ٿ��^B��@�n��3@&d�N�!?�F;5�,�@���x�ٿ(�g���@o85v14@�M��5�!?�x���%�@^�x%�ٿu�q���@+Vs���3@qX�n(�!?���ҹ�@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@���a�ٿ� ߸D�@V:[��3@�#�_&�!?��|E۴@Y�>TƘٿ������@c��B}�3@�a�Q�!?�)Q)�@Y�>TƘٿ������@c��B}�3@�a�Q�!?�)Q)�@Y�>TƘٿ������@c��B}�3@�a�Q�!?�)Q)�@��gcL�ٿ���h��@�l�"�3@p�.��!?��.>�@��gcL�ٿ���h��@�l�"�3@p�.��!?��.>�@��gcL�ٿ���h��@�l�"�3@p�.��!?��.>�@]�};ԙٿ����@S��� 4@ �k�!?�^��]}�@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@젮��ٿa��~i�@gE�D��3@��?�P�!?���)��@.�ŢR�ٿ�#�$��@àrg��3@�<��F�!?��5Q��@.�ŢR�ٿ�#�$��@àrg��3@�<��F�!?��5Q��@.�ŢR�ٿ�#�$��@àrg��3@�<��F�!?��5Q��@.�ŢR�ٿ�#�$��@àrg��3@�<��F�!?��5Q��@.�ŢR�ٿ�#�$��@àrg��3@�<��F�!?��5Q��@���u��ٿ"���g^�@�A_��3@��=��!?Pe��'�@��Z��ٿ�LX��@�Y�6�3@F�Ci�!?���mc�@��Z��ٿ�LX��@�Y�6�3@F�Ci�!?���mc�@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@,�=�ӡٿ�% �o��@U�Sk�3@xf��Q�!?�p�}�ɴ@���ٿ�@6����@�V>��3@T0#e�!?����@Է��+�ٿ��i/S�@|�+��3@k��dS�!?!G�vcW�@~��ŝٿ�H�`�@�l�;��3@�t�p�!?��CN�6�@���\�ٿp*m����@�4w��3@&䩞s�!?Q�E�n��@���\�ٿp*m����@�4w��3@&䩞s�!?Q�E�n��@D���ژٿޫ���+�@�.��3@�@ُ!?3�#��w�@D���ژٿޫ���+�@�.��3@�@ُ!?3�#��w�@D���ژٿޫ���+�@�.��3@�@ُ!?3�#��w�@D���ژٿޫ���+�@�.��3@�@ُ!?3�#��w�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@�q>�ٿ/|�6��@���9��3@adr�ڏ!?Z��~�@��ٿ�mf���@Ŏ����3@K��&�!?R-)P삵@��Ie�ٿ�V%�<�@�	m��3@ :���!?�"*!��@�O�s�ٿ������@U�%��3@��C#W�!?rԬ�C�@���s�ٿ|t��W�@�m�� �3@�;����!?��oRl�@���R�ٿ}�2��@Mz4��3@i؟ϸ�!?;�elO�@~��lj�ٿ��Ҿ��@��5���3@���MK�!?����e	�@~��lj�ٿ��Ҿ��@��5���3@���MK�!?����e	�@~��lj�ٿ��Ҿ��@��5���3@���MK�!?����e	�@~��lj�ٿ��Ҿ��@��5���3@���MK�!?����e	�@�B��ٿ�%]���@!8y�z�3@f���~�!?��Lb�&�@�B��ٿ�%]���@!8y�z�3@f���~�!?��Lb�&�@u/Ǒ�ٿ͙��`�@bPJN�3@��-]�!?�p��R�@Qg�Иٿ�Ͻ<�,�@�d|~y�3@B�O��!?W���n�@Qg�Иٿ�Ͻ<�,�@�d|~y�3@B�O��!?W���n�@Qg�Иٿ�Ͻ<�,�@�d|~y�3@B�O��!?W���n�@Qg�Иٿ�Ͻ<�,�@�d|~y�3@B�O��!?W���n�@Qg�Иٿ�Ͻ<�,�@�d|~y�3@B�O��!?W���n�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@��N��ٿ�V#!K�@Ʊ�\�3@-THH�!?�^��,�@�z�m��ٿG�]���@Y�<I��3@���VJ�!??�Z��@�z�m��ٿG�]���@Y�<I��3@���VJ�!??�Z��@�z�m��ٿG�]���@Y�<I��3@���VJ�!??�Z��@�z�m��ٿG�]���@Y�<I��3@���VJ�!??�Z��@�z�m��ٿG�]���@Y�<I��3@���VJ�!??�Z��@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@k.l�ٿt�!VA��@�q�u�3@��r�!?�:����@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@�2�p�ٿ�U(}�@�]
�=�3@P��Y��!?��r�+�@#��s�ٿ?<����@E4���3@�S�x�!?t4�Po��@1%���ٿZ,b����@g<�7��3@��	[��!?�rB���@1%���ٿZ,b����@g<�7��3@��	[��!?�rB���@1%���ٿZ,b����@g<�7��3@��	[��!?�rB���@1%���ٿZ,b����@g<�7��3@��	[��!?�rB���@���O�ٿ�k����@����>�3@U�Zi�!?..���g�@���O�ٿ�k����@����>�3@U�Zi�!?..���g�@���O�ٿ�k����@����>�3@U�Zi�!?..���g�@����K�ٿ 2��4�@bx���3@pH��X�!?�2���w�@����K�ٿ 2��4�@bx���3@pH��X�!?�2���w�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@a� ��ٿ������@�A>}g�3@�}�Aa�!?�����?�@��%_�ٿJ��"cA�@�O@p�3@���Lf�!?ُA�ű�@��%_�ٿJ��"cA�@�O@p�3@���Lf�!?ُA�ű�@��%_�ٿJ��"cA�@�O@p�3@���Lf�!?ُA�ű�@��%_�ٿJ��"cA�@�O@p�3@���Lf�!?ُA�ű�@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@���W�ٿ�o�Z��@��t5�4@�bS�#�!?v�)E�ٴ@�1�"�ٿ��/���@��C-�3@v�W�X�!?j����@�1�"�ٿ��/���@��C-�3@v�W�X�!?j����@Y;�ٿה\Y�8�@����3@�r�!?=j���s�@Y;�ٿה\Y�8�@����3@�r�!?=j���s�@�~>�B�ٿ�[�1�W�@6��;	�3@��N��!?������@�~>�B�ٿ�[�1�W�@6��;	�3@��N��!?������@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@��8�#�ٿ���t�3�@^�`$�3@��0�!?oXq��@�FF0�ٿ�I��y��@��h�3@�pW��!?<}y7B��@�FF0�ٿ�I��y��@��h�3@�pW��!?<}y7B��@�FF0�ٿ�I��y��@��h�3@�pW��!?<}y7B��@�ƌPC�ٿ^��w�S�@%i�R��3@ӶrY�!?/6a�Zy�@�ƌPC�ٿ^��w�S�@%i�R��3@ӶrY�!?/6a�Zy�@�جt֜ٿ�cQ �@�&����3@R�:r��!?,K��H�@��}��ٿ���1%��@� ��3@�oV��!?�m�
�@>Hө�ٿ�{���@���@`�3@�J����!?�<��˴@>Hө�ٿ�{���@���@`�3@�J����!?�<��˴@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@H��B�ٿ&m[)��@AME��3@�j���!?&
��@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@Cw��_�ٿ�缝
��@`����4@��C@��!?�:�h�Ŵ@�^@�ٿ69I#2>�@G,�q�3@������!?C�����@�^@�ٿ69I#2>�@G,�q�3@������!?C�����@�^@�ٿ69I#2>�@G,�q�3@������!?C�����@��;4�ٿ��'��@O�&t��3@-�QM؏!?s�vʨ�@��;4�ٿ��'��@O�&t��3@-�QM؏!?s�vʨ�@��;4�ٿ��'��@O�&t��3@-�QM؏!?s�vʨ�@��;4�ٿ��'��@O�&t��3@-�QM؏!?s�vʨ�@���'�ٿn��C��@F�Y�Y�3@$��U�!?8�-'�@���'�ٿn��C��@F�Y�Y�3@$��U�!?8�-'�@���'�ٿn��C��@F�Y�Y�3@$��U�!?8�-'�@�#pR��ٿ�琪���@%�Pe��3@�cø�!?U"6��ʹ@zt�c�ٿ�i�Po�@�q���3@&�[^�!?@���@zt�c�ٿ�i�Po�@�q���3@&�[^�!?@���@zt�c�ٿ�i�Po�@�q���3@&�[^�!?@���@|�Ǎ�ٿ�p����@�>h�3@IY���!?�=Q ��@|�Ǎ�ٿ�p����@�>h�3@IY���!?�=Q ��@|�Ǎ�ٿ�p����@�>h�3@IY���!?�=Q ��@|�Ǎ�ٿ�p����@�>h�3@IY���!?�=Q ��@|�Ǎ�ٿ�p����@�>h�3@IY���!?�=Q ��@X/�u�ٿ��د�y�@�S�U�3@wݨ[Y�!?y�H)ģ�@X/�u�ٿ��د�y�@�S�U�3@wݨ[Y�!?y�H)ģ�@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@��W��ٿf5�ª��@e�Q��3@_�u�!?B~.ʴ@H�
T��ٿDZc��*�@��5��3@��'b�!?.x�޴@�L{�S�ٿ �f7>~�@uù[.�3@�̚k�!?o�����@�L{�S�ٿ �f7>~�@uù[.�3@�̚k�!?o�����@�H�ٿ��~cK��@Ns���3@$���!?�u�״�@�H�ٿ��~cK��@Ns���3@$���!?�u�״�@�H�ٿ��~cK��@Ns���3@$���!?�u�״�@�H�ٿ��~cK��@Ns���3@$���!?�u�״�@�H�ٿ��~cK��@Ns���3@$���!?�u�״�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@���w��ٿ��H���@�(���3@�s� l�!?0��n�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@O��}�ٿ;Z8/�@�qZIn�3@�hm8�!?!#h��>�@��R�ٿ(�����@�b��>�3@�m�b�!?L"�Tش@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@���{�ٿ[�[s!��@ѓ>%0�3@)�|�}�!?6��s���@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@�dj�ٿ4VDS��@���L�3@�[7�K�!?{1x�  �@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@a�,di�ٿ��R����@v���3@�g��u�!?(�h�1�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@7fy 
�ٿ3�{���@:,����3@Z8����!?�K+�F�@Q�	n�ٿO��DO)�@��r�j�3@��f�#�!?��6ݢZ�@/��#M�ٿ�*��a9�@Imۡ��3@a =v@�!?��xL�@/��#M�ٿ�*��a9�@Imۡ��3@a =v@�!?��xL�@/��#M�ٿ�*��a9�@Imۡ��3@a =v@�!?��xL�@/��#M�ٿ�*��a9�@Imۡ��3@a =v@�!?��xL�@/��#M�ٿ�*��a9�@Imۡ��3@a =v@�!?��xL�@~7{��ٿ���;��@{a=��3@�J�u�!?X�_g�@�)AS�ٿ��L���@#�� ��3@]���!?�ϫ"'�@�)AS�ٿ��L���@#�� ��3@]���!?�ϫ"'�@�\]Y�ٿ����@�����3@c�vg�!?�Hմ@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�7K�ٿFV2@�@�&�3@S���r�!?�	�2��@�!
*�ٿ�7?��@�9d��3@�k�R�!?,�7���@PF���ٿ�PLI)�@Ï�P��3@��c��!?C�d��@PF���ٿ�PLI)�@Ï�P��3@��c��!?C�d��@PF���ٿ�PLI)�@Ï�P��3@��c��!?C�d��@R�),�ٿ�dnv��@b�Oy�4@�e�j�!?����´@R�),�ٿ�dnv��@b�Oy�4@�e�j�!?����´@���	E�ٿU>��M�@0�0?4@��B:�!?�a\Nδ@���	E�ٿU>��M�@0�0?4@��B:�!?�a\Nδ@���	E�ٿU>��M�@0�0?4@��B:�!?�a\Nδ@���	E�ٿU>��M�@0�0?4@��B:�!?�a\Nδ@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@�I1@�ٿ*�bͦU�@�gmҮ�3@L6�U�!?
r���@Ɖ�=�ٿ*��ǋ��@�]<"�3@�~�T�!?��Y��@Ɖ�=�ٿ*��ǋ��@�]<"�3@�~�T�!?��Y��@�v;�Y�ٿ?!��$��@$�*,�3@j����!?)�U�}�@�Ѿ�ʔٿU��?�@Z��� 4@U�A��!?۞����@�V�B��ٿ���xN�@<c.f4@�$d�!?����<*�@�V�B��ٿ���xN�@<c.f4@�$d�!?����<*�@��lT�ٿr~��D��@��� 4@��w�,�!?s���l̴@����k�ٿy��؇�@Ϳ����3@a��	N�!?"Ah�B�@W�p���ٿu����@e�G�,�3@9E�3�!?ze�Xkִ@�9�j��ٿE���=�@H�Ǌn 4@ИiL�!?�`��Ǵ@�9�j��ٿE���=�@H�Ǌn 4@ИiL�!?�`��Ǵ@�9�j��ٿE���=�@H�Ǌn 4@ИiL�!?�`��Ǵ@�9�j��ٿE���=�@H�Ǌn 4@ИiL�!?�`��Ǵ@�9�j��ٿE���=�@H�Ǌn 4@ИiL�!?�`��Ǵ@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@ d����ٿk�{؍.�@�����4@���T"�!?�����@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@��	���ٿ�����@h[S�3@Za���!?]�A]b�@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@�T���ٿ��?
���@b:oa�3@�K>�U�!?�H_V��@��$zE�ٿ/���@��p<��3@��v�0�!?c{*v�W�@��$zE�ٿ/���@��p<��3@��v�0�!?c{*v�W�@��$zE�ٿ/���@��p<��3@��v�0�!?c{*v�W�@��$zE�ٿ/���@��p<��3@��v�0�!?c{*v�W�@3Ɯ웑ٿ,<Ƿ��@J����3@�N���!?`�Rb�K�@3Ɯ웑ٿ,<Ƿ��@J����3@�N���!?`�Rb�K�@3Ɯ웑ٿ,<Ƿ��@J����3@�N���!?`�Rb�K�@�� �ٿL����E�@n�UH�4@���!?�(I�?�@�'\���ٿ��څ3&�@U�'J�3@o����!?��K���@�'\���ٿ��څ3&�@U�'J�3@o����!?��K���@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@�T���ٿ#NFRP?�@�/Y ��3@MGTC�!?w~�BT�@.K��\�ٿ�t9�ݵ�@�ygN�3@s��!? ��"��@�?a�x�ٿ��D#5�@:1�"��3@~i��<�!?0�d�Q]�@�?a�x�ٿ��D#5�@:1�"��3@~i��<�!?0�d�Q]�@�?a�x�ٿ��D#5�@:1�"��3@~i��<�!?0�d�Q]�@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@ŰP�ٿ�^�I�:�@j�YV�3@&�*U�!?z��$��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�܅w��ٿe"z��I�@%�����3@�@��/�!?���P��@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@�����ٿ����@PK��^�3@Q�?i�!?AQ�WZA�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@c5Dr��ٿХ�]�@d��3@)aQM�!?�X��{&�@QO�PٿeWg��@�mlF��3@8Qr�!?�l�6��@QO�PٿeWg��@�mlF��3@8Qr�!?�l�6��@QO�PٿeWg��@�mlF��3@8Qr�!?�l�6��@QO�PٿeWg��@�mlF��3@8Qr�!?�l�6��@�^�Ie�ٿ�`���@0����3@>��E�!?K��x�@9Ʉ:�ٿ`���V�@̅?z�3@�`�I?�!?z���K��@9Ʉ:�ٿ`���V�@̅?z�3@�`�I?�!?z���K��@�g{S��ٿh2�����@������3@<�胐!?_KLD��@�g{S��ٿh2�����@������3@<�胐!?_KLD��@�g{S��ٿh2�����@������3@<�胐!?_KLD��@�Y�|�ٿ�y�|i�@iŮ�y�3@�Nh)�!?���H��@�Y�|�ٿ�y�|i�@iŮ�y�3@�Nh)�!?���H��@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@��k�W�ٿ��y'U��@Sly�Z�3@d�����!?������@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@Ċ�a�ٿn|;F�@�0���3@��3�R�!?*��?���@��d�ٿI��Vm�@��A;�3@�A�~�!?�{v�@��d�ٿI��Vm�@��A;�3@�A�~�!?�{v�@��d�ٿI��Vm�@��A;�3@�A�~�!?�{v�@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@r"h�/�ٿ	t�����@�)"1��3@!B�4(�!?�I'�~ݴ@h� �ٿ�Ys���@�v'"�3@&L��!?�^2�{�@c�+ѭ�ٿ�K	��@H���)�3@l�	�!?Q`d��@c�+ѭ�ٿ�K	��@H���)�3@l�	�!?Q`d��@m5����ٿ����ų�@��F� �3@�i����!?Ҥ�Շ�@m5����ٿ����ų�@��F� �3@�i����!?Ҥ�Շ�@m5����ٿ����ų�@��F� �3@�i����!?Ҥ�Շ�@m5����ٿ����ų�@��F� �3@�i����!?Ҥ�Շ�@m5����ٿ����ų�@��F� �3@�i����!?Ҥ�Շ�@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@�k��5�ٿ���=J�@Vh��3@�aߎR�!?A,�����@��Aٿ;�/R!��@b�8��3@輳oo�!?�����@��Aٿ;�/R!��@b�8��3@輳oo�!?�����@��Aٿ;�/R!��@b�8��3@輳oo�!?�����@��Aٿ;�/R!��@b�8��3@輳oo�!?�����@�ض�A�ٿl���b��@�`���3@�A�/��!?�=��@�ض�A�ٿl���b��@�`���3@�A�/��!?�=��@�ض�A�ٿl���b��@�`���3@�A�/��!?�=��@�ض�A�ٿl���b��@�`���3@�A�/��!?�=��@�ض�A�ٿl���b��@�`���3@�A�/��!?�=��@�,��֎ٿ�Λ����@q�ŗo�3@��|�V�!?Q
����@�,��֎ٿ�Λ����@q�ŗo�3@��|�V�!?Q
����@�,��֎ٿ�Λ����@q�ŗo�3@��|�V�!?Q
����@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@���֑ٿ](�M�@[ �34@

�k�!?U���@��c�s�ٿ�\����@Omq�g�3@i����!?���:�@�f���ٿ����E�@!\�M��3@�����!?i/�`�@�f���ٿ����E�@!\�M��3@�����!?i/�`�@�f���ٿ����E�@!\�M��3@�����!?i/�`�@����T�ٿ�3l��@DUC��3@�((X%�!?�������@����T�ٿ�3l��@DUC��3@�((X%�!?�������@�{��ٿߊ$�Z4�@�-
�Q�3@��ĕ�!?����e6�@�{��ٿߊ$�Z4�@�-
�Q�3@��ĕ�!?����e6�@�{��ٿߊ$�Z4�@�-
�Q�3@��ĕ�!?����e6�@�{��ٿߊ$�Z4�@�-
�Q�3@��ĕ�!?����e6�@�{��ٿߊ$�Z4�@�-
�Q�3@��ĕ�!?����e6�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@]�.U��ٿ�*�l���@i�����3@�*S)�!?j��c�@������ٿ�
{-I�@�=s�3@O����!?��s���@������ٿ�
{-I�@�=s�3@O����!?��s���@�!9
P�ٿUWl�^��@ ����3@�)�H�!?�����i�@�!9
P�ٿUWl�^��@ ����3@�)�H�!?�����i�@�!/8�ٿ_�����@tGR�8�3@PX~y�!?@%"��@�!/8�ٿ_�����@tGR�8�3@PX~y�!?@%"��@�!/8�ٿ_�����@tGR�8�3@PX~y�!?@%"��@�!/8�ٿ_�����@tGR�8�3@PX~y�!?@%"��@�!/8�ٿ_�����@tGR�8�3@PX~y�!?@%"��@��E���ٿ��m��@�@�Y��w�3@ȥ��s�!?��ŧ���@��E���ٿ��m��@�@�Y��w�3@ȥ��s�!?��ŧ���@��E���ٿ��m��@�@�Y��w�3@ȥ��s�!?��ŧ���@��E���ٿ��m��@�@�Y��w�3@ȥ��s�!?��ŧ���@���BH�ٿNX�8�@�yA���3@
���o�!? �){��@���BH�ٿNX�8�@�yA���3@
���o�!? �){��@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@\�X��ٿ���v�@��1e�4@��+�!?��	16ߵ@S,�W��ٿ�o�j���@D�b"�4@�\1��!?X�(����@Fb��3�ٿv��Ŵ�@r��9��3@7cu�!?�y�Wف�@Fb��3�ٿv��Ŵ�@r��9��3@7cu�!?�y�Wف�@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@�Q5N�ٿ���y7�@�����3@�,"�O�!?Nڬ ��@��ިL�ٿ۶���@]���3@�lB��!?'�ӄ ��@��ިL�ٿ۶���@]���3@�lB��!?'�ӄ ��@��ިL�ٿ۶���@]���3@�lB��!?'�ӄ ��@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@{AW��ٿ�F=���@��(V>�3@u.���!?C �c�j�@�̡zc�ٿr�yc��@�()Ye�3@�+�Z�!?M'C�@�̡zc�ٿr�yc��@�()Ye�3@�+�Z�!?M'C�@���ٿ�]c���@�K�:�3@"i ���!?�ߐĩ�@���Z�ٿ�?]\=��@M�+���3@"Zא!?��8�h@�@���Z�ٿ�?]\=��@M�+���3@"Zא!?��8�h@�@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@�G�z�ٿ.9�\�k�@����3@��jt�!?�>����@x�;؂�ٿ.��f�@ך|��	4@[\�j)�!?j�$�3�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@i%�f�ٿE��5:�@��14@DQsQV�!?��,�WA�@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@��x�%�ٿ�y�s�Q�@�ܴ�o�3@LΌ�c�!?��鴴@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@���ٿ�_l����@�D����3@�NǙN�!?>����ٴ@ɘ�>A�ٿ��i&C��@y0.%�3@A�>n�!?�2vtд@�g��
�ٿ�/���@#3��u�3@�9��P�!?�{wJ&�@�g��
�ٿ�/���@#3��u�3@�9��P�!?�{wJ&�@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@ 3����ٿ�#�����@+b�x�3@r|�z��!?��}+���@s��ؗٿ����~��@����3@�5�_��!?N"�����@s��ؗٿ����~��@����3@�5�_��!?N"�����@s��ؗٿ����~��@����3@�5�_��!?N"�����@s��ؗٿ����~��@����3@�5�_��!?N"�����@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@uky�L�ٿy�Ѯ��@�^�#I�3@���F�!?]@��-�@n�	��ٿ �*i���@�P��>4@�����!?��ѡ��@�#Gb��ٿ���t��@�%cx_�3@���!?��R�H��@�#Gb��ٿ���t��@�%cx_�3@���!?��R�H��@�#Gb��ٿ���t��@�%cx_�3@���!?��R�H��@�#Gb��ٿ���t��@�%cx_�3@���!?��R�H��@�#Gb��ٿ���t��@�%cx_�3@���!?��R�H��@�h�Qc�ٿ"�z[�@I�Ty�4@�1�]�!?��E8��@��m4Ɲٿ��T�t�@����4@��O�!�!?�=���@��m4Ɲٿ��T�t�@����4@��O�!�!?�=���@��m4Ɲٿ��T�t�@����4@��O�!�!?�=���@��m4Ɲٿ��T�t�@����4@��O�!�!?�=���@ѹM:��ٿ��l����@��9��3@5�'誐!?�>�����@ѹM:��ٿ��l����@��9��3@5�'誐!?�>�����@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@6����ٿ��@��@x�%���3@�X�<��!?S�)��@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@�m�7ڝٿ� ]�.��@���zB�3@�9,ې!?��|E�@L��-�ٿ��&	���@ȵ6��3@��(�ِ!?z�:L��@L��-�ٿ��&	���@ȵ6��3@��(�ِ!?z�:L��@L��-�ٿ��&	���@ȵ6��3@��(�ِ!?z�:L��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@�m���ٿ{Z�s�A�@�b���3@[z��t�!?�TJ��@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@��s{�ٿA;�:_��@(k�%�3@ZV�|�!?N�J&�˴@�v.��ٿ��)oZo�@��%�#�3@s��{�!?Ͱp�!�@�v.��ٿ��)oZo�@��%�#�3@s��{�!?Ͱp�!�@�v.��ٿ��)oZo�@��%�#�3@s��{�!?Ͱp�!�@�v.��ٿ��)oZo�@��%�#�3@s��{�!?Ͱp�!�@8�$��ٿd� r���@}�`1 4@G�+L�!?������@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@��}f�ٿD�8���@2kw�4@�O���!?O 6�n�@TD�h�ٿ��ă��@�Wч��3@3 �'�!?B������@TD�h�ٿ��ă��@�Wч��3@3 �'�!?B������@z?�dj�ٿ+���B�@�&�~�4@�����!?|��] Ҵ@z?�dj�ٿ+���B�@�&�~�4@�����!?|��] Ҵ@z?�dj�ٿ+���B�@�&�~�4@�����!?|��] Ҵ@�x�#�ٿuțN��@���3�3@���l-�!?�c��C�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@.�� �ٿn���$�@T�UL�3@�b2��!?S��~�@��!mښٿ+��z�@�̳��3@�)~��!?њ;S=ʴ@��!mښٿ+��z�@�̳��3@�)~��!?њ;S=ʴ@��!mښٿ+��z�@�̳��3@�)~��!?њ;S=ʴ@��!mښٿ+��z�@�̳��3@�)~��!?њ;S=ʴ@��!mښٿ+��z�@�̳��3@�)~��!?њ;S=ʴ@��~ɺ�ٿ
s8�)�@L����3@�B���!?d����۴@�=5Q�ٿG+���@@�qӚ�3@M�����!?^���״@�=5Q�ٿG+���@@�qӚ�3@M�����!?^���״@M�T)��ٿ�d����@[�6Γ�3@n
�Qa�!?3Q����@M�T)��ٿ�d����@[�6Γ�3@n
�Qa�!?3Q����@M�T)��ٿ�d����@[�6Γ�3@n
�Qa�!?3Q����@B4I}��ٿR9j��@]�e	��3@����!?x�!@mɴ@B4I}��ٿR9j��@]�e	��3@����!?x�!@mɴ@��Cі�ٿpv���@�>i��3@a�EY7�!?5�yƖ�@��Cі�ٿpv���@�>i��3@a�EY7�!?5�yƖ�@��Cі�ٿpv���@�>i��3@a�EY7�!?5�yƖ�@��Cі�ٿpv���@�>i��3@a�EY7�!?5�yƖ�@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@��{Ɨٿ����w�@�T��3@���Y�!?������@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@e��j^�ٿ>q����@mds���3@�#�]h�!?E�3T'��@jiib��ٿ�_�����@�oH)�3@�p/���!?>�i7h�@��3�ٿ��f����@�p>G�3@p�|�;�!?�kM�Y�@��3�ٿ��f����@�p>G�3@p�|�;�!?�kM�Y�@��3�ٿ��f����@�p>G�3@p�|�;�!?�kM�Y�@��3�ٿ��f����@�p>G�3@p�|�;�!?�kM�Y�@"2��
�ٿ���_��@j�u��3@ɔ�؏!?J�Ź+'�@"2��
�ٿ���_��@j�u��3@ɔ�؏!?J�Ź+'�@"2��
�ٿ���_��@j�u��3@ɔ�؏!?J�Ź+'�@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@������ٿ���T��@����3@FY�)Q�!?d���9Ĵ@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@O�h(k�ٿP�$E�w�@��$x�3@��4�H�!?n.=�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@�wE��ٿ/i�[7)�@]�{��3@��!?E��QƦ�@8�2$ڏٿ�a��>�@u4F�3@t4}P/�!?1���ݴ@8�2$ڏٿ�a��>�@u4F�3@t4}P/�!?1���ݴ@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@�؏2�ٿ(��oY0�@{��4@Bhu_��!?���u:R�@V�<�5�ٿ G<f\,�@镎��3@LN��!?Y�b3���@68�;O�ٿ�D�po��@O��|=�3@jĚ��!?����@68�;O�ٿ�D�po��@O��|=�3@jĚ��!?����@68�;O�ٿ�D�po��@O��|=�3@jĚ��!?����@���.�ٿ�@��a��@�b*R4�3@$���!?�K�d�@�~�	�ٿ,���@�%���3@a��D��!?aws���@�~�	�ٿ,���@�%���3@a��D��!?aws���@��U��ٿ�q��Xz�@��>��3@����!?0Z��A�@��U��ٿ�q��Xz�@��>��3@����!?0Z��A�@��U��ٿ�q��Xz�@��>��3@����!?0Z��A�@I)�p!�ٿ����@ݚ��u�3@W�ic8�!?�\��w�@I)�p!�ٿ����@ݚ��u�3@W�ic8�!?�\��w�@I)�p!�ٿ����@ݚ��u�3@W�ic8�!?�\��w�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@�����ٿ�w䋩g�@=�ǰp�3@�p��j�!?P�9�e6�@Q��זٿj�� ��@E�L��3@n�B#�!?��5z�@Q��זٿj�� ��@E�L��3@n�B#�!?��5z�@7����ٿE��l"W�@� 9��3@�I>��!?�;���@7����ٿE��l"W�@� 9��3@�I>��!?�;���@7����ٿE��l"W�@� 9��3@�I>��!?�;���@7����ٿE��l"W�@� 9��3@�I>��!?�;���@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@��Θ�ٿ�R���1�@sg����3@���ٟ�!?/���qĵ@�zȿD�ٿ��8JV�@�
�u�3@���UY�!?�m�z�@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@�X<�v�ٿ��o����@��?N�3@��N���!?������@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@Q�VW�ٿz�u9L��@�cdg��3@(�bq�!?K2�kʴ@�.UD��ٿkvv�n�@טf���3@BL��9�!?%��>\�@�.UD��ٿkvv�n�@טf���3@BL��9�!?%��>\�@�.UD��ٿkvv�n�@טf���3@BL��9�!?%��>\�@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@����ٿ�p��N�@�.v!�3@9!��q�!?������@u��X3�ٿq$����@���h�3@�E.{�!?�(�`�Ǵ@]��-��ٿ�Wo�c�@! ����3@/�S�B�!?\N;�d��@]��-��ٿ�Wo�c�@! ����3@/�S�B�!?\N;�d��@�����ٿ��K��@�S����3@�)�t��!?<�"Īִ@���<�ٿ��6s��@���ð�3@���2�!?����@���<�ٿ��6s��@���ð�3@���2�!?����@���<�ٿ��6s��@���ð�3@���2�!?����@�L�ٿb���-[�@V]�~�3@Z��:�!?ܾЅ�@�L�ٿb���-[�@V]�~�3@Z��:�!?ܾЅ�@�L�ٿb���-[�@V]�~�3@Z��:�!?ܾЅ�@�L�ٿb���-[�@V]�~�3@Z��:�!?ܾЅ�@�L�ٿb���-[�@V]�~�3@Z��:�!?ܾЅ�@�3��ٿ#ۡ�\�@Sp�z 4@��J�!?ٯU K�@�3��ٿ#ۡ�\�@Sp�z 4@��J�!?ٯU K�@�3��ٿ#ۡ�\�@Sp�z 4@��J�!?ٯU K�@�3��ٿ#ۡ�\�@Sp�z 4@��J�!?ٯU K�@r���T�ٿ���Ѓ��@ix�J�3@�L�;�!?\{M��õ@g'���ٿ�Uw��@3�n���3@���F�!?���w;�@g'���ٿ�Uw��@3�n���3@���F�!?���w;�@g'���ٿ�Uw��@3�n���3@���F�!?���w;�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��qh�ٿt���:�@�U��_�3@}"��e�!?���P�@��z��ٿ-ټ\I�@�t3v4@,��5�!?�|�l]�@����ٿ���w �@�qɦ�4@���J�!?�s��#��@����ٿ���w �@�qɦ�4@���J�!?�s��#��@����ٿ���w �@�qɦ�4@���J�!?�s��#��@����ٿ���w �@�qɦ�4@���J�!?�s��#��@����ٿ���w �@�qɦ�4@���J�!?�s��#��@����ٿ���w �@�qɦ�4@���J�!?�s��#��@5�Ӝ�ٿ���R.�@�� �4@�p�)�!?x�aiRߵ@5�Ӝ�ٿ���R.�@�� �4@�p�)�!?x�aiRߵ@5�Ӝ�ٿ���R.�@�� �4@�p�)�!?x�aiRߵ@5�Ӝ�ٿ���R.�@�� �4@�p�)�!?x�aiRߵ@�Bh�ٿ�sW[��@�<�R�	4@"G5֏!?U�>r�s�@�Q��ٿ�Jt0rp�@���o��3@���ڏ!?u� ����@�Q��ٿ�Jt0rp�@���o��3@���ڏ!?u� ����@�Q��ٿ�Jt0rp�@���o��3@���ڏ!?u� ����@q�A$��ٿ�Pٌ3�@ ���3@��A�V�!?g�r�eA�@q�A$��ٿ�Pٌ3�@ ���3@��A�V�!?g�r�eA�@q�A$��ٿ�Pٌ3�@ ���3@��A�V�!?g�r�eA�@��g@$�ٿ
�"���@�<9���3@c��+�!?-ȥ��S�@��g@$�ٿ
�"���@�<9���3@c��+�!?-ȥ��S�@��g@$�ٿ
�"���@�<9���3@c��+�!?-ȥ��S�@�x�"�ٿ0)_��N�@e�Rz�4@6�ջ�!?�L0 ؔ�@�x�"�ٿ0)_��N�@e�Rz�4@6�ջ�!?�L0 ؔ�@�x�"�ٿ0)_��N�@e�Rz�4@6�ջ�!?�L0 ؔ�@�x�"�ٿ0)_��N�@e�Rz�4@6�ջ�!?�L0 ؔ�@�]�Kٿp�t���@cB��3@�F�[�!?�<�S���@����Ԗٿ�}Oj��@�Sr�H�3@���C�!?�W�<µ@����Ԗٿ�}Oj��@�Sr�H�3@���C�!?�W�<µ@����Ԗٿ�}Oj��@�Sr�H�3@���C�!?�W�<µ@����Ԗٿ�}Oj��@�Sr�H�3@���C�!?�W�<µ@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@��B<?�ٿ@I��d�@c�TĊ�3@�+��!?6�Q��(�@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@�+&�ٿ&>:e���@�xb��3@]�P�G�!?��<��@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@Q�H��ٿ:����@٣E���3@��B�!?Gς޴@el���ٿ,w���@lB.�3@���"4�!?�Y��=Y�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@���`n�ٿh��@�2�c�3@2�O��!?Y�>�z�@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@] գ�ٿ{�U��@r�>�U�3@����k�!?)_���@"t+6ƚٿ"#���@R�Sɞ�3@���7��!?4ʤ�u��@E��!"�ٿNP
��@k�0v��3@6y_�!?�?1�@O���<�ٿ\�lq0�@H�&3T�3@d,��$�!?����
�@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@^Z����ٿ:Z�����@q�p+.�3@�bc��!?M[E���@f�̵�ٿ2n���-�@#���V�3@np�|c�!?�d����@f�̵�ٿ2n���-�@#���V�3@np�|c�!?�d����@���Zŏٿ���
�@;+��3@"+��<�!?|&K.lb�@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@Wf����ٿR/�V��@�3݇4@b��e�!?�l܉3��@~|"=�ٿ`A�I���@���t4@ ����!?l^��Ĵ@~|"=�ٿ`A�I���@���t4@ ����!?l^��Ĵ@L) �"�ٿ��az�@�3��3@'�}s�!?q��v�@L) �"�ٿ��az�@�3��3@'�}s�!?q��v�@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@SNO6�ٿ����)��@�����3@���*x�!?�8� �@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�,��ٿ6�^�>��@J�����3@,�l=,�!?(5�+�V�@�J��ٿ�(K<��@����4@�-�!?u��ߠ	�@�J��ٿ�(K<��@����4@�-�!?u��ߠ	�@�J��ٿ�(K<��@����4@�-�!?u��ߠ	�@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@m�mX"�ٿ<<.�$�@������3@`��܎�!?Q�aC�Ѵ@�-`���ٿ.35�w`�@��(�Q�3@4�i�!?Ҁ�g���@�-`���ٿ.35�w`�@��(�Q�3@4�i�!?Ҁ�g���@�-`���ٿ.35�w`�@��(�Q�3@4�i�!?Ҁ�g���@�-`���ٿ.35�w`�@��(�Q�3@4�i�!?Ҁ�g���@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@ACbÚٿ�'s�U�@��N�3@�I�p�!?�n�GS�@{좖ٿwug7q�@ �;���3@R�i*��!?��5���@{좖ٿwug7q�@ �;���3@R�i*��!?��5���@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@3܎"�ٿ������@}px]�3@�ݦ�Q�!?"�+��@�ڊ��ٿ��P�?��@����3@�P:m�!?���ѝ��@�ڊ��ٿ��P�?��@����3@�P:m�!?���ѝ��@�?����ٿM�g:�@���J�3@������!?��	PpG�@�?����ٿM�g:�@���J�3@������!?��	PpG�@�?����ٿM�g:�@���J�3@������!?��	PpG�@����ٿ������@�@���3@C�(8t�!?�hʫ0�@����ٿ������@�@���3@C�(8t�!?�hʫ0�@����ٿ������@�@���3@C�(8t�!?�hʫ0�@����ٿ������@�@���3@C�(8t�!?�hʫ0�@�����ٿ"/2=���@��L�M�3@$�p<�!?�j���z�@��枺�ٿ���ع�@�N��A�3@*��]�!?Mt��a�@��枺�ٿ���ع�@�N��A�3@*��]�!?Mt��a�@��פ��ٿ�w�jX��@�osX��3@�ixI�!?D+j�yM�@��פ��ٿ�w�jX��@�osX��3@�ixI�!?D+j�yM�@��פ��ٿ�w�jX��@�osX��3@�ixI�!?D+j�yM�@��פ��ٿ�w�jX��@�osX��3@�ixI�!?D+j�yM�@��פ��ٿ�w�jX��@�osX��3@�ixI�!?D+j�yM�@j΍vA�ٿ�Y�m��@��6�N 4@0*7G�!?��?>= �@j΍vA�ٿ�Y�m��@��6�N 4@0*7G�!?��?>= �@ٻ�n*�ٿ�O C��@��*��4@��/�!?�)��Ǵ@ٻ�n*�ٿ�O C��@��*��4@��/�!?�)��Ǵ@ٻ�n*�ٿ�O C��@��*��4@��/�!?�)��Ǵ@ٻ�n*�ٿ�O C��@��*��4@��/�!?�)��Ǵ@ٻ�n*�ٿ�O C��@��*��4@��/�!?�)��Ǵ@��j�_�ٿ��:���@�ج��3@�J�BL�!?3z̝���@��j�_�ٿ��:���@�ج��3@�J�BL�!?3z̝���@cs�ٿ2UW_�;�@����3@��D;�!?��Q��T�@Eu��ٿ����7��@�=-K��3@��WU��!?����	�@1���ٿ2b�*���@G���+�3@�t�&L�!?��K`ش@1���ٿ2b�*���@G���+�3@�t�&L�!?��K`ش@1���ٿ2b�*���@G���+�3@�t�&L�!?��K`ش@1���ٿ2b�*���@G���+�3@�t�&L�!?��K`ش@��đٿ��H�#�@Q�d�3@g=Ӏp�!?�Y^S���@M�y�ٿ1X�0�m�@N���3@U@�x�!?��@�Y�@M�y�ٿ1X�0�m�@N���3@U@�x�!?��@�Y�@�$i"�ٿ������@9��/��3@�}`�x�!?��ٷ��@�$i"�ٿ������@9��/��3@�}`�x�!?��ٷ��@M����ٿ{��S2�@\PΨW�3@�S����!?��@���@[��R��ٿ�6����@��z���3@E�$�;�!?�����t�@[��R��ٿ�6����@��z���3@E�$�;�!?�����t�@[��R��ٿ�6����@��z���3@E�$�;�!?�����t�@[��R��ٿ�6����@��z���3@E�$�;�!?�����t�@[��R��ٿ�6����@��z���3@E�$�;�!?�����t�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@�����ٿ�Nf¬�@_��{�3@T�i�B�!?�2�38n�@��݈��ٿo;�6��@��u&�3@�E���!?JOt@��݈��ٿo;�6��@��u&�3@�E���!?JOt@��݈��ٿo;�6��@��u&�3@�E���!?JOt@��݈��ٿo;�6��@��u&�3@�E���!?JOt@��݈��ٿo;�6��@��u&�3@�E���!?JOt@�e��ٿ�>����@#5j��3@�+Zq�!?w��,5�@�e��ٿ�>����@#5j��3@�+Zq�!?w��,5�@�e��ٿ�>����@#5j��3@�+Zq�!?w��,5�@�e��ٿ�>����@#5j��3@�+Zq�!?w��,5�@���C��ٿ��� �@���P �3@'���q�!?ң���5�@���C��ٿ��� �@���P �3@'���q�!?ң���5�@���C��ٿ��� �@���P �3@'���q�!?ң���5�@�~ 8��ٿ��%
;�@?���(�3@�#�^�!?��W�}f�@�~ 8��ٿ��%
;�@?���(�3@�#�^�!?��W�}f�@�~ 8��ٿ��%
;�@?���(�3@�#�^�!?��W�}f�@�~ 8��ٿ��%
;�@?���(�3@�#�^�!?��W�}f�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@�a����ٿ������@�-4��3@�/?�r�!?��?h�`�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@]Hp+q�ٿ['�����@�g7��3@;��`�!?4���'T�@:N:,�ٿ\�"ݬ�@��h��3@:���!?��Lx�@:N:,�ٿ\�"ݬ�@��h��3@:���!?��Lx�@:N:,�ٿ\�"ݬ�@��h��3@:���!?��Lx�@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@��5	K�ٿ��L�c�@kp��3@g�ʏ!?U�<�y��@�;�Q�ٿ ��h��@n�'X��3@t ��!?�g�е@�;�Q�ٿ ��h��@n�'X��3@t ��!?�g�е@�;�Q�ٿ ��h��@n�'X��3@t ��!?�g�е@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�B�Ėٿ�
��3�@���Q��3@�E��A�!?�U�5(�@�fQHE�ٿ���:
�@(��M��3@֍",�!?��۫��@�fQHE�ٿ���:
�@(��M��3@֍",�!?��۫��@�fQHE�ٿ���:
�@(��M��3@֍",�!?��۫��@re��ٿtu4;�@̧ؒ��3@rh3��!?x��p���@re��ٿtu4;�@̧ؒ��3@rh3��!?x��p���@~�e�ٿ�CC)�@C��*V�3@̉����!?�rN��@�mE���ٿ����A��@���F��3@�	4��!?�gx�6�@�mE���ٿ����A��@���F��3@�	4��!?�gx�6�@v�dժ�ٿ��eG2��@H�5��3@���+�!?�ۅ:�@v�dժ�ٿ��eG2��@H�5��3@���+�!?�ۅ:�@v�dժ�ٿ��eG2��@H�5��3@���+�!?�ۅ:�@v�dժ�ٿ��eG2��@H�5��3@���+�!?�ۅ:�@v�dժ�ٿ��eG2��@H�5��3@���+�!?�ۅ:�@6��`��ٿ�y�6���@Rәg�3@��kQ�!?5l�أ�@6��`��ٿ�y�6���@Rәg�3@��kQ�!?5l�أ�@6��`��ٿ�y�6���@Rәg�3@��kQ�!?5l�أ�@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@NT�x,�ٿ��0�1�@�n����3@(86r<�!?�=Tz���@�e3*��ٿuKc)��@O8 ��3@�xbYg�!?�契���@�e3*��ٿuKc)��@O8 ��3@�xbYg�!?�契���@�e3*��ٿuKc)��@O8 ��3@�xbYg�!?�契���@����ٿjsWX�@����3@��0#�!?p���4Y�@����ٿjsWX�@����3@��0#�!?p���4Y�@f-F�ӎٿ1����@��Y�a�3@d��$��!?�ˋx[v�@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@|,��
�ٿ
1�uؼ�@���#z4@=�͠�!?/&ܫ��@�L�$L�ٿ<���<�@["&D��3@7��g�!?-'�M�\�@�L�$L�ٿ<���<�@["&D��3@7��g�!?-'�M�\�@�L�$L�ٿ<���<�@["&D��3@7��g�!?-'�M�\�@[tP*F�ٿ������@)J�-��3@<%<Đ!?C�P��@7�c�ڕٿ|�ұ���@#>�ݕ�3@h�s�!?�ܷ���@��я�ٿ�)���]�@PG�aE�3@�#�T��!?�q��m��@��я�ٿ�)���]�@PG�aE�3@�#�T��!?�q��m��@��я�ٿ�)���]�@PG�aE�3@�#�T��!?�q��m��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@!�&8��ٿ�7)s���@��弎�3@�<��Z�!?I��-��@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@���T��ٿ��^Gc�@�3��k�3@��?�g�!?�5�ۺK�@kXT��ٿ��c`u�@橛���3@�i�~��!?)Ġ�i�@kXT��ٿ��c`u�@橛���3@�i�~��!?)Ġ�i�@kXT��ٿ��c`u�@橛���3@�i�~��!?)Ġ�i�@$=�W�ٿrE��ii�@���	�3@f��.�!?n��I`�@$=�W�ٿrE��ii�@���	�3@f��.�!?n��I`�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@"���ٿ�m�{��@Lb�y�3@>����!?�7[zr�@�GG�ړٿ�5X[�P�@����3@|��f�!?v�X�7�@�xë�ٿ�p�mav�@� ��n�3@^s�:=�!?vh�a�[�@ڏ�y��ٿs��'��@5΢�X�3@�	G_9�!?2�#荕�@ڏ�y��ٿs��'��@5΢�X�3@�	G_9�!?2�#荕�@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@v��U��ٿ@�v!n��@�f�E��3@�Ӧi�!?�+W��@m�l��ٿs���	��@~$����3@�g��!?xꚤ'��@�H�R�ٿ����@��z���3@v����!?���S�@��Y�ٿ��*���@�7� ��3@��%�!?{DS'��@��Y�ٿ��*���@�7� ��3@��%�!?{DS'��@��Y�ٿ��*���@�7� ��3@��%�!?{DS'��@��
��ٿb�Oi/
�@r�y��3@Y��_�!?�]�n�ϴ@��
��ٿb�Oi/
�@r�y��3@Y��_�!?�]�n�ϴ@��
��ٿb�Oi/
�@r�y��3@Y��_�!?�]�n�ϴ@��
��ٿb�Oi/
�@r�y��3@Y��_�!?�]�n�ϴ@��
��ٿb�Oi/
�@r�y��3@Y��_�!?�]�n�ϴ@���g �ٿ����@���3@�[�H�!?����+�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@0���ٿ8����@��f��3@�pFc�!?��C�(�@"���ٿ�d��@J?yY�3@A���!?G�ei�ʴ@"���ٿ�d��@J?yY�3@A���!?G�ei�ʴ@"���ٿ�d��@J?yY�3@A���!?G�ei�ʴ@"���ٿ�d��@J?yY�3@A���!?G�ei�ʴ@0暓 �ٿ|u�r<�@��MT7�3@
Uo��!?I�ϴ@�%A�ٿ���e�@f�3���3@��9�a�!?2����۴@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@Q����ٿˮ��X�@�����3@�;J9A�!?�XA�]�@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@��3�ٿ�˗�9��@Z쁄��3@���!?����G��@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@���y.�ٿ m����@����3@�q���!?Youg���@H���җٿA /�]�@���\�3@8)�TT�!?H%�Zx�@H���җٿA /�]�@���\�3@8)�TT�!?H%�Zx�@H���җٿA /�]�@���\�3@8)�TT�!?H%�Zx�@����іٿ�����@����3@�@���!?�c�<��@����іٿ�����@����3@�@���!?�c�<��@oh(h��ٿͼ� ��@�@D.�3@��~�!?�H�	���@oh(h��ٿͼ� ��@�@D.�3@��~�!?�H�	���@oh(h��ٿͼ� ��@�@D.�3@��~�!?�H�	���@oh(h��ٿͼ� ��@�@D.�3@��~�!?�H�	���@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�_Q'[�ٿ0#H�i�@�f���3@��(Ð!?N���?�@�}e�ٿۨX%q�@-W�~I�3@oHS��!?���&a�@�}e�ٿۨX%q�@-W�~I�3@oHS��!?���&a�@��̕ٿ=a:�S��@����4@���~�!?�45��˵@��̕ٿ=a:�S��@����4@���~�!?�45��˵@��̕ٿ=a:�S��@����4@���~�!?�45��˵@��̕ٿ=a:�S��@����4@���~�!?�45��˵@��̕ٿ=a:�S��@����4@���~�!?�45��˵@��̕ٿ=a:�S��@����4@���~�!?�45��˵@���țٿY]��@�;�O�4@��%ɰ�!?4B}�@�',��ٿ��e����@������3@Z�$�!?he�obԴ@�',��ٿ��e����@������3@Z�$�!?he�obԴ@1��P�ٿ���J�@���4�3@n$[��!?ϥ��ô@1��P�ٿ���J�@���4�3@n$[��!?ϥ��ô@1��P�ٿ���J�@���4�3@n$[��!?ϥ��ô@Ip,Ѭ�ٿ�p�~�@�6~6�3@|�Z
�!?�?5�3o�@Ip,Ѭ�ٿ�p�~�@�6~6�3@|�Z
�!?�?5�3o�@Ip,Ѭ�ٿ�p�~�@�6~6�3@|�Z
�!?�?5�3o�@Ip,Ѭ�ٿ�p�~�@�6~6�3@|�Z
�!?�?5�3o�@Ip,Ѭ�ٿ�p�~�@�6~6�3@|�Z
�!?�?5�3o�@�ų��ٿ��<.�I�@��1=�3@)��<Y�!?�����մ@��9�ٿ�������@���t��3@7gg?n�!?CY���@��9�ٿ�������@���t��3@7gg?n�!?CY���@v6�ٿ�p��1�@�PU 4@G��aU�!?��t�!�@v6�ٿ�p��1�@�PU 4@G��aU�!?��t�!�@v6�ٿ�p��1�@�PU 4@G��aU�!?��t�!�@v6�ٿ�p��1�@�PU 4@G��aU�!?��t�!�@�C8D$�ٿ�PC��@|�i��3@`����!?��%�F��@�C8D$�ٿ�PC��@|�i��3@`����!?��%�F��@kH�ϔٿ@ Z��@���U�3@���@�!?�r��@kH�ϔٿ@ Z��@���U�3@���@�!?�r��@kH�ϔٿ@ Z��@���U�3@���@�!?�r��@kH�ϔٿ@ Z��@���U�3@���@�!?�r��@���a�ٿO����@����L�3@�H����!?�S J�@���a�ٿO����@����L�3@�H����!?�S J�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�K�k6�ٿD)H�D�@��3�I�3@�[��#�!?�f�v�e�@�D�Kܙٿ/CWn�@ta%b��3@1�oȁ!?����H�@�D�Kܙٿ/CWn�@ta%b��3@1�oȁ!?����H�@�:�Y�ٿ��� ��@UD�Y|�3@�d?�-�!?��z	%�@�:�Y�ٿ��� ��@UD�Y|�3@�d?�-�!?��z	%�@�q��ǖٿ	���@�,��_�3@�T*���!?�MU��D�@�q��ǖٿ	���@�,��_�3@�T*���!?�MU��D�@�q��ǖٿ	���@�,��_�3@�T*���!?�MU��D�@�q��ǖٿ	���@�,��_�3@�T*���!?�MU��D�@�q��ǖٿ	���@�,��_�3@�T*���!?�MU��D�@/�;3�ٿ�ū}��@�p��n�3@{�T�@�!?�y��ȴ@/�;3�ٿ�ū}��@�p��n�3@{�T�@�!?�y��ȴ@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@��]>Ӗٿ;*��y�@{�j'��3@�(�n�!?l�X�5�@m��p��ٿ���q���@��E�4@�j�A4�!?׿+�[w�@m��p��ٿ���q���@��E�4@�j�A4�!?׿+�[w�@m��p��ٿ���q���@��E�4@�j�A4�!?׿+�[w�@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@�&�z��ٿs-�| ��@���3�3@��+�c�!?�8���´@"`�Ƙٿz��pV�@��Tχ4@�`p�!?�`Ɋn۴@"`�Ƙٿz��pV�@��Tχ4@�`p�!?�`Ɋn۴@"`�Ƙٿz��pV�@��Tχ4@�`p�!?�`Ɋn۴@y�*��ٿ|��ܭ\�@���4@����7�!?b���@y�*��ٿ|��ܭ\�@���4@����7�!?b���@�A��	�ٿ'a[��F�@����4@��f6Y�!?����Q��@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@��A�Ӕٿ\�R��@K�A��4@_��f�!?�:�]Q�@p�;h�ٿ"����@�O����3@� T%D�!?������@p�;h�ٿ"����@�O����3@� T%D�!?������@p�;h�ٿ"����@�O����3@� T%D�!?������@����/�ٿ�/��R��@�G��3@�+E^��!?��|{��@=mT��ٿU����@��OPl�3@F��>�!?�d��B�@
4X�'�ٿ̪Y�*h�@Y1M !�3@;	lQ�!?����@
4X�'�ٿ̪Y�*h�@Y1M !�3@;	lQ�!?����@
4X�'�ٿ̪Y�*h�@Y1M !�3@;	lQ�!?����@� �lƌٿ��r�C��@�s����3@�C�c�!?�[L��@�ά��ٿH�HE���@p�/;�3@�8�.�!?�(A'�@�ά��ٿH�HE���@p�/;�3@�8�.�!?�(A'�@�ά��ٿH�HE���@p�/;�3@�8�.�!?�(A'�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@o�s��ٿU��n��@�����3@�Ϝ�w�!?`��۱�@ˇ(ʓٿ��r�q�@k[r��3@�`�칐!?����C�@x�b2�ٿ�#(�p�@�u�9(�3@�0c[�!?�"� ��@K��(-�ٿ�����!�@	��B�3@0���!?U7��s��@K��(-�ٿ�����!�@	��B�3@0���!?U7��s��@ ���ٿa�jN�{�@T��V�3@��A�u�!?�V�P��@ ���ٿa�jN�{�@T��V�3@��A�u�!?�V�P��@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�iޏ�ٿ��~N��@���\b�3@���ʐ!?u�7i�@�#�m��ٿ������@;����3@'����!?��W��@�#�m��ٿ������@;����3@'����!?��W��@�#�m��ٿ������@;����3@'����!?��W��@By�3��ٿ'l�,[)�@�`��)�3@C���(�!?��B#�@By�3��ٿ'l�,[)�@�`��)�3@C���(�!?��B#�@By�3��ٿ'l�,[)�@�`��)�3@C���(�!?��B#�@��xD�ٿ�j&��Z�@�����3@	C�1�!?@ƳH�C�@��xD�ٿ�j&��Z�@�����3@	C�1�!?@ƳH�C�@��xD�ٿ�j&��Z�@�����3@	C�1�!?@ƳH�C�@��(�ٿ��٥u��@qO�f��3@P�Ca��!?#�10�&�@	8|��ٿ���7m�@���7{�3@34
ӏ!?zuN�M�@	8|��ٿ���7m�@���7{�3@34
ӏ!?zuN�M�@	8|��ٿ���7m�@���7{�3@34
ӏ!?zuN�M�@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@�r�C��ٿ�[A	C�@�Kӽ�3@�a�U��!?��ة���@Y¬�2�ٿqG�a�@�;9�O�3@�`���!?��U��@Y¬�2�ٿqG�a�@�;9�O�3@�`���!?��U��@Y¬�2�ٿqG�a�@�;9�O�3@�`���!?��U��@Y¬�2�ٿqG�a�@�;9�O�3@�`���!?��U��@Y¬�2�ٿqG�a�@�;9�O�3@�`���!?��U��@b<���ٿ�e[�'I�@(&�Ǥ�3@�fi!?�z�XM��@b<���ٿ�e[�'I�@(&�Ǥ�3@�fi!?�z�XM��@���z�ٿbX��/�@�g��4@��C�$�!?�ȭm���@���z�ٿbX��/�@�g��4@��C�$�!?�ȭm���@���z�ٿbX��/�@�g��4@��C�$�!?�ȭm���@���z�ٿbX��/�@�g��4@��C�$�!?�ȭm���@ih�p��ٿ�8��@.���4@�1�A\�!?P��f� �@C܊x�ٿAz}iR�@)}��3@�P��!?���'v�@C܊x�ٿAz}iR�@)}��3@�P��!?���'v�@C܊x�ٿAz}iR�@)}��3@�P��!?���'v�@C܊x�ٿAz}iR�@)}��3@�P��!?���'v�@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@�_��ٿ��7K���@^�ɐ��3@�Yϸ��!?�Y��;��@Z���ٿOA=����@��v���3@�RZϐ!?ݳT$�'�@�gz1N�ٿ�Iq�o�@th�{�3@���Ő!?�F)J��@�gz1N�ٿ�Iq�o�@th�{�3@���Ő!?�F)J��@��b��ٿ�A6*3�@I�D:2�3@"�� �!?�)�SFq�@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@�8.K�ٿ�pco]5�@��p%�3@^�.���!?�ʯ���@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@d^��c�ٿ����@9@�D4@|5x-�!?=����@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@+��t�ٿ�^���&�@�Y��04@�O�$q�!?�+�՜Ѵ@X��#�ٿ��R!��@[�j��3@L��ZS�!?���vv�@X��#�ٿ��R!��@[�j��3@L��ZS�!?���vv�@X��#�ٿ��R!��@[�j��3@L��ZS�!?���vv�@X��#�ٿ��R!��@[�j��3@L��ZS�!?���vv�@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@H+�թ�ٿ+O�&V�@h|���3@�BAZY�!?�/�Jڴ@)x�ޓٿP����@G� "�3@�H��&�!?��Q�_�@�ʊ���ٿ��J�5��@wZ/��3@�EӘ�!?w1>2��@��ɦ�ٿڐ��Y7�@4���4�3@��i�!?�H�¾6�@��ɦ�ٿڐ��Y7�@4���4�3@��i�!?�H�¾6�@��ɦ�ٿڐ��Y7�@4���4�3@��i�!?�H�¾6�@}��z�ٿ��j8M�@5�z�N�3@�ٚ�׏!?��`�#�@}��z�ٿ��j8M�@5�z�N�3@�ٚ�׏!?��`�#�@}��z�ٿ��j8M�@5�z�N�3@�ٚ�׏!?��`�#�@}��z�ٿ��j8M�@5�z�N�3@�ٚ�׏!?��`�#�@}��z�ٿ��j8M�@5�z�N�3@�ٚ�׏!?��`�#�@��b	�ٿ;�ֈ��@��`ӷ�3@o�*�!?&��%�N�@��]=\�ٿ�Ϯ�=�@0G���3@@#��!?�^Eڵx�@��]=\�ٿ�Ϯ�=�@0G���3@@#��!?�^Eڵx�@:��<�ٿ/��@p��@�U�1r4@��zg��!?)�����@�����ٿ��.S��@�����3@�&�(�!?QO>V��@�����ٿ��.S��@�����3@�&�(�!?QO>V��@�����ٿ��.S��@�����3@�&�(�!?QO>V��@�����ٿ��.S��@�����3@�&�(�!?QO>V��@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@���=1�ٿ���K���@�Sk/h�3@�O���!?m�>�ɴ@��UB�ٿ������@Ԅ�M �3@?	O���!?��]���@��UB�ٿ������@Ԅ�M �3@?	O���!?��]���@�t��L�ٿ����t�@X����3@v��$�!?b1���@�t��L�ٿ����t�@X����3@v��$�!?b1���@�t��L�ٿ����t�@X����3@v��$�!?b1���@�t��L�ٿ����t�@X����3@v��$�!?b1���@��Ar1�ٿ����-<�@��L{�3@G�m��!?r�-��@��Ar1�ٿ����-<�@��L{�3@G�m��!?r�-��@��Ar1�ٿ����-<�@��L{�3@G�m��!?r�-��@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@��4dĕٿM�,�!�@H�p�&�3@�LJH�!?}S��5�@���n�ٿ���X�@��_���3@Mǒ\�!?��>/��@���n�ٿ���X�@��_���3@Mǒ\�!?��>/��@���n�ٿ���X�@��_���3@Mǒ\�!?��>/��@�K��ǔٿ�_˗��@��l��3@���!?��'����@�K��ǔٿ�_˗��@��l��3@���!?��'����@�K��ǔٿ�_˗��@��l��3@���!?��'����@�K��ǔٿ�_˗��@��l��3@���!?��'����@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@%s;�n�ٿ�o�o'�@���!��3@*�8#�!?HYG��ڴ@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@��s���ٿ��@6S�@��N�X�3@� �mY�!?�$�� +�@���A�ٿ�񦼑��@3!G$C�3@u��k�!?x~r�@���A�ٿ�񦼑��@3!G$C�3@u��k�!?x~r�@���A�ٿ�񦼑��@3!G$C�3@u��k�!?x~r�@���A�ٿ�񦼑��@3!G$C�3@u��k�!?x~r�@P7pƖٿ��26I��@��k���3@�F� ��!?͸,��@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@2���ٿ��ٗȏ�@������3@��(j�!?��c�-�@m�G�זٿ������@u�߶�3@a�EAA�!?� ����@m�G�זٿ������@u�߶�3@a�EAA�!?� ����@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@�7��ٿ��s(h}�@�X�2��3@�"6�!?�a���>�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@͑���ٿ�A"<ǁ�@0r��3@a�E�5�!?\�[�1$�@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@�L�X�ٿ� g��@���GU�3@֝�8q�!?m��?᪵@��@�:�ٿr��5��@s��3�3@ᰃ��!?�9�M�&�@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@v�K?{�ٿǤ[���@����3@o)�oF�!?��B��@��츛ٿm�3�X�@� A�3@��`(��!?�k�+��@-���1�ٿ�(��_�@dW�P�3@U9�p�!?琜���@-���1�ٿ�(��_�@dW�P�3@U9�p�!?琜���@�G|=��ٿT&S⨪�@�[^��3@=���t�!?�y=|"��@�G|=��ٿT&S⨪�@�[^��3@=���t�!?�y=|"��@�G|=��ٿT&S⨪�@�[^��3@=���t�!?�y=|"��@�G|=��ٿT&S⨪�@�[^��3@=���t�!?�y=|"��@P]�c�ٿ�a7O���@�w�R�3@4uM�R�!?�-s�&�@	�ٿ�k�=�K�@qT0��3@�rҙP�!?����N%�@	�ٿ�k�=�K�@qT0��3@�rҙP�!?����N%�@	�ٿ�k�=�K�@qT0��3@�rҙP�!?����N%�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@���L �ٿ����d��@�ak���3@[¿ꖐ!?g�@�Z)�@��$"Z�ٿ��7���@�z��3@���a�!?���|&�@��$"Z�ٿ��7���@�z��3@���a�!?���|&�@��$"Z�ٿ��7���@�z��3@���a�!?���|&�@��$"Z�ٿ��7���@�z��3@���a�!?���|&�@+t���ٿ	 ��!�@��%���3@�� g�!?X��O��@+t���ٿ	 ��!�@��%���3@�� g�!?X��O��@`Nu��ٿٗ�x,�@���kF�3@�6]���!?r	�B+z�@`Nu��ٿٗ�x,�@���kF�3@�6]���!?r	�B+z�@`Nu��ٿٗ�x,�@���kF�3@�6]���!?r	�B+z�@`Nu��ٿٗ�x,�@���kF�3@�6]���!?r	�B+z�@`Nu��ٿٗ�x,�@���kF�3@�6]���!?r	�B+z�@?�.�ٿrܶ0���@�=����3@��Lf�!?D�*�&�@?�.�ٿrܶ0���@�=����3@��Lf�!?D�*�&�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�PV���ٿ���RL�@k��A,�3@O�T��!?Q�*1�@�l�ėٿ���ԟ=�@Ԓ���3@���=p�!?hsa�!�@�,��&�ٿ��
7�@^c���3@��B�!?�_�Ф�@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�ء/ٝٿ�ڀ����@���ZK�3@��v<�!?U\�׵@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�C�/"�ٿTG:�I��@R%^��3@m���!?������@�W�Q�ٿ{	e��D�@'`b�|�3@�Ys̅�!?��)��@�W�Q�ٿ{	e��D�@'`b�|�3@�Ys̅�!?��)��@�W�Q�ٿ{	e��D�@'`b�|�3@�Ys̅�!?��)��@�W�Q�ٿ{	e��D�@'`b�|�3@�Ys̅�!?��)��@�Vm��ٿ	b�ȵ��@we����3@�8�V4�!?$v���ش@�Vm��ٿ	b�ȵ��@we����3@�8�V4�!?$v���ش@��9���ٿ���6���@D���3@n\JF��!?/E���@��9���ٿ���6���@D���3@n\JF��!?/E���@��9���ٿ���6���@D���3@n\JF��!?/E���@��9���ٿ���6���@D���3@n\JF��!?/E���@��9���ٿ���6���@D���3@n\JF��!?/E���@��9���ٿ���6���@D���3@n\JF��!?/E���@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@�֝�˕ٿ)�B���@'���3@.�J�!?:K�GV)�@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@|ᖷ��ٿ(��O�@�W��	�3@l�G�!?,�}���@x��!M�ٿP]�t���@3U�g:�3@�Ţ4�!?��7�ϴ@x��!M�ٿP]�t���@3U�g:�3@�Ţ4�!?��7�ϴ@x��!M�ٿP]�t���@3U�g:�3@�Ţ4�!?��7�ϴ@x��!M�ٿP]�t���@3U�g:�3@�Ţ4�!?��7�ϴ@�DK�ٿ�Y�D�@�&��3@��Uc�!?0pO*>��@S�ԶՔٿ�]!���@��W`��3@���b�!?��wW�@S�ԶՔٿ�]!���@��W`��3@���b�!?��wW�@S�ԶՔٿ�]!���@��W`��3@���b�!?��wW�@q�ě�ٿ����0�@�Q�3W�3@�j�Y�!?���p�@�?��.�ٿB�
����@�!	n�3@"�E�x�!?�f���N�@�?��.�ٿB�
����@�!	n�3@"�E�x�!?�f���N�@�?��.�ٿB�
����@�!	n�3@"�E�x�!?�f���N�@�?��.�ٿB�
����@�!	n�3@"�E�x�!?�f���N�@�$��/�ٿ��o��@�mHx��3@3�/ː!?��6��W�@�$��/�ٿ��o��@�mHx��3@3�/ː!?��6��W�@�$��/�ٿ��o��@�mHx��3@3�/ː!?��6��W�@�$��/�ٿ��o��@�mHx��3@3�/ː!?��6��W�@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@�@7$��ٿҞJ@��@W�|j�3@K�=��!?t�����@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@��L���ٿ��FxR'�@.*J�5�3@�pwzn�!?r=�+�R�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@���ٿm�4=��@�#B�@�3@�`T�!?��і�@��a�c�ٿ���F��@�(@�3@��`T�!?��nw�:�@��a�c�ٿ���F��@�(@�3@��`T�!?��nw�:�@��a�c�ٿ���F��@�(@�3@��`T�!?��nw�:�@��a�c�ٿ���F��@�(@�3@��`T�!?��nw�:�@��{xʔٿ�:K���@������3@f	�T�!?���� �@��{xʔٿ�:K���@������3@f	�T�!?���� �@��{xʔٿ�:K���@������3@f	�T�!?���� �@��{xʔٿ�:K���@������3@f	�T�!?���� �@��{xʔٿ�:K���@������3@f	�T�!?���� �@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�ҿ�@�ٿ.h�i��@x�B���3@��s�'�!?�1�>�@�$V�ٿ�O��@�Sv��3@�O���!?��Mkm�@�$V�ٿ�O��@�Sv��3@�O���!?��Mkm�@�$V�ٿ�O��@�Sv��3@�O���!?��Mkm�@�$V�ٿ�O��@�Sv��3@�O���!?��Mkm�@�-��ٿ1@>~��@�4:>��3@b)�B�!?��Sq��@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@�ZZG�ٿN��G?�@/�����3@��P��!?Z".�w�@��|ˑٿ��l\�0�@��<���3@l0��=�!?\��Tc}�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@/e��y�ٿ`mP=��@�n?i�3@��+�I�!?�)D�c�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@����ٿ�B]�O�@���f{�3@l���B�!?�-��7�@�&b���ٿ߉��S��@�
�r�3@y�4{-�!?m)��#�@�-57�ٿ�2�BG~�@}��ue�3@5,�E��!?ȕ
����@�-57�ٿ�2�BG~�@}��ue�3@5,�E��!?ȕ
����@�-57�ٿ�2�BG~�@}��ue�3@5,�E��!?ȕ
����@�d�G*�ٿ���4�@���&��3@%(	z�!?,?�콎�@|���ٿUb+\!�@�n[��3@M|c!^�!?s��xM��@|���ٿUb+\!�@�n[��3@M|c!^�!?s��xM��@�H���ٿ�q���P�@"/�z�3@$�}��!?8������@�H���ٿ�q���P�@"/�z�3@$�}��!?8������@����ٿ�׀Ο�@,R�y�3@Y�[��!?;�B9N��@����ٿ�׀Ο�@,R�y�3@Y�[��!?;�B9N��@�L�*˕ٿ!����G�@(��N��3@�g_I��!?r�`PqM�@�&4`ݕٿW��i��@���6�3@f y�a�!?U�)oM	�@�y�j�ٿ�D��h��@_\u
�3@@*Ç�!?�D5��$�@�y�j�ٿ�D��h��@_\u
�3@@*Ç�!?�D5��$�@J����ٿ2	S�M.�@��V��3@&y��h�!?~����!�@J����ٿ2	S�M.�@��V��3@&y��h�!?~����!�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@�����ٿA��Mg�@%LG��4@��t�!?T6��n�@!90�ٿI_��"C�@E�LV=�3@i!X�f�!?͇�ɵ@!90�ٿI_��"C�@E�LV=�3@i!X�f�!?͇�ɵ@��<�ٿ�_s%B�@����M�3@��j��!?����j�@��<�ٿ�_s%B�@����M�3@��j��!?����j�@��<�ٿ�_s%B�@����M�3@��j��!?����j�@1�5,�ٿ{t����@����
�3@٘Rΐ!?֘Yu��@1�5,�ٿ{t����@����
�3@٘Rΐ!?֘Yu��@1�5,�ٿ{t����@����
�3@٘Rΐ!?֘Yu��@1�5,�ٿ{t����@����
�3@٘Rΐ!?֘Yu��@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@�:_�ٿf�tO���@s�C���3@4@�V��!?Up
�F>�@~9m�"�ٿ����8��@Op�)��3@y�&�c�!?�1}��)�@~9m�"�ٿ����8��@Op�)��3@y�&�c�!?�1}��)�@~9m�"�ٿ����8��@Op�)��3@y�&�c�!?�1}��)�@~9m�"�ٿ����8��@Op�)��3@y�&�c�!?�1}��)�@ҧ51�ٿ� ���H�@�J#�3@vN����!?�.lS�@ҧ51�ٿ� ���H�@�J#�3@vN����!?�.lS�@ҧ51�ٿ� ���H�@�J#�3@vN����!?�.lS�@ҧ51�ٿ� ���H�@�J#�3@vN����!?�.lS�@ҧ51�ٿ� ���H�@�J#�3@vN����!?�.lS�@q�g��ٿ�F�!��@(��8�3@���n�!?�=���@q�g��ٿ�F�!��@(��8�3@���n�!?�=���@�x�+,�ٿ�����@�%�V�3@k�3��!?"�k��@�x�+,�ٿ�����@�%�V�3@k�3��!?"�k��@�x�+,�ٿ�����@�%�V�3@k�3��!?"�k��@}���ٿ�B~��@1����3@�B�!?w��`^�@}���ٿ�B~��@1����3@�B�!?w��`^�@}���ٿ�B~��@1����3@�B�!?w��`^�@}���ٿ�B~��@1����3@�B�!?w��`^�@}���ٿ�B~��@1����3@�B�!?w��`^�@}���ٿ�B~��@1����3@�B�!?w��`^�@��P��ٿ�ǅ��j�@�>����3@��d6��!?3_U�&�@��P��ٿ�ǅ��j�@�>����3@��d6��!?3_U�&�@��P��ٿ�ǅ��j�@�>����3@��d6��!?3_U�&�@��P��ٿ�ǅ��j�@�>����3@��d6��!?3_U�&�@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@ed����ٿ~���
Y�@��V֙�3@ْ���!?m����@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@��⛱�ٿ���"~�@��(�y�3@��O�!?��3?���@�X���ٿC����l�@Kz���3@g��DZ�!?�-N=�5�@w_����ٿ/����w�@b��a��3@E�!?{0���r�@w_����ٿ/����w�@b��a��3@E�!?{0���r�@w_����ٿ/����w�@b��a��3@E�!?{0���r�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@�}y�ٿ;�eIm��@6$
 ��3@`�(i�!?:�ŋ�@C�5�ٿ�!ӱh>�@1�xV�3@B6S�E�!?#b&��@����ٿj�!��@�D�X�3@�%�Y�!?%���e�@(UP�ٿ	�)�N�@8���3@�IdgY�!?V��q��@(UP�ٿ	�)�N�@8���3@�IdgY�!?V��q��@(UP�ٿ	�)�N�@8���3@�IdgY�!?V��q��@z�+���ٿ��6��@����Y�3@���!�!?	��0�@7�+��ٿ�D���@������3@�����!?���	��@2�U�W�ٿ�8��ߕ�@n/\�H�3@R�#��!?���@2�U�W�ٿ�8��ߕ�@n/\�H�3@R�#��!?���@2�U�W�ٿ�8��ߕ�@n/\�H�3@R�#��!?���@jtv@�ٿ�M����@n�=�3@�/v;+�!? � |���@jtv@�ٿ�M����@n�=�3@�/v;+�!? � |���@jtv@�ٿ�M����@n�=�3@�/v;+�!? � |���@jtv@�ٿ�M����@n�=�3@�/v;+�!? � |���@jtv@�ٿ�M����@n�=�3@�/v;+�!? � |���@I�2h��ٿ�>B��J�@�k"��3@(±Y�!?�꼌�̵@��k���ٿt�mP#��@̦�o`�3@&)�2I�!?ͯ��L��@��k���ٿt�mP#��@̦�o`�3@&)�2I�!?ͯ��L��@ӗu�ٿ	"7�}\�@�w?���3@�U�ˏ!?�."���@ӗu�ٿ	"7�}\�@�w?���3@�U�ˏ!?�."���@ p;�ٿ���ư�@��>��3@\5 �!?��C��G�@{�U��ٿ����c�@������3@����@�!?άbzD�@{�U��ٿ����c�@������3@����@�!?άbzD�@{�U��ٿ����c�@������3@����@�!?άbzD�@mO��3�ٿ��cs�@�ӣ��3@���Ώ!?m�K���@mO��3�ٿ��cs�@�ӣ��3@���Ώ!?m�K���@mO��3�ٿ��cs�@�ӣ��3@���Ώ!?m�K���@��խ�ٿ����@gy�r��3@Z�,n@�!?'���­�@��խ�ٿ����@gy�r��3@Z�,n@�!?'���­�@��խ�ٿ����@gy�r��3@Z�,n@�!?'���­�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@��pn�ٿ�m��K�@b�!�f�3@b�g�!?�uJ�`/�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@=��H�ٿ�����%�@�Q���3@¿�w��!?��^�@d.'�יٿD�-.a�@Q1S�3@
K����!?��Gh&Ѵ@d.'�יٿD�-.a�@Q1S�3@
K����!?��Gh&Ѵ@d.'�יٿD�-.a�@Q1S�3@
K����!?��Gh&Ѵ@���ҟ�ٿ���)��@�Ӭr��3@
�&�Y�!?�OY:5�@�T
�N�ٿD" ys�@떭U��3@��S/<�!?x���Z�@�T
�N�ٿD" ys�@떭U��3@��S/<�!?x���Z�@�T
�N�ٿD" ys�@떭U��3@��S/<�!?x���Z�@�T
�N�ٿD" ys�@떭U��3@��S/<�!?x���Z�@�T
�N�ٿD" ys�@떭U��3@��S/<�!?x���Z�@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@r�B�ٿ��� ī�@��{-��3@AbO�B�!?��豴@Ew^�ٿ�j����@�,=�3@���B�!? A(0��@Ew^�ٿ�j����@�,=�3@���B�!? A(0��@Ew^�ٿ�j����@�,=�3@���B�!? A(0��@Ew^�ٿ�j����@�,=�3@���B�!? A(0��@Ew^�ٿ�j����@�,=�3@���B�!? A(0��@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@.pTٿ�pG�H�@i�cy4@������!?l�Eִܼ@�����ٿZ&c��@����4@$SPXB�!?�%��@�*�ѝ�ٿI�,�@Q},G��3@���h��!?�{�^}<�@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��h̗ٿ�EGn3%�@l06մ�3@�|�!?wۃ���@��,�ٿI�����@��(�{�3@u�E��!?�hwUt�@��,�ٿI�����@��(�{�3@u�E��!?�hwUt�@>��̛�ٿS(��@������3@#ۗ,o�!?P���Ch�@>��̛�ٿS(��@������3@#ۗ,o�!?P���Ch�@>��̛�ٿS(��@������3@#ۗ,o�!?P���Ch�@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@I�I�ٿ�KG����@ඪ/��3@�{=�l�!?j�\g���@��'WQ�ٿp�ۅ�@�KH��3@�l7~�!?��xu�@��'WQ�ٿp�ۅ�@�KH��3@�l7~�!?��xu�@�r,�^�ٿ�����@���"�3@�L�E�!?��P.�@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@w�~=�ٿ#]eF/�@yE����3@�z�v�!?��NR��@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@05�o�ٿ�c��8:�@z���3@kc�,6�!?�2���ƴ@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@���3h�ٿOn4��@��p"V�3@`Hs�9�!?p��q~�@۷�ٿ�Q��xQ�@�]]UK�3@�!!{��!?7��@�j11�ٿ��x.�@+O�R�3@��>�!?���g�@�j11�ٿ��x.�@+O�R�3@��>�!?���g�@�0�m$�ٿ���3��@�}�kK4@�����!?K����ٴ@���ڸ�ٿ��Q!k�@Cy�5�3@�=��C�!?Vùy��@���ڸ�ٿ��Q!k�@Cy�5�3@�=��C�!?Vùy��@���ڸ�ٿ��Q!k�@Cy�5�3@�=��C�!?Vùy��@���ڸ�ٿ��Q!k�@Cy�5�3@�=��C�!?Vùy��@���ڸ�ٿ��Q!k�@Cy�5�3@�=��C�!?Vùy��@�ì�ٿW��>��@�6A���3@H� O�!?�[�~��@�ì�ٿW��>��@�6A���3@H� O�!?�[�~��@�ì�ٿW��>��@�6A���3@H� O�!?�[�~��@�ì�ٿW��>��@�6A���3@H� O�!?�[�~��@�ì�ٿW��>��@�6A���3@H� O�!?�[�~��@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@���e�ٿ�F��?��@�Q���3@��>*�!?������@��Y��ٿ�'�h��@	܁��3@�����!?%��/�@��Y��ٿ�'�h��@	܁��3@�����!?%��/�@��Y��ٿ�'�h��@	܁��3@�����!?%��/�@@-/���ٿ�Nٞή�@�c.,��3@��gZ\�!?:9��lX�@@-/���ٿ�Nٞή�@�c.,��3@��gZ\�!?:9��lX�@@-/���ٿ�Nٞή�@�c.,��3@��gZ\�!?:9��lX�@�Acx��ٿ�q�M/�@4М$G�3@-I��V�!?���`���@�Acx��ٿ�q�M/�@4М$G�3@-I��V�!?���`���@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@����ɝٿ����&�@$;�Ǳ4@��{���!?�H$�� �@��9�ʎٿB.wNx�@��0�4@�D�^�!?������@��PF�ٿ�E��f�@݁|�4@�_�;\�!? �� Y��@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@ڨ��=�ٿB�e]���@����3@L��KN�!?����䡴@�	��Ȓٿ%o�^h��@7��k��3@#��W�!?�1��	u�@�	��Ȓٿ%o�^h��@7��k��3@#��W�!?�1��	u�@�	��Ȓٿ%o�^h��@7��k��3@#��W�!?�1��	u�@�	��Ȓٿ%o�^h��@7��k��3@#��W�!?�1��	u�@�	��Ȓٿ%o�^h��@7��k��3@#��W�!?�1��	u�@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@�M]'�ٿu���v��@Ѭ�to�3@+Β�!?z����@#�3�ٿ�r��@p�����3@N�Q�o�!?��/i��@#�3�ٿ�r��@p�����3@N�Q�o�!?��/i��@#�3�ٿ�r��@p�����3@N�Q�o�!?��/i��@#�3�ٿ�r��@p�����3@N�Q�o�!?��/i��@�����ٿߍ�2��@c��:�3@u&>�N�!?��؛2:�@�����ٿߍ�2��@c��:�3@u&>�N�!?��؛2:�@�����ٿߍ�2��@c��:�3@u&>�N�!?��؛2:�@�����ٿߍ�2��@c��:�3@u&>�N�!?��؛2:�@�����ٿߍ�2��@c��:�3@u&>�N�!?��؛2:�@�``)��ٿ�mH�$�@EU����3@��l�!?a�8�Ƶ@�``)��ٿ�mH�$�@EU����3@��l�!?a�8�Ƶ@�``)��ٿ�mH�$�@EU����3@��l�!?a�8�Ƶ@�``)��ٿ�mH�$�@EU����3@��l�!?a�8�Ƶ@�``)��ٿ�mH�$�@EU����3@��l�!?a�8�Ƶ@�Q�A�ٿ��ƽ$��@�a���3@#��A��!?h�[Z��@�Q�A�ٿ��ƽ$��@�a���3@#��A��!?h�[Z��@����͐ٿ�@H|�@��B��3@�wJ��!?�'��B��@����͐ٿ�@H|�@��B��3@�wJ��!?�'��B��@����͐ٿ�@H|�@��B��3@�wJ��!?�'��B��@����͐ٿ�@H|�@��B��3@�wJ��!?�'��B��@�e���ٿ,�PJU�@p��^4@���Ѡ�!?*����д@�e���ٿ,�PJU�@p��^4@���Ѡ�!?*����д@�e���ٿ,�PJU�@p��^4@���Ѡ�!?*����д@�e���ٿ,�PJU�@p��^4@���Ѡ�!?*����д@��^*�ٿi�/���@*i�4@�>����!?�ʹ�%��@��^*�ٿi�/���@*i�4@�>����!?�ʹ�%��@��^*�ٿi�/���@*i�4@�>����!?�ʹ�%��@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@��7���ٿ-����@8�GA@�3@q��q��!?������@%�1���ٿ�7L�0��@�ّ�$�3@��I)�!?�(k�1�@%�1���ٿ�7L�0��@�ّ�$�3@��I)�!?�(k�1�@%�1���ٿ�7L�0��@�ّ�$�3@��I)�!?�(k�1�@%�1���ٿ�7L�0��@�ّ�$�3@��I)�!?�(k�1�@%�1���ٿ�7L�0��@�ّ�$�3@��I)�!?�(k�1�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@��1�ٿ�3��4f�@���s�3@
���,�!?�)2�#�@�C���ٿ+�����@���UP�3@�tn;�!?��&xw(�@�C���ٿ+�����@���UP�3@�tn;�!?��&xw(�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@I|_�O�ٿB�{��@�U����3@K��$ُ!?�o�8.�@���,u�ٿ����@�l����3@�/K��!?����O´@���,u�ٿ����@�l����3@�/K��!?����O´@53�ۗٿ���n�@[���9�3@��l4��!?�x[�z�@53�ۗٿ���n�@[���9�3@��l4��!?�x[�z�@53�ۗٿ���n�@[���9�3@��l4��!?�x[�z�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@�&	��ٿV�Q����@�����3@����!?>�O'=�@bt)�O�ٿ(+(�\~�@GT)<��3@-%W�!?�~�BZ�@bt)�O�ٿ(+(�\~�@GT)<��3@-%W�!?�~�BZ�@�*��K�ٿ�sz`)��@�<�+��3@ԇѩ��!?�� Bд@�*��K�ٿ�sz`)��@�<�+��3@ԇѩ��!?�� Bд@�.��ٿ%S*.r��@3d����3@"��!?�5 մ@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@��@!��ٿc��osj�@���3@�C+�!?��ݵ�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@W�-&�ٿg)�{�@�k/�1�3@mM�CB�!?*�R�O�@g�xZ�ٿ�{؂ ��@Xai���3@��>�,�!?:�/oɃ�@g�xZ�ٿ�{؂ ��@Xai���3@��>�,�!?:�/oɃ�@g�xZ�ٿ�{؂ ��@Xai���3@��>�,�!?:�/oɃ�@g�xZ�ٿ�{؂ ��@Xai���3@��>�,�!?:�/oɃ�@�r"�h�ٿ��Cj�@m68��3@�ߌ�+�!?X�+O �@�r"�h�ٿ��Cj�@m68��3@�ߌ�+�!?X�+O �@��h�ٿy3���@7���.�3@8�H�!?F�H�Ҡ�@��h�ٿy3���@7���.�3@8�H�!?F�H�Ҡ�@�+ւ'�ٿ�4f�c�@�	.���3@��O��!?t��w뮵@�O3~��ٿ��z�l��@�9"ş�3@�\9�!?ы���@�O3~��ٿ��z�l��@�9"ş�3@�\9�!?ы���@�O3~��ٿ��z�l��@�9"ş�3@�\9�!?ы���@V�
�<�ٿԅ6p��@A�ޤ,4@h�mBf�!?iՃ�O��@&��Ɛٿ��b��_�@S��8B�3@J9bX�!?��of��@�@�C�ٿ0H�KG�@���͎4@�؆L�!?H�iY	8�@�@�C�ٿ0H�KG�@���͎4@�؆L�!?H�iY	8�@�@�C�ٿ0H�KG�@���͎4@�؆L�!?H�iY	8�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@S^��ٿ'Ҥ}�@�%���3@>��6�!?AR�@���k�ٿ�h ^(�@���
��3@��(�!?bSm{̿�@���k�ٿ�h ^(�@���
��3@��(�!?bSm{̿�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@������ٿ �.���@R����4@����!?�pE�@:k'��ٿ�[�~о�@J���	�3@���q�!?���Z�W�@:k'��ٿ�[�~о�@J���	�3@���q�!?���Z�W�@��L.�ٿ�t��|�@=p'�4@��ȓ�!?��J�4x�@��L.�ٿ�t��|�@=p'�4@��ȓ�!?��J�4x�@��L.�ٿ�t��|�@=p'�4@��ȓ�!?��J�4x�@�r#��ٿE���@�@=��4@o���f�!?�|n�ݴ@�r#��ٿE���@�@=��4@o���f�!?�|n�ݴ@�r#��ٿE���@�@=��4@o���f�!?�|n�ݴ@�r#��ٿE���@�@=��4@o���f�!?�|n�ݴ@�r#��ٿE���@�@=��4@o���f�!?�|n�ݴ@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@	BXe�ٿ�N=�q�@%{޳��3@&-�K�!?!^�ϡ��@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@2��࡝ٿt?&��@����.�3@ q�:�!?ۅ3n3̴@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@���8 �ٿ�4���@b]]:��3@
^��O�!?�r�i�@��Ҙٿ�B�ӂ�@�C����3@�ǲ��!?^CN^J�@��Ҙٿ�B�ӂ�@�C����3@�ǲ��!?^CN^J�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��Ԅ��ٿix�x�@�5���3@⿬�3�!?�JX=̎�@��v^�ٿa����G�@��[t�3@��(�!?x���t{�@��v^�ٿa����G�@��[t�3@��(�!?x���t{�@��v^�ٿa����G�@��[t�3@��(�!?x���t{�@��v^�ٿa����G�@��[t�3@��(�!?x���t{�@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��D�b�ٿ�-����@�띵��3@ �P��!?	A
�5ĵ@��{)^�ٿ���nR��@�����3@ٯ����!?q}�эW�@��{)^�ٿ���nR��@�����3@ٯ����!?q}�эW�@����2�ٿ��lh�f�@���*�3@���XK�!?L�>Ya�@����2�ٿ��lh�f�@���*�3@���XK�!?L�>Ya�@����2�ٿ��lh�f�@���*�3@���XK�!?L�>Ya�@����2�ٿ��lh�f�@���*�3@���XK�!?L�>Ya�@]�w&��ٿ/8�/���@"q��3@��W��!?���6�@]�w&��ٿ/8�/���@"q��3@��W��!?���6�@]�w&��ٿ/8�/���@"q��3@��W��!?���6�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�9j�:�ٿTU���@�(
��3@�8���!?�_ߌ�D�@�d��ٿd�	�P�@��/@�3@f��ː!?Rj�=;�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@Y򎂮�ٿ5A܏���@��]�o�3@�:�#`�!?��;Q4�@F��6��ٿ�@���@��p�E�3@�=�!?)[�2Q��@F��6��ٿ�@���@��p�E�3@�=�!?)[�2Q��@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@;��w�ٿ�������@M �lX4@�0|�K�!?��5��S�@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�KfD��ٿ>��+��@�*L��4@M�!�m�!?��ܑ4��@�7�W �ٿ�.��K��@R�7ب�3@ے�,�!?�4񩣵�@�7�W �ٿ�.��K��@R�7ب�3@ے�,�!?�4񩣵�@�7�W �ٿ�.��K��@R�7ب�3@ے�,�!?�4񩣵�@�7�W �ٿ�.��K��@R�7ب�3@ے�,�!?�4񩣵�@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@nC~�ٿ�X"��Z�@����k�3@S�ߵE�!?c�#���@��;���ٿ
8���@��R�T�3@9 w�#�!?����@��;���ٿ
8���@��R�T�3@9 w�#�!?����@��;���ٿ
8���@��R�T�3@9 w�#�!?����@��;���ٿ
8���@��R�T�3@9 w�#�!?����@:j4���ٿC�$sT�@I6y�
�3@	�D�!?K�G�@5y�ٿ��c&���@�=���3@����2�!?-��T�@��b�J�ٿmS��і�@�I�o=�3@泉&u�!?�!'����@��b�J�ٿmS��і�@�I�o=�3@泉&u�!?�!'����@��b�J�ٿmS��і�@�I�o=�3@泉&u�!?�!'����@��b�J�ٿmS��і�@�I�o=�3@泉&u�!?�!'����@��b�J�ٿmS��і�@�I�o=�3@泉&u�!?�!'����@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@��D.��ٿ�yel"��@������3@&��b�!?Hd���7�@���ٿ�h����@~�Ǫ�4@�S}���!?0��5�@���ٿ�h����@~�Ǫ�4@�S}���!?0��5�@���ٿ�h����@~�Ǫ�4@�S}���!?0��5�@���w��ٿ�Y�� �@Y{j�Q�3@��|��!?}����;�@���w��ٿ�Y�� �@Y{j�Q�3@��|��!?}����;�@�V��Зٿ�HU'�@l�Q��3@pwb���!?�Z�=�@O�FӚٿ�0wU��@����S 4@b�q�`�!?�g�v��@�_�D��ٿ8j[�W�@9���4@����`�!?W�DuM�@�_�D��ٿ8j[�W�@9���4@����`�!?W�DuM�@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@.(Tc��ٿ�H�Ȗ��@Ji�<��3@�(�8��!?݆W��״@�f�v(�ٿ9qi�@�Z�Ų�3@��5N��!?VZX�Bݴ@�f�v(�ٿ9qi�@�Z�Ų�3@��5N��!?VZX�Bݴ@�f�v(�ٿ9qi�@�Z�Ų�3@��5N��!?VZX�Bݴ@�f�v(�ٿ9qi�@�Z�Ų�3@��5N��!?VZX�Bݴ@�f�v(�ٿ9qi�@�Z�Ų�3@��5N��!?VZX�Bݴ@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@}�N�2�ٿd<�^Ci�@)��J�3@�eY��!?'ν�x�@��7��ٿ�|
2_(�@j,��n�3@����!?Vd�H�@��7��ٿ�|
2_(�@j,��n�3@����!?Vd�H�@��zh��ٿ�\�Q��@��Ӛ��3@k�I�{�!?�c�D%�@��zh��ٿ�\�Q��@��Ӛ��3@k�I�{�!?�c�D%�@�K�x$�ٿ��T�e�@���=�3@˄#�Q�!?����@�@�=�8�ٿE��J
�@���� �3@'�x?8�!?	^׶F۵@�0h�}�ٿ��kJ2�@F[.�3@|�8+�!?,���!�@�0h�}�ٿ��kJ2�@F[.�3@|�8+�!?,���!�@�0h�}�ٿ��kJ2�@F[.�3@|�8+�!?,���!�@f��O�ٿ�aR��@ν���3@&wgN�!?�h�	6��@f��O�ٿ�aR��@ν���3@&wgN�!?�h�	6��@f��O�ٿ�aR��@ν���3@&wgN�!?�h�	6��@D����ٿr������@�� m��3@?��C�!?�2!�r��@�%����ٿ~�Z�բ�@:���3@ʦ�W%�!?��~bɴ@�%����ٿ~�Z�բ�@:���3@ʦ�W%�!?��~bɴ@©_'�ٿ�"��6v�@�Q�V �3@_�u�!?k�B2+8�@���ٿ��v�<�@�]��3@q)'�1�!?���!b�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@	'C�ٿe+ 
��@8����3@]�ea�!?٬/�@��睗ٿ���Pi��@�p����3@tٴ�Ώ!?�C�Ӵ@��睗ٿ���Pi��@�p����3@tٴ�Ώ!?�C�Ӵ@]���E�ٿ(J��D�@�cb�3@خ�濏!?��zW��@]���E�ٿ(J��D�@�cb�3@خ�濏!?��zW��@]���E�ٿ(J��D�@�cb�3@خ�濏!?��zW��@�Y�T�ٿ`�Ћ���@.�{4@��!?]�:��@�7���ٿY��武�@���3@�/w"L�!?�bYAյ@H��a��ٿ�אؿ��@�j_�3@Y_�3�!?�)o_�ѵ@H��a��ٿ�אؿ��@�j_�3@Y_�3�!?�)o_�ѵ@q9Be��ٿ�~����@���|��3@K-g"x�!?⴦���@q9Be��ٿ�~����@���|��3@K-g"x�!?⴦���@q9Be��ٿ�~����@���|��3@K-g"x�!?⴦���@G��^{�ٿ��|C\�@��Le�3@�V�M��!?�
�G�@G��^{�ٿ��|C\�@��Le�3@�V�M��!?�
�G�@G��^{�ٿ��|C\�@��Le�3@�V�M��!?�
�G�@G��^{�ٿ��|C\�@��Le�3@�V�M��!?�
�G�@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@�����ٿ�t��@(�s�f�3@\�.f�!?d6�7��@��N&�ٿ��am]M�@�X�H�3@�5�7��!?ل�V��@��N&�ٿ��am]M�@�X�H�3@�5�7��!?ل�V��@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@��r#4�ٿ�jֽ;�@�=��l�3@���~8�!?�ι�{R�@6 e83�ٿ-n|�?�@��Y��3@
�j�!?��馎�@6 e83�ٿ-n|�?�@��Y��3@
�j�!?��馎�@6 e83�ٿ-n|�?�@��Y��3@
�j�!?��馎�@ ی)��ٿ�YG��@��(4@����!?P��?޴@�Np�ٿ�7�_*w�@S�����3@�X��Ð!?�{_�d�@�Np�ٿ�7�_*w�@S�����3@�X��Ð!?�{_�d�@�Np�ٿ�7�_*w�@S�����3@�X��Ð!?�{_�d�@59����ٿ����@����3@�i5��!?�|�֙�@@��S̗ٿA�#�@���ܕ�3@�R�K�!?��_�|M�@@��S̗ٿA�#�@���ܕ�3@�R�K�!?��_�|M�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@~_���ٿD��qD�@U�T���3@y��c��!?oov^�	�@���ٿ�N{b](�@���u��3@�H�4�!? ��n�%�@���ٿ�N{b](�@���u��3@�H�4�!? ��n�%�@���ٿ�N{b](�@���u��3@�H�4�!? ��n�%�@���ٿ�N{b](�@���u��3@�H�4�!? ��n�%�@���ٿ�N{b](�@���u��3@�H�4�!? ��n�%�@d��MP�ٿM�����@�c���3@VP8�!??h�4)��@d��MP�ٿM�����@�c���3@VP8�!??h�4)��@d��MP�ٿM�����@�c���3@VP8�!??h�4)��@�69�ٿe��%3>�@i����3@*��Lo�!?�(s��D�@�69�ٿe��%3>�@i����3@*��Lo�!?�(s��D�@�8�6�ٿ���l׷�@T'�3@F�ӈ��!?`Bɿk^�@�8�6�ٿ���l׷�@T'�3@F�ӈ��!?`Bɿk^�@�8�6�ٿ���l׷�@T'�3@F�ӈ��!?`Bɿk^�@�8�6�ٿ���l׷�@T'�3@F�ӈ��!?`Bɿk^�@�8�6�ٿ���l׷�@T'�3@F�ӈ��!?`Bɿk^�@dz�O��ٿ�T�a0�@yf����3@�?�Ə!?d\��n�@dz�O��ٿ�T�a0�@yf����3@�?�Ə!?d\��n�@dz�O��ٿ�T�a0�@yf����3@�?�Ə!?d\��n�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�A�3N�ٿ 'h��@���U4@�8ޡ�!?DCW�w�@�q��p�ٿ~D��@o�@���V�3@d��-�!?֪���_�@�q��p�ٿ~D��@o�@���V�3@d��-�!?֪���_�@�q��p�ٿ~D��@o�@���V�3@d��-�!?֪���_�@斵׳�ٿ8T��L8�@4���_�3@�#�(��!?��Ħ��@斵׳�ٿ8T��L8�@4���_�3@�#�(��!?��Ħ��@斵׳�ٿ8T��L8�@4���_�3@�#�(��!?��Ħ��@斵׳�ٿ8T��L8�@4���_�3@�#�(��!?��Ħ��@斵׳�ٿ8T��L8�@4���_�3@�#�(��!?��Ħ��@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����ٿA��,C�@��B��3@�ޮ�!?���g�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@����i�ٿ)�Z1�@��q4@�N/�"�!?A.��y�@�;H��ٿ ����@;ZFe��3@o%QH.�!?o��Ma�@�;H��ٿ ����@;ZFe��3@o%QH.�!?o��Ma�@�;H��ٿ ����@;ZFe��3@o%QH.�!?o��Ma�@(�U�ٿ���KF@�@��']�3@:����!?փ��+ҵ@(�U�ٿ���KF@�@��']�3@:����!?փ��+ҵ@(�U�ٿ���KF@�@��']�3@:����!?փ��+ҵ@(�U�ٿ���KF@�@��']�3@:����!?փ��+ҵ@(�U�ٿ���KF@�@��']�3@:����!?փ��+ҵ@���g�ٿ��?�lz�@AӇ���3@JT�7��!?1�`��@�*��+�ٿ��y��@�LI�� 4@V<)V�!?�6�e�7�@�*��+�ٿ��y��@�LI�� 4@V<)V�!?�6�e�7�@�*��+�ٿ��y��@�LI�� 4@V<)V�!?�6�e�7�@Lɖ�M�ٿz`�K���@��B:�3@�����!?��Y�|�@��a��ٿ�(���@o�"�4@�r���!?��p��@��a��ٿ�(���@o�"�4@�r���!?��p��@��a��ٿ�(���@o�"�4@�r���!?��p��@��a��ٿ�(���@o�"�4@�r���!?��p��@ 05쁕ٿ�ɳd���@��_�R4@�?���!?�>�ƴ@ 05쁕ٿ�ɳd���@��_�R4@�?���!?�>�ƴ@ 05쁕ٿ�ɳd���@��_�R4@�?���!?�>�ƴ@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@u$Li��ٿ�?�3�@f�,\U4@K�C{��!?#�_*{��@��
_�ٿ�����@��8���3@�x�s�!?U��6��@��
_�ٿ�����@��8���3@�x�s�!?U��6��@��
_�ٿ�����@��8���3@�x�s�!?U��6��@��
_�ٿ�����@��8���3@�x�s�!?U��6��@��
_�ٿ�����@��8���3@�x�s�!?U��6��@mfD]��ٿC�����@�cқ��3@�K��j�!?�cyÁ�@mfD]��ٿC�����@�cқ��3@�K��j�!?�cyÁ�@mfD]��ٿC�����@�cқ��3@�K��j�!?�cyÁ�@mfD]��ٿC�����@�cқ��3@�K��j�!?�cyÁ�@mfD]��ٿC�����@�cқ��3@�K��j�!?�cyÁ�@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��TB<�ٿ�(�3Ծ�@[l�2��3@~���/�!?U�}�Aе@��`�ٿ�ѹ����@V��r=�3@r����!?ɓ_�L �@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���b�ٿ�5�.�2�@�S1�� 4@Lն4�!?���I��@���wf�ٿ�H9��n�@b�*Gx4@�j��!?O0�t�@
� w�ٿ�J#�4�@π���3@�Tj��!?d. i�@
� w�ٿ�J#�4�@π���3@�Tj��!?d. i�@
� w�ٿ�J#�4�@π���3@�Tj��!?d. i�@
� w�ٿ�J#�4�@π���3@�Tj��!?d. i�@
� w�ٿ�J#�4�@π���3@�Tj��!?d. i�@���Ďٿ��2�5��@�,�U
�3@�f	��!?u��1�q�@���Ďٿ��2�5��@�,�U
�3@�f	��!?u��1�q�@���Ďٿ��2�5��@�,�U
�3@�f	��!?u��1�q�@���Ďٿ��2�5��@�,�U
�3@�f	��!?u��1�q�@���Ďٿ��2�5��@�,�U
�3@�f	��!?u��1�q�@?db>�ٿt��s�b�@t��o�3@�O�_�!?� ����@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@�Aa�ٿsT`?:a�@e���R4@���<�!?c�@��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@������ٿ@���]�@��	Y��3@����!?�uфM��@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@VDP���ٿ�*�t�@��[�3@z�Is�!?L�{�;�@xٯ��ٿL���2��@�����3@~�]R�!?�;�&;�@�x�x�ٿvZQ�>�@��X���3@#bAd�!?�e���t�@�x�x�ٿvZQ�>�@��X���3@#bAd�!?�e���t�@�x�x�ٿvZQ�>�@��X���3@#bAd�!?�e���t�@�x�x�ٿvZQ�>�@��X���3@#bAd�!?�e���t�@bY*�N�ٿ�@���@�d��8�3@�B[@�!?�i=�$�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�[�1J�ٿ���C�@��3YB�3@��1B�!?�tM�1�@�A��ٿ��8)5��@E}�3@O>�ו�!?q��>�a�@�A��ٿ��8)5��@E}�3@O>�ו�!?q��>�a�@� s2�ٿ�)J+�@�.�?x4@���Đ!?!�F!e�@� s2�ٿ�)J+�@�.�?x4@���Đ!?!�F!e�@� s2�ٿ�)J+�@�.�?x4@���Đ!?!�F!e�@�K�zv�ٿ���@�߷d4@������!?�KK��@�K�zv�ٿ���@�߷d4@������!?�KK��@�K�zv�ٿ���@�߷d4@������!?�KK��@�K�zv�ٿ���@�߷d4@������!?�KK��@��X�ٿ�k�]���@���A�4@�#��!?��MF�6�@z	
�ŕٿ$�����@���Cf�3@���d�!?�Q�=��@z	
�ŕٿ$�����@���Cf�3@���d�!?�Q�=��@?��ӛٿX7�{��@甎_�4@^��e�!?J�ﳵ@?��ӛٿX7�{��@甎_�4@^��e�!?J�ﳵ@?��ӛٿX7�{��@甎_�4@^��e�!?J�ﳵ@?��ӛٿX7�{��@甎_�4@^��e�!?J�ﳵ@?��ӛٿX7�{��@甎_�4@^��e�!?J�ﳵ@���G��ٿq.��r��@̓)��4@���!?>pHРӴ@M�uD��ٿF��p4��@l?*w��3@СqH�!?�	�妴@M�uD��ٿF��p4��@l?*w��3@СqH�!?�	�妴@M�uD��ٿF��p4��@l?*w��3@СqH�!?�	�妴@M�uD��ٿF��p4��@l?*w��3@СqH�!?�	�妴@g�MQh�ٿ'm�m.I�@2�|�C4@㉒w(�!?�̔��y�@g�MQh�ٿ'm�m.I�@2�|�C4@㉒w(�!?�̔��y�@g�MQh�ٿ'm�m.I�@2�|�C4@㉒w(�!?�̔��y�@g�MQh�ٿ'm�m.I�@2�|�C4@㉒w(�!?�̔��y�@g�MQh�ٿ'm�m.I�@2�|�C4@㉒w(�!?�̔��y�@�N:B�ٿ�RWY��@Z��k 4@B�����!?�C���@�N:B�ٿ�RWY��@Z��k 4@B�����!?�C���@�N:B�ٿ�RWY��@Z��k 4@B�����!?�C���@�N:B�ٿ�RWY��@Z��k 4@B�����!?�C���@w�b��ٿ��+��@W�#h��3@�KL�!?�\\�⭴@w�b��ٿ��+��@W�#h��3@�KL�!?�\\�⭴@W)�{��ٿ��=� ��@���R��3@�&�碐!?Sy!~K��@�W�9�ٿH�wl�"�@VP�>��3@������!?a�Â0�@�W�9�ٿH�wl�"�@VP�>��3@������!?a�Â0�@�W�9�ٿH�wl�"�@VP�>��3@������!?a�Â0�@�W�9�ٿH�wl�"�@VP�>��3@������!?a�Â0�@�W�9�ٿH�wl�"�@VP�>��3@������!?a�Â0�@���պ�ٿ1��3I�@�|�B��3@�� \|�!?}�����@���պ�ٿ1��3I�@�|�B��3@�� \|�!?}�����@���պ�ٿ1��3I�@�|�B��3@�� \|�!?}�����@3�����ٿ���?G�@�Y�1`�3@�?��Z�!?��IzM�@3�����ٿ���?G�@�Y�1`�3@�?��Z�!?��IzM�@3�����ٿ���?G�@�Y�1`�3@�?��Z�!?��IzM�@3�����ٿ���?G�@�Y�1`�3@�?��Z�!?��IzM�@3�����ٿ���?G�@�Y�1`�3@�?��Z�!?��IzM�@��|��ٿ���)&��@c�*��3@�� ��!?�9�^bĵ@��|��ٿ���)&��@c�*��3@�� ��!?�9�^bĵ@���ٿ�I����@�I;�A�3@Ґ��!?Ez�<�Q�@���ٿ�I����@�I;�A�3@Ґ��!?Ez�<�Q�@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@��$ Ɵٿ�=�#���@�e�rA�3@5 �j�!?��n�O��@o�~�ٿ*�
����@�OW�3@\~k��!?�y����@�.^�ٿٌ��~��@�����3@_T`P�!?K�?���@�.^�ٿٌ��~��@�����3@_T`P�!?K�?���@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@�`$�p�ٿ�"tx�$�@��=���3@��M_�!?d�b
:��@����ٿb&��:��@�����3@�_F�?�!?d2m���@����ٿb&��:��@�����3@�_F�?�!?d2m���@����ٿb&��:��@�����3@�_F�?�!?d2m���@����ٿb&��:��@�����3@�_F�?�!?d2m���@����ٿb&��:��@�����3@�_F�?�!?d2m���@+�hE�ٿo�@՜�@ �`��3@:kO �!?����@+�hE�ٿo�@՜�@ �`��3@:kO �!?����@:��4�ٿ�؇��@'�5�3@��6W�!?{3���"�@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@?�Z�5�ٿ�o�5���@�cì��3@̟̄2�!?�K���@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@����؛ٿ�>�Ϣ�@��}n�3@��ʷ��!?�\���´@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@F`.�ʘٿK	�)�@C��b�3@�fYs�!?�j���@''*��ٿ�eL���@�����3@�u�S��!?n�~����@''*��ٿ�eL���@�����3@�u�S��!?n�~����@�=�R�ٿy�[n��@���8�3@	._ϻ�!?���s��@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@���7�ٿ����ܼ�@�����3@��z�A�!?%�o���@
��Y<�ٿǑt����@��_��3@iy���!?�jٴ?�@
��Y<�ٿǑt����@��_��3@iy���!?�jٴ?�@
��Y<�ٿǑt����@��_��3@iy���!?�jٴ?�@
��Y<�ٿǑt����@��_��3@iy���!?�jٴ?�@��u�l�ٿJ�EdB��@^��;��3@X���!?������@��u�l�ٿJ�EdB��@^��;��3@X���!?������@��u�l�ٿJ�EdB��@^��;��3@X���!?������@�m�ܕٿ^�i��
�@�k}6�3@n��c��!?Q�۷��@�m�ܕٿ^�i��
�@�k}6�3@n��c��!?Q�۷��@�m�ܕٿ^�i��
�@�k}6�3@n��c��!?Q�۷��@�m�ܕٿ^�i��
�@�k}6�3@n��c��!?Q�۷��@�<�,�ٿ:���s�@�a<��3@�:l4�!?�;=����@�M�ٿ�;k���@R���[�3@�l�Y�!?�2�&��@�M�ٿ�;k���@R���[�3@�l�Y�!?�2�&��@��FV��ٿ�6��!��@<p����3@�U��=�!?d��YV�@�Mgl�ٿ5��y�@��4@c�8�!?���1��@�Mgl�ٿ5��y�@��4@c�8�!?���1��@�Mgl�ٿ5��y�@��4@c�8�!?���1��@�Mgl�ٿ5��y�@��4@c�8�!?���1��@�!��ٿ��9�]��@�Q��4@_����!?���z�@�!��ٿ��9�]��@�Q��4@_����!?���z�@�!��ٿ��9�]��@�Q��4@_����!?���z�@�!��ٿ��9�]��@�Q��4@_����!?���z�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�F��ٿh�KI]N�@@I���3@n5(=�!?R�{�u�@�C�Q�ٿ&���A�@�k����3@�Ja瀐!?q]����@�C�Q�ٿ&���A�@�k����3@�Ja瀐!?q]����@�C�Q�ٿ&���A�@�k����3@�Ja瀐!?q]����@�C�Q�ٿ&���A�@�k����3@�Ja瀐!?q]����@�C�Q�ٿ&���A�@�k����3@�Ja瀐!?q]����@�Ej�ٿ4�����@��n��3@Ĭv�Ӑ!?(Y�Z��@����ٿ��>���@��p9��3@�O��!?и�4W�@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@	G�䋛ٿi9�-��@�'B�_�3@L�b	��!?��m�$��@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@���"�ٿkXZá�@�lg�3@����<�!?ލ�sNY�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@�xH��ٿs�pZ��@��m�x�3@�4p0?�!?��8D4�@cK���ٿ�܈���@�|��n�3@wӍ[�!?
�i��y�@cK���ٿ�܈���@�|��n�3@wӍ[�!?
�i��y�@X:x(��ٿtO�s��@ϴ.	 4@
cE�U�!?�1�Kw��@X:x(��ٿtO�s��@ϴ.	 4@
cE�U�!?�1�Kw��@X:x(��ٿtO�s��@ϴ.	 4@
cE�U�!?�1�Kw��@c��`�ٿ&���]��@F��3Z4@'bXy�!?M�W� �@c��`�ٿ&���]��@F��3Z4@'bXy�!?M�W� �@c��`�ٿ&���]��@F��3Z4@'bXy�!?M�W� �@c��`�ٿ&���]��@F��3Z4@'bXy�!?M�W� �@c��`�ٿ&���]��@F��3Z4@'bXy�!?M�W� �@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�p ��ٿ�Y�W-=�@��O���3@���O��!?,b����@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@�G���ٿ���A��@�ް�3@0��p�!?d�H@�j�@��2���ٿ=��3y��@�����3@����!?כ�(́�@��2���ٿ=��3y��@�����3@����!?כ�(́�@��2���ٿ=��3y��@�����3@����!?כ�(́�@��2���ٿ=��3y��@�����3@����!?כ�(́�@��2���ٿ=��3y��@�����3@����!?כ�(́�@���`8�ٿo[�$��@�;D���3@��W"�!?�%=[��@���`8�ٿo[�$��@�;D���3@��W"�!?�%=[��@���`8�ٿo[�$��@�;D���3@��W"�!?�%=[��@���`8�ٿo[�$��@�;D���3@��W"�!?�%=[��@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@Ƒ�I�ٿ�!*����@'���W�3@RC�a�!?�=c���@�����ٿ��xu;�@�>�h��3@��p]�!?~+mA�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@�>Y��ٿ��Ҵ�-�@M���3@��=Hb�!?-�ҳ~�@T�V�+�ٿ�=���[�@��ë�3@XE�<�!? �ߜc�@T�V�+�ٿ�=���[�@��ë�3@XE�<�!? �ߜc�@T�V�+�ٿ�=���[�@��ë�3@XE�<�!? �ߜc�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@?bB,��ٿM�C�V�@l5Y�4@� 
1l�!?mȅ�U�@���}s�ٿe���y��@*+�4@%���p�!?���
g�@���}s�ٿe���y��@*+�4@%���p�!?���
g�@���}s�ٿe���y��@*+�4@%���p�!?���
g�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@�%�ۖٿ<ٻ�%�@(�7	��3@����p�!?�J?��b�@��6�ޏٿ��㧳��@��3� 4@��'�C�!?=^l}�V�@i�!�ٿ@Z�A�@'ll�3@��}�V�!?�S�|�@i�!�ٿ@Z�A�@'ll�3@��}�V�!?�S�|�@i�!�ٿ@Z�A�@'ll�3@��}�V�!?�S�|�@i�!�ٿ@Z�A�@'ll�3@��}�V�!?�S�|�@i�!�ٿ@Z�A�@'ll�3@��}�V�!?�S�|�@�BW֍ٿN֡=�<�@�����3@K�u���!?h6R���@!��M��ٿ�XF��!�@m�I�	�3@]5�ԏ!?H�6\[�@!��M��ٿ�XF��!�@m�I�	�3@]5�ԏ!?H�6\[�@]�-�4�ٿ��&�j�@l�"���3@PcT��!?"�Z����@]�-�4�ٿ��&�j�@l�"���3@PcT��!?"�Z����@]�-�4�ٿ��&�j�@l�"���3@PcT��!?"�Z����@^��V��ٿd@/�Lf�@O�0��3@ǚ�h�!?��(:#=�@^��V��ٿd@/�Lf�@O�0��3@ǚ�h�!?��(:#=�@�h��i�ٿz<�*�@i�#��3@!6�No�!?L�^U��@�h��i�ٿz<�*�@i�#��3@!6�No�!?L�^U��@W#\9��ٿ�N�:¬�@��/9�3@�\���!?���h�@W#\9��ٿ�N�:¬�@��/9�3@�\���!?���h�@W#\9��ٿ�N�:¬�@��/9�3@�\���!?���h�@W#\9��ٿ�N�:¬�@��/9�3@�\���!?���h�@W#\9��ٿ�N�:¬�@��/9�3@�\���!?���h�@o���ٿ%��u-��@�����3@����!?�y5��)�@�h�9�ٿ~��OF��@��_0�3@/ �� �!?�V���@�h�9�ٿ~��OF��@��_0�3@/ �� �!?�V���@�h�9�ٿ~��OF��@��_0�3@/ �� �!?�V���@�h�9�ٿ~��OF��@��_0�3@/ �� �!?�V���@�h�9�ٿ~��OF��@��_0�3@/ �� �!?�V���@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@d��Eܗٿ��/ >�@kP'�	�3@��J!�!?�8�mѫ�@�f��z�ٿ��*io��@�o�K�3@�u�e�!?�7~$�:�@�f��z�ٿ��*io��@�o�K�3@�u�e�!?�7~$�:�@�f��z�ٿ��*io��@�o�K�3@�u�e�!?�7~$�:�@�f��z�ٿ��*io��@�o�K�3@�u�e�!?�7~$�:�@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@*�/���ٿXQ��c�@��Ą>�3@"��_�!?Ő�3��@K �5�ٿ�����@�@}��!�3@����=�!?|>K�⦵@K �5�ٿ�����@�@}��!�3@����=�!?|>K�⦵@K �5�ٿ�����@�@}��!�3@����=�!?|>K�⦵@K �5�ٿ�����@�@}��!�3@����=�!?|>K�⦵@�܌��ٿ��c����@�"�`�3@nm�f�!?���Lu�@�܌��ٿ��c����@�"�`�3@nm�f�!?���Lu�@˥>�ٿ��g���@e���4@�G[��!?�De�a�@˥>�ٿ��g���@e���4@�G[��!?�De�a�@˥>�ٿ��g���@e���4@�G[��!?�De�a�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@M�H��ٿ�4~$�d�@Z��f��3@�j�g�!?=��Wzk�@���m��ٿ,�1��K�@�3�ϋ�3@����[�!?����|#�@�Jb��ٿ��@���@���u;�3@����U�!?���ܴ@�Jb��ٿ��@���@���u;�3@����U�!?���ܴ@�Jb��ٿ��@���@���u;�3@����U�!?���ܴ@�Jb��ٿ��@���@���u;�3@����U�!?���ܴ@�Jb��ٿ��@���@���u;�3@����U�!?���ܴ@܅
��ٿ��!� 5�@�����3@u�|k��!?�V��@܅
��ٿ��!� 5�@�����3@u�|k��!?�V��@܅
��ٿ��!� 5�@�����3@u�|k��!?�V��@܅
��ٿ��!� 5�@�����3@u�|k��!?�V��@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@9�WH1�ٿ2�da�u�@��\f��3@K�l�_�!?H#.�b�@yZVO��ٿ�u�3}�@�
�`�4@�����!?���ڵZ�@yZVO��ٿ�u�3}�@�
�`�4@�����!?���ڵZ�@�jLU�ٿ.M�{��@�|���3@܃���!?�QIA�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@\뿰�ٿ4�5��*�@�Yn�m�3@h�A��!?l�0�m�@��@�ٿi[& m�@'��D�3@�N��w�!?z8b��$�@��@�ٿi[& m�@'��D�3@�N��w�!?z8b��$�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@�,�>:�ٿ=p�l%�@��J��3@��c?�!?|��RI�@;��d=�ٿ9V"3�@߻���3@	3.{�!?jI_d[�@;��d=�ٿ9V"3�@߻���3@	3.{�!?jI_d[�@;��d=�ٿ9V"3�@߻���3@	3.{�!?jI_d[�@;��d=�ٿ9V"3�@߻���3@	3.{�!?jI_d[�@�8�X͏ٿ}ܑ2z��@Lk;]4@�&:�!?����ݒ�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@�G��ٿ������@ߺO=4@	�+�&�!?&ry��#�@����ٿ�-@|�T�@1rօ�3@@��I�!?��h	o��@����ٿ�-@|�T�@1rօ�3@@��I�!?��h	o��@~�g�ٿz4�l�@Su�
��3@�kmI�!?��*la��@ ��m3�ٿ{5so��@<*��y�3@��)i_�!?y閟"��@ ��m3�ٿ{5so��@<*��y�3@��)i_�!?y閟"��@ ��m3�ٿ{5so��@<*��y�3@��)i_�!?y閟"��@ ��m3�ٿ{5so��@<*��y�3@��)i_�!?y閟"��@�k�dݖٿ�UwxD�@n,|f�3@: P�h�!?r~w�Q�@�k�dݖٿ�UwxD�@n,|f�3@: P�h�!?r~w�Q�@�k�dݖٿ�UwxD�@n,|f�3@: P�h�!?r~w�Q�@���伏ٿz� R2��@�:-y��3@��2L�!?���Cj��@���伏ٿz� R2��@�:-y��3@��2L�!?���Cj��@��3D��ٿgf��#i�@����3@F$ 7�!?0���@��3D��ٿgf��#i�@����3@F$ 7�!?0���@��3D��ٿgf��#i�@����3@F$ 7�!?0���@̮��ٿ�d1Ȍ�@���4@����!?G�[��@̮��ٿ�d1Ȍ�@���4@����!?G�[��@̮��ٿ�d1Ȍ�@���4@����!?G�[��@̮��ٿ�d1Ȍ�@���4@����!?G�[��@̮��ٿ�d1Ȍ�@���4@����!?G�[��@b�)q��ٿ�mA��@Y&�[��3@�gky�!?�%�bv�@b�)q��ٿ�mA��@Y&�[��3@�gky�!?�%�bv�@��W;�ٿu��M���@��; ��3@�e��!?w�F���@��W;�ٿu��M���@��; ��3@�e��!?w�F���@AZ���ٿ���RY[�@teO���3@8־1�!?��k�l�@�Zta��ٿv6H���@�F��W�3@;����!?�v�m�A�@�Zta��ٿv6H���@�F��W�3@;����!?�v�m�A�@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@�@E�i�ٿ�t���S�@dYGJ��3@�S�Ð!?���t��@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@��6'�ٿɣi�CF�@M�0��3@��ΐ!?��+ę�@����ٿ�����@u�'���3@Y����!?���˵@����ٿ�����@u�'���3@Y����!?���˵@����ٿ�����@u�'���3@Y����!?���˵@����ٿ�����@u�'���3@Y����!?���˵@�4�(�ٿχ�����@5��B��3@�m>��!?���싵@-
[���ٿ��(`��@ƝPQ�3@>;�oǐ!?:�;Iv��@k�gu�ٿI���v��@�.��x�3@���N8�!?O���@k�gu�ٿI���v��@�.��x�3@���N8�!?O���@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@R�PA)�ٿ)������@�Rn��3@,�y�"�!?I5cل�@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��*�ٿ~�`ۿp�@��p;�3@���#�!?�3�[���@��Р�ٿ cѿO��@%7j��3@��!qF�!?q�}X[�@��Р�ٿ cѿO��@%7j��3@��!qF�!?q�}X[�@��Р�ٿ cѿO��@%7j��3@��!qF�!?q�}X[�@��Р�ٿ cѿO��@%7j��3@��!qF�!?q�}X[�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@B)�>˖ٿ/m����@��4@�[��?�!?����-O�@�1M8Кٿ���r��@�Z���3@�y�?�!?FG�^Ѵ@�;*���ٿ���P��@��]�8�3@�YE�!?��7 ���@�;*���ٿ���P��@��]�8�3@�YE�!?��7 ���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@VȨ�ٿ���{��@�¨�44@[���;�!? ��|���@_��%��ٿ�h�&���@���# 4@o���!?����@@hO��ٿ�)����@��D���3@�#����!?|i˭���@@hO��ٿ�)����@��D���3@�#����!?|i˭���@@hO��ٿ�)����@��D���3@�#����!?|i˭���@@hO��ٿ�)����@��D���3@�#����!?|i˭���@@hO��ٿ�)����@��D���3@�#����!?|i˭���@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@G�M���ٿ�Hf�Q�@ �R��3@д�-a�!?B(;�ݴ@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@+?>Ŗٿ��\���@o<��i�3@��g�\�!?�.�[��@��Ji+�ٿ�1�����@�&��z�3@��O �!?�F
��"�@��Ji+�ٿ�1�����@�&��z�3@��O �!?�F
��"�@��l��ٿB���2�@ixM�� 4@���B�!?e���o�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@��ǝٿ�����H�@���:��3@���W�!?3��ܕF�@G��a�ٿ�mI��d�@�8.���3@�tEa�!?+�sT��@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@�|%�ٿ�Ņ�ؑ�@E����3@�T ��!?�9���/�@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@b8涛ٿ�n�#� �@���t��3@�1v�!�!?n
R-��@Ɋ��)�ٿ{D�a���@*4��.�3@�Ҁ��!?�%��*�@Ɋ��)�ٿ{D�a���@*4��.�3@�Ҁ��!?�%��*�@Ɋ��)�ٿ{D�a���@*4��.�3@�Ҁ��!?�%��*�@������ٿ�̪|���@�o׎��3@S�x,�!?�(�/_�@	Qv��ٿ�g����@�"��3@��:w�!?ށ���$�@	Qv��ٿ�g����@�"��3@��:w�!?ށ���$�@	Qv��ٿ�g����@�"��3@��:w�!?ށ���$�@	Qv��ٿ�g����@�"��3@��:w�!?ށ���$�@,^!��ٿZ��/zY�@Ӌo���3@b?�㑐!?�(誴@,^!��ٿZ��/zY�@Ӌo���3@b?�㑐!?�(誴@,^!��ٿZ��/zY�@Ӌo���3@b?�㑐!?�(誴@ȕ��_�ٿP�} ��@����3@�F���!?�JX�Ԓ�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@[�s �ٿ��#9�@���"��3@"\Ga�!?d�n8�@�X3Ğٿ��:��)�@�h�G�3@��sm�!?_4�m��@�X3Ğٿ��:��)�@�h�G�3@��sm�!?_4�m��@�X3Ğٿ��:��)�@�h�G�3@��sm�!?_4�m��@�X3Ğٿ��:��)�@�h�G�3@��sm�!?_4�m��@�X3Ğٿ��:��)�@�h�G�3@��sm�!?_4�m��@6�� t�ٿDV����@��5R�3@������!?	/�|���@Z�1�ٿ�Q�2���@�e��o�3@����\�!?�����ִ@	vm�2�ٿ�q�)���@����f�3@^����!?C(�C)D�@	vm�2�ٿ�q�)���@����f�3@^����!?C(�C)D�@E���ُٿ�-��I��@P�z��3@�p��!?�iR���@�����ٿ���4:H�@K1��3@ԥ�:�!?�bhZ�@�����ٿ���4:H�@K1��3@ԥ�:�!?�bhZ�@�����ٿ���4:H�@K1��3@ԥ�:�!?�bhZ�@�����ٿ���4:H�@K1��3@ԥ�:�!?�bhZ�@�F��e�ٿq��	���@���}3�3@��]a�!?.����@�F��e�ٿq��	���@���}3�3@��]a�!?.����@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�?i��ٿ������@wC�/�3@���67�!?�t�
1�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�oN�ٿ�dS.^3�@���3@@Q��'�!?InZ#5b�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@�6yR�ٿ~$�Q�@k�&��3@��X�!?�U�_!�@��Pb�ٿ88;����@��D��3@��8��!?g�6�@��Pb�ٿ88;����@��D��3@��8��!?g�6�@��Pb�ٿ88;����@��D��3@��8��!?g�6�@��Pb�ٿ88;����@��D��3@��8��!?g�6�@��Pb�ٿ88;����@��D��3@��8��!?g�6�@U�J���ٿhy�]N�@>�8��3@�Xӏ��!?ч̧/�@U�J���ٿhy�]N�@>�8��3@�Xӏ��!?ч̧/�@U�J���ٿhy�]N�@>�8��3@�Xӏ��!?ч̧/�@U�J���ٿhy�]N�@>�8��3@�Xӏ��!?ч̧/�@�ȴ��ٿ- ��bJ�@z��ͯ�3@�~�e��!?�*�	^�@�ȴ��ٿ- ��bJ�@z��ͯ�3@�~�e��!?�*�	^�@�/�Z�ٿy�YQ0N�@%��m�3@�c�Z@�!?0!�;�ϴ@�/�Z�ٿy�YQ0N�@%��m�3@�c�Z@�!?0!�;�ϴ@�/�Z�ٿy�YQ0N�@%��m�3@�c�Z@�!?0!�;�ϴ@0(b5��ٿ�v�o�@,�[˽�3@���I�!?��8�ش@0h����ٿ����C�@��Z��3@�Iþf�!?�}:)�@��h��ٿ�6T�I��@�'��v�3@���[��!?}��y�P�@%��ѕٿ�rH.���@����3@�gN�V�!??GP�(�@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@iR�ٿ�9�����@�yP�\�3@�6��!?k��=�ʹ@�#���ٿ�^|Z4��@�x+�4@��B
.�!?ˢ%/\��@�#���ٿ�^|Z4��@�x+�4@��B
.�!?ˢ%/\��@�#���ٿ�^|Z4��@�x+�4@��B
.�!?ˢ%/\��@�R��˓ٿ�l�`��@���V�3@j{|�!?c�G�_��@�R��˓ٿ�l�`��@���V�3@j{|�!?c�G�_��@:�0�{�ٿH��;6�@~�����3@Z1�B��!?8�8�	��@:�0�{�ٿH��;6�@~�����3@Z1�B��!?8�8�	��@:�0�{�ٿH��;6�@~�����3@Z1�B��!?8�8�	��@:�0�{�ٿH��;6�@~�����3@Z1�B��!?8�8�	��@:�0�{�ٿH��;6�@~�����3@Z1�B��!?8�8�	��@^׭���ٿ�c%����@2��j�3@�L��N�!?x�oC4۴@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@Fފ�|�ٿ�N�`�H�@��xZ�3@	_���!?:s����@�Փ���ٿ3&��R��@�}
��3@�U��4�!?������@�Փ���ٿ3&��R��@�}
��3@�U��4�!?������@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@#�o}1�ٿ����F�@'����3@�d�;��!?�}�`�ȴ@g���ٿ������@@�@�m�3@\�|B�!?�޿���@g���ٿ������@@�@�m�3@\�|B�!?�޿���@g���ٿ������@@�@�m�3@\�|B�!?�޿���@g���ٿ������@@�@�m�3@\�|B�!?�޿���@g���ٿ������@@�@�m�3@\�|B�!?�޿���@g���ٿ������@@�@�m�3@\�|B�!?�޿���@y�tϚٿ�ML�.�@k���V�3@e%�Ve�!?�`��@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@J��ٿ�eP���@mhL��3@��Eq�!?�,Ӕ�@m��e�ٿ{�"0�@���=Y�3@���t�!?2�
ɴ@m��e�ٿ{�"0�@���=Y�3@���t�!?2�
ɴ@m��e�ٿ{�"0�@���=Y�3@���t�!?2�
ɴ@�����ٿ�w(�"�@�	K͓�3@��jy�!?	�����@�����ٿ�w(�"�@�	K͓�3@��jy�!?	�����@�����ٿ�w(�"�@�	K͓�3@��jy�!?	�����@�����ٿ�w(�"�@�	K͓�3@��jy�!?	�����@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@�$�ol�ٿm��K��@��x���3@S/����!?�98H�W�@_�㓸�ٿWY����@uTâ��3@�|zHT�!?����Hv�@_�㓸�ٿWY����@uTâ��3@�|zHT�!?����Hv�@_�㓸�ٿWY����@uTâ��3@�|zHT�!?����Hv�@_�㓸�ٿWY����@uTâ��3@�|zHT�!?����Hv�@_�㓸�ٿWY����@uTâ��3@�|zHT�!?����Hv�@�X��ٿ//y��@f�ѣ�3@D���=�!?�� Ѻ�@�X��ٿ//y��@f�ѣ�3@D���=�!?�� Ѻ�@]���S�ٿn�K���@4.I��3@��/��!?�:���ʹ@]���S�ٿn�K���@4.I��3@��/��!?�:���ʹ@]���S�ٿn�K���@4.I��3@��/��!?�:���ʹ@]���S�ٿn�K���@4.I��3@��/��!?�:���ʹ@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@�!ۤ=�ٿ׭`����@��19<�3@��9~/�!?)d�;Q�@i�V��ٿ(�s�$}�@�}I�3@��^��!?�<�,ƴ@i�V��ٿ(�s�$}�@�}I�3@��^��!?�<�,ƴ@i�V��ٿ(�s�$}�@�}I�3@��^��!?�<�,ƴ@�>�;�ٿUܝTS�@׏_���3@�&�?�!?�C����@s��綒ٿ.b�����@��^�3@��d��!?2굀��@s��綒ٿ.b�����@��^�3@��d��!?2굀��@s��綒ٿ.b�����@��^�3@��d��!?2굀��@s��綒ٿ.b�����@��^�3@��d��!?2굀��@Q61c�ٿ�?���@�5��3@;V����!?.�FS1�@Q61c�ٿ�?���@�5��3@;V����!?.�FS1�@Q61c�ٿ�?���@�5��3@;V����!?.�FS1�@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@���O(�ٿm�!V��@l6y���3@;+�!?�h����@j��՘ٿ�vb���@3aX���3@_�=��!?�:9��s�@j��՘ٿ�vb���@3aX���3@_�=��!?�:9��s�@j��՘ٿ�vb���@3aX���3@_�=��!?�:9��s�@j��՘ٿ�vb���@3aX���3@_�=��!?�:9��s�@czO��ٿ�H-�Q�@N ��M�3@6��"��!?V���tS�@czO��ٿ�H-�Q�@N ��M�3@6��"��!?V���tS�@���X�ٿ�OO���@g]��/4@���r��!?�?`1!*�@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@<�4��ٿ�\0!��@w�Gm�3@H�N�!?�鈘��@�^�q�ٿN��0���@=���+�3@�ڛ9�!?A��\���@?WFkw�ٿ���h:�@\6�̷�3@�:#R<�!?�r�3��@��L�ߙٿe|ѯ�n�@�����3@0���!?{$���Q�@�d�ތ�ٿ���p2��@�N,b��3@hg�ga�!?�-yM�´@�d�ތ�ٿ���p2��@�N,b��3@hg�ga�!?�-yM�´@����ٿ�U4ry�@�I/��3@=Ԃ|)�!?� b���@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@ԯ��ٿ�u6�`��@+��3@Ē>m�!?�[�l��@�7˖�ٿB�E � �@c+�h�3@K|+9�!?�wl ��@�7˖�ٿB�E � �@c+�h�3@K|+9�!?�wl ��@�7˖�ٿB�E � �@c+�h�3@K|+9�!?�wl ��@�%Ɠ
�ٿ-���2v�@K�"�+�3@Hs�!?H�x�E��@�%Ɠ
�ٿ-���2v�@K�"�+�3@Hs�!?H�x�E��@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���)��ٿ�_]�q�@٪>��3@�ih8�!?\w�BV�@���M�ٿK�J��Q�@��kq�4@`��U4�!?緘n$�@���M�ٿK�J��Q�@��kq�4@`��U4�!?緘n$�@5_pM��ٿ�9�]&�@������3@譥�j�!?5K�ИN�@5_pM��ٿ�9�]&�@������3@譥�j�!?5K�ИN�@5_pM��ٿ�9�]&�@������3@譥�j�!?5K�ИN�@��?��ٿo4$X)��@����3@� �`��!?B��;.�@��[ʛٿ؅�-X��@�f��l�3@�;�O�!?B5̃�B�@��[ʛٿ؅�-X��@�f��l�3@�;�O�!?B5̃�B�@�m
0�ٿ��3 ���@8���3@��:{�!?��5`�@�m
0�ٿ��3 ���@8���3@��:{�!?��5`�@�m
0�ٿ��3 ���@8���3@��:{�!?��5`�@�m
0�ٿ��3 ���@8���3@��:{�!?��5`�@����ٿS�����@E;w(�3@�Z.�!?��.T��@����ٿS�����@E;w(�3@�Z.�!?��.T��@����ٿS�����@E;w(�3@�Z.�!?��.T��@����ٿS�����@E;w(�3@�Z.�!?��.T��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@�2��ٿ��~�ś�@���3@&/�BL�!?2�Q�o��@k��ٿ)��*�z�@�e��3@���Rx�!?;��ZL\�@k��ٿ)��*�z�@�e��3@���Rx�!?;��ZL\�@�q�ٿ���CC��@�}S�P�3@��~���!?	�&$]��@�q�ٿ���CC��@�}S�P�3@��~���!?	�&$]��@�q�ٿ���CC��@�}S�P�3@��~���!?	�&$]��@�q�ٿ���CC��@�}S�P�3@��~���!?	�&$]��@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@/�p�ٿ'�[a�@�tT�4@\�Ɣ6�!?FZ�.�@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@�g_9��ٿ�������@��2��3@=����!?!�����@SB��%�ٿ�;9*2t�@��2 4@Cp�RN�!?���$���@BL�0�ٿ��p]p�@&^-9��3@�}V�!?��H(��@BL�0�ٿ��p]p�@&^-9��3@�}V�!?��H(��@�	��l�ٿ�{' N�@i��Q��3@��cb�!?�019r�@�	��l�ٿ�{' N�@i��Q��3@��cb�!?�019r�@����ȍٿ�8.�E��@�?��5�3@W����!?8j�0G�@��ݎٿ2��20�@���Ff�3@A2���!?x��1��@��ݎٿ2��20�@���Ff�3@A2���!?x��1��@��ݎٿ2��20�@���Ff�3@A2���!?x��1��@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��<h��ٿS&B���@�nn%�4@K�p�S�!?P#n֍�@��rE>�ٿ��+��@�k��3@(	Q�@�!?sZ��70�@��rE>�ٿ��+��@�k��3@(	Q�@�!?sZ��70�@��rE>�ٿ��+��@�k��3@(	Q�@�!?sZ��70�@pč�g�ٿW�N2�w�@��3���3@�EP$�!?n��~���@��،��ٿ�����@�k�3@P�g�!?J���er�@��،��ٿ�����@�k�3@P�g�!?J���er�@��،��ٿ�����@�k�3@P�g�!?J���er�@��،��ٿ�����@�k�3@P�g�!?J���er�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@�:p��ٿDz�R�@�4䙒�3@k�-0?�!?��F�@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@3���ٿ�u��[�@�\�;'�3@1����!?T�H5&��@��u��ٿ�(��0��@��;�3@��\�!?E4�6��@��u��ٿ�(��0��@��;�3@��\�!?E4�6��@DK'e��ٿ��-���@#��3@�)V0�!?4b��л�@DK'e��ٿ��-���@#��3@�)V0�!?4b��л�@DK'e��ٿ��-���@#��3@�)V0�!?4b��л�@DK'e��ٿ��-���@#��3@�)V0�!?4b��л�@DK'e��ٿ��-���@#��3@�)V0�!?4b��л�@�����ٿڶ9��п@f*!v��3@{
� �!?64��0�@�����ٿڶ9��п@f*!v��3@{
� �!?64��0�@�����ٿڶ9��п@f*!v��3@{
� �!?64��0�@�����ٿڶ9��п@f*!v��3@{
� �!?64��0�@�]�'��ٿ?x` �}�@���|�3@���R��!?���u�@�]�'��ٿ?x` �}�@���|�3@���R��!?���u�@�e!�ٿD��|��@��U�3@F��|ӏ!?�SQ�Dٵ@�e!�ٿD��|��@��U�3@F��|ӏ!?�SQ�Dٵ@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@�NOe>�ٿ�u�]�@�H~A4@��uC�!?s���a�@���ᇚٿ�A�i���@�[�R�3@+���}�!?�)�OY�@���<�ٿĝoS��@�^c�3@���K�!?�)0Z��@���<�ٿĝoS��@�^c�3@���K�!?�)0Z��@ԮTH�ٿ�ͤF��@�ُM�3@l#1�!?�ʻ�d��@ԮTH�ٿ�ͤF��@�ُM�3@l#1�!?�ʻ�d��@X�0�O�ٿd�(��@�"@��3@\'W�W�!?R�m.�ܴ@X�0�O�ٿd�(��@�"@��3@\'W�W�!?R�m.�ܴ@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@R:\��ٿF�CV�?�@U�Q�3@3��9�!?��~���@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@N:yi�ٿr� ���@G�@��3@/�H�f�!?�LE��Ӵ@,�Љ�ٿ������@R��
��3@�F�q�!?&W�8�@,�Љ�ٿ������@R��
��3@�F�q�!?&W�8�@,�Љ�ٿ������@R��
��3@�F�q�!?&W�8�@,�Љ�ٿ������@R��
��3@�F�q�!?&W�8�@�8�ѯ�ٿ��U�w�@���W�3@�S�%~�!?�&E���@�8�ѯ�ٿ��U�w�@���W�3@�S�%~�!?�&E���@�8�ѯ�ٿ��U�w�@���W�3@�S�%~�!?�&E���@�8�ѯ�ٿ��U�w�@���W�3@�S�%~�!?�&E���@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@N�*�`�ٿG���`��@�SQa�3@;�S1�!?�E&)?�@',�W��ٿkR\#]��@ ��[�3@���0��!?Y+��к�@Z6��Ȕٿ	i���C�@��h��3@��=�b�!?~��|}��@�h�ّٿ���@V��@P��^�3@�[��W�!?�N�g�@�h�ّٿ���@V��@P��^�3@�[��W�!?�N�g�@�h�ّٿ���@V��@P��^�3@�[��W�!?�N�g�@�h�ّٿ���@V��@P��^�3@�[��W�!?�N�g�@�h�ّٿ���@V��@P��^�3@�[��W�!?�N�g�@�FU�Бٿ����E�@������3@#�O}��!?d�����@�z�s�ٿMn!��@�z�#44@z��׎�!?8��]X�@�z�s�ٿMn!��@�z�#44@z��׎�!?8��]X�@�z�s�ٿMn!��@�z�#44@z��׎�!?8��]X�@��ܫy�ٿ����ȯ�@�T�0�3@F��v�!?&�B1�@��ܫy�ٿ����ȯ�@�T�0�3@F��v�!?&�B1�@��ܫy�ٿ����ȯ�@�T�0�3@F��v�!?&�B1�@��ܫy�ٿ����ȯ�@�T�0�3@F��v�!?&�B1�@��ܫy�ٿ����ȯ�@�T�0�3@F��v�!?&�B1�@G�KYՑٿ'N\֑��@�a���3@�;��M�!?��F�t�@G�KYՑٿ'N\֑��@�a���3@�;��M�!?��F�t�@G�KYՑٿ'N\֑��@�a���3@�;��M�!?��F�t�@�Y��ٿ�E����@��gY��3@�XDB�!?UIE4xt�@�8RY�ٿ�l��@�=ɉ4@�h��?�!?M���ĵ@�8RY�ٿ�l��@�=ɉ4@�h��?�!?M���ĵ@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@g*�~��ٿI�,}���@��^�3@�ha��!?���M׮�@������ٿ{WF����@7�Ƅ��3@�ڇ��!?���&��@�ne�ٿ�����@3���3@�k=m�!?���e7��@�ne�ٿ�����@3���3@�k=m�!?���e7��@�ne�ٿ�����@3���3@�k=m�!?���e7��@�ne�ٿ�����@3���3@�k=m�!?���e7��@�ne�ٿ�����@3���3@�k=m�!?���e7��@�u����ٿ<����{�@���)��3@��-ߐ!?z��/]�@�;N�ٿ��b���@����3@�~��l�!?C0���@�;N�ٿ��b���@����3@�~��l�!?C0���@�;N�ٿ��b���@����3@�~��l�!?C0���@�uj)�ٿV-k�?�@�up��4@��i�z�!?�i�<޴@�uj)�ٿV-k�?�@�up��4@��i�z�!?�i�<޴@�uj)�ٿV-k�?�@�up��4@��i�z�!?�i�<޴@�����ٿ婖3���@����4@�|R�!?�b�=(�@�x�7m�ٿ1�K�:�@���4@S\a��!?�������@�x�7m�ٿ1�K�:�@���4@S\a��!?�������@`nL�#�ٿ8�3�/�@R����3@M���!?�iQд@`nL�#�ٿ8�3�/�@R����3@M���!?�iQд@�h��`�ٿ�*�d�@�j�=��3@Օ�ڏ!?�����#�@�h��`�ٿ�*�d�@�j�=��3@Օ�ڏ!?�����#�@�h��`�ٿ�*�d�@�j�=��3@Օ�ڏ!?�����#�@�h��`�ٿ�*�d�@�j�=��3@Օ�ڏ!?�����#�@�g�s_�ٿ�(T%�@�P����3@::z�Տ!?a�\Cz�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@5R�p��ٿ�[��@$��$9�3@?�x�!?�Ńp�>�@�n�Q�ٿ�R$&:�@�.L�3@u2W>A�!?�H��p�@�n�Q�ٿ�R$&:�@�.L�3@u2W>A�!?�H��p�@�n�Q�ٿ�R$&:�@�.L�3@u2W>A�!?�H��p�@��R		�ٿ�J�1K�@mL�G�3@��p�!?'�t»´@��R		�ٿ�J�1K�@mL�G�3@��p�!?'�t»´@��R		�ٿ�J�1K�@mL�G�3@��p�!?'�t»´@��R		�ٿ�J�1K�@mL�G�3@��p�!?'�t»´@��R		�ٿ�J�1K�@mL�G�3@��p�!?'�t»´@��sH�ٿ�n����@M��e��3@S���!?��K��ŵ@��sH�ٿ�n����@M��e��3@S���!?��K��ŵ@��sH�ٿ�n����@M��e��3@S���!?��K��ŵ@��sH�ٿ�n����@M��e��3@S���!?��K��ŵ@��C��ٿ��p�D�@y��>�3@�M��!?�����@��C��ٿ��p�D�@y��>�3@�M��!?�����@��C��ٿ��p�D�@y��>�3@�M��!?�����@=�}3��ٿ�����@N���4@�(�aG�!?=Ww$�@=�}3��ٿ�����@N���4@�(�aG�!?=Ww$�@��Δ�ٿgWX?�@9-����3@���Pu�!?/B�_F�@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@1Q�Մ�ٿ�Zu|��@��BLR�3@{���!?*��õ@�|	QőٿN�����@G�px�3@���5�!?^3BW,�@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�?�/�ٿi��ǥ��@�(���3@EE�($�!?J�:��@�yڣ��ٿ��q����@wS@���3@�N}��!?׈g�\ŵ@�yڣ��ٿ��q����@wS@���3@�N}��!?׈g�\ŵ@�yڣ��ٿ��q����@wS@���3@�N}��!?׈g�\ŵ@�yڣ��ٿ��q����@wS@���3@�N}��!?׈g�\ŵ@�yڣ��ٿ��q����@wS@���3@�N}��!?׈g�\ŵ@�����ٿd��t�X�@ϴ%�.�3@Z=�;�!?�f��-�@�����ٿd��t�X�@ϴ%�.�3@Z=�;�!?�f��-�@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@<�E��ٿ���6���@�؃m��3@l[.Ny�!?���δ@DG�ٿE�CM��@$�$���3@����Ð!? ����N�@DG�ٿE�CM��@$�$���3@����Ð!? ����N�@DG�ٿE�CM��@$�$���3@����Ð!? ����N�@DG�ٿE�CM��@$�$���3@����Ð!? ����N�@rb�V<�ٿ������@\i��4@��׈�!?.����4�@��rE��ٿ�9׃��@���,4@玈��!?
�7��@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@��@�w�ٿm3�M�)�@�t�T�4@Бf6��!?���|���@V����ٿ�t� �0�@٥����3@�Bd�!?>�)α�@j�ٿ������@�_QG�3@��&�<�!?����v�@j�ٿ������@�_QG�3@��&�<�!?����v�@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@���牓ٿ��O��@�T�3@�X��L�!?���Y �@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@	�6�Ǎٿ�V���@zΙH�4@����Y�!?r������@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�7�ٿT�ZFxK�@��Ob�4@$i�G�!?�����u�@�BW3�ٿ�(8E��@P2h<4@w��~�!?���U!��@�BW3�ٿ�(8E��@P2h<4@w��~�!?���U!��@�BW3�ٿ�(8E��@P2h<4@w��~�!?���U!��@�BW3�ٿ�(8E��@P2h<4@w��~�!?���U!��@�BW3�ٿ�(8E��@P2h<4@w��~�!?���U!��@9ې ��ٿ4���X�@��v4@����!?���/�@���ی�ٿ>0l��Y�@Og\/� 4@�<�8M�!?C�{ݴ@$�v���ٿ�2��"�@���E�3@�f�v�!?�<BO�@$�v���ٿ�2��"�@���E�3@�f�v�!?�<BO�@�x	�ٿ�2�nX�@h�?ۦ4@ᥡ�u�!?����B�@�x	�ٿ�2�nX�@h�?ۦ4@ᥡ�u�!?����B�@�x	�ٿ�2�nX�@h�?ۦ4@ᥡ�u�!?����B�@lgE�ؒٿZ-�G5[�@���4@��֤.�!?�O^�@��N/=�ٿh���@�V��u4@�L55�!?{K��ִ@��N/=�ٿh���@�V��u4@�L55�!?{K��ִ@��N/=�ٿh���@�V��u4@�L55�!?{K��ִ@��N/=�ٿh���@�V��u4@�L55�!?{K��ִ@��N/=�ٿh���@�V��u4@�L55�!?{K��ִ@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@�L��^�ٿ�m�ߞb�@��k_4@ߎf�b�!?a�t���@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@*Vu�\�ٿ��*��@�P��l�3@qe�=�!?����T�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@[eHHE�ٿ�V<mM�@�?A��3@_K|w�!?�q�k�@uq6�ٿ=�h��@P�E�x�3@�>��Ə!?��e%s^�@,�T�ٿ����|�@9D�,�4@Y��J�!?O,ԼPT�@,�T�ٿ����|�@9D�,�4@Y��J�!?O,ԼPT�@�>�`5�ٿ2�%���@@�Y���3@�âw��!?-����@�>�`5�ٿ2�%���@@�Y���3@�âw��!?-����@�>�`5�ٿ2�%���@@�Y���3@�âw��!?-����@�>�`5�ٿ2�%���@@�Y���3@�âw��!?-����@�f�<k�ٿIz�vE�@=|@�4�3@�����!?�cJAB�@���}��ٿ!�� �X�@O�.8��3@�?sr�!?/^�I��@���}��ٿ!�� �X�@O�.8��3@�?sr�!?/^�I��@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@�QX��ٿ��U�1�@4\���3@:���!?���mv�@x�Heؙٿ��D|T��@$�A�T�3@�OU�!?�VS ?�@x�Heؙٿ��D|T��@$�A�T�3@�OU�!?�VS ?�@x�Heؙٿ��D|T��@$�A�T�3@�OU�!?�VS ?�@��/)ǛٿdQ�L]��@}��0��3@�ncb��!?��g|��@�u�XG�ٿZ1s�b�@&=����3@K�W�}�!?�ߪk�@�u�XG�ٿZ1s�b�@&=����3@K�W�}�!?�ߪk�@����ٿ��+r�\�@4VZ}�4@�P���!?�5���@����ٿ��+r�\�@4VZ}�4@�P���!?�5���@����_�ٿ��&8`�@Yg�U�4@u�"𢡄!?@��8vӴ@����_�ٿ��&8`�@Yg�U�4@u�"𢡄!?@��8vӴ@����_�ٿ��&8`�@Yg�U�4@u�"𢡄!?@��8vӴ@�]iOR�ٿR2x�\�@ٯ� 4@�D��!?P����5�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@4W�>K�ٿ����f�@�l�1
4@��cp�!?���!�@p�OC�ٿ{g�:@ �@���6� 4@�z\�C�!?��U1�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@�����ٿ#��U��@��-
4@ 7��M�!?�5*�Zg�@���/3�ٿ�d,��@=PE��4@4[��x�!?	�b䀵@���/3�ٿ�d,��@=PE��4@4[��x�!?	�b䀵@���/3�ٿ�d,��@=PE��4@4[��x�!?	�b䀵@���/3�ٿ�d,��@=PE��4@4[��x�!?	�b䀵@�ǔٿwRS���@O��3@�����!?��n�~�@s�(��ٿ�����@ �N��3@�!S�#�!?|s$�E�@s�(��ٿ�����@ �N��3@�!S�#�!?|s$�E�@s�(��ٿ�����@ �N��3@�!S�#�!?|s$�E�@s�(��ٿ�����@ �N��3@�!S�#�!?|s$�E�@���3��ٿ4OU�Hp�@{X�p�3@s�I�!?���Ĵ@���3��ٿ4OU�Hp�@{X�p�3@s�I�!?���Ĵ@���3��ٿ4OU�Hp�@{X�p�3@s�I�!?���Ĵ@���3��ٿ4OU�Hp�@{X�p�3@s�I�!?���Ĵ@��曙�ٿ~��A0�@��D�3@��f�!?Ձ�����@��曙�ٿ~��A0�@��D�3@��f�!?Ձ�����@��曙�ٿ~��A0�@��D�3@��f�!?Ձ�����@��曙�ٿ~��A0�@��D�3@��f�!?Ձ�����@o+���ٿ�!�4�C�@�����3@ꌨԻ�!?LUaB��@o+���ٿ�!�4�C�@�����3@ꌨԻ�!?LUaB��@o+���ٿ�!�4�C�@�����3@ꌨԻ�!?LUaB��@o+���ٿ�!�4�C�@�����3@ꌨԻ�!?LUaB��@�+E��ٿ��R\��@a��ȼ4@���$�!?>��F�.�@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@TF6�ٿZיγ�@�O���3@���_�!?��!���@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@D��[Ҕٿ�b�(q^�@+_��R�3@a�]Y�!?���،�@�!ޘٿ���M��@�C����3@���D4�!?6&��Or�@�!ޘٿ���M��@�C����3@���D4�!?6&��Or�@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@�zw��ٿiq����@.�e��3@�̾W��!?>�D���@5�Bⵙٿ�h~L��@�ߘ��3@t�Uv�!?�ي��v�@5�Bⵙٿ�h~L��@�ߘ��3@t�Uv�!?�ي��v�@5�Bⵙٿ�h~L��@�ߘ��3@t�Uv�!?�ي��v�@5�Bⵙٿ�h~L��@�ߘ��3@t�Uv�!?�ي��v�@5�Bⵙٿ�h~L��@�ߘ��3@t�Uv�!?�ي��v�@��궉�ٿ��ыV+�@�f ���3@r{	.R�!?������@��궉�ٿ��ыV+�@�f ���3@r{	.R�!?������@�J���ٿ_o�Je�@p9��q�3@�EThC�!?����ӵ@QM��V�ٿ���pW�@��z��3@��M�%�!?�����L�@QM��V�ٿ���pW�@��z��3@��M�%�!?�����L�@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@�tH��ٿ�E�t�|�@�w�h�3@ީs�^�!?t'}:)ϴ@IM�f��ٿ��[1$�@w�����3@����!?�nPh��@IM�f��ٿ��[1$�@w�����3@����!?�nPh��@IM�f��ٿ��[1$�@w�����3@����!?�nPh��@,��	[�ٿ�X(m�R�@��o/}�3@l��$�!?���(�@,��	[�ٿ�X(m�R�@��o/}�3@l��$�!?���(�@?K{?_�ٿ���_���@L]���3@�"���!?:�m���@?K{?_�ٿ���_���@L]���3@�"���!?:�m���@�H3ݗٿ�e��b�@wU�3@0K�#�!?�oS�#�@�T��̗ٿމ�����@��4�3@l=z��!?��$bf�@�T��̗ٿމ�����@��4�3@l=z��!?��$bf�@�T��̗ٿމ�����@��4�3@l=z��!?��$bf�@�T��̗ٿމ�����@��4�3@l=z��!?��$bf�@�T��̗ٿމ�����@��4�3@l=z��!?��$bf�@E���;�ٿL\	"�@�=���3@�NFCؐ!?�Clд@��r�;�ٿp������@��u��4@0Y�Α�!?���Up�@��r�;�ٿp������@��u��4@0Y�Α�!?���Up�@��r�;�ٿp������@��u��4@0Y�Α�!?���Up�@��r�;�ٿp������@��u��4@0Y�Α�!?���Up�@X8jT�ٿ0�}���@ ��3�3@7ӂߞ�!?�ٗ�0�@X8jT�ٿ0�}���@ ��3�3@7ӂߞ�!?�ٗ�0�@X8jT�ٿ0�}���@ ��3�3@7ӂߞ�!?�ٗ�0�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@��8��ٿ��0�;�@Z�����3@�5u=,�!?l�,�
~�@%p�ڳ�ٿL��2�@{�C���3@��#i�!?�Q���@%p�ڳ�ٿL��2�@{�C���3@��#i�!?�Q���@%p�ڳ�ٿL��2�@{�C���3@��#i�!?�Q���@�oRڐٿ)k�@�We��3@��w�!?��s��@�oRڐٿ)k�@�We��3@��w�!?��s��@�O�ۣ�ٿk���S�@�^E�3@wC�hΐ!?���:��@�y6�h�ٿ̟}HI��@2o@Z�3@�\ө�!?
�C����@�y6�h�ٿ̟}HI��@2o@Z�3@�\ө�!?
�C����@�y6�h�ٿ̟}HI��@2o@Z�3@�\ө�!?
�C����@�y6�h�ٿ̟}HI��@2o@Z�3@�\ө�!?
�C����@�IH�q�ٿ��D�U�@���_�3@^6����!?�E�9�ɴ@�IH�q�ٿ��D�U�@���_�3@^6����!?�E�9�ɴ@.�3y�ٿFbb]��@r˂��3@Z����!?�z��p�@.�3y�ٿFbb]��@r˂��3@Z����!?�z��p�@�+�Ɏ�ٿ��׸���@ͅb���3@���=�!?)M88��@�+�Ɏ�ٿ��׸���@ͅb���3@���=�!?)M88��@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@M��̚ٿ�y2���@F"�V��3@1�6�2�!?2��p�]�@�aOE��ٿ�㑛{�@�6�г�3@��<�8�!?E���(�@�aOE��ٿ�㑛{�@�6�г�3@��<�8�!?E���(�@�aOE��ٿ�㑛{�@�6�г�3@��<�8�!?E���(�@�aOE��ٿ�㑛{�@�6�г�3@��<�8�!?E���(�@�aOE��ٿ�㑛{�@�6�г�3@��<�8�!?E���(�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@nJޚ �ٿ2]����@��E��4@�=���!?�T��\�@�~[/��ٿ�i](u��@R�H?��3@F!�!?��Zb�@�~[/��ٿ�i](u��@R�H?��3@F!�!?��Zb�@�~[/��ٿ�i](u��@R�H?��3@F!�!?��Zb�@�~[/��ٿ�i](u��@R�H?��3@F!�!?��Zb�@�~[/��ٿ�i](u��@R�H?��3@F!�!?��Zb�@GY��ٿ����@�fP���3@.��Ə!?R�# <X�@GY��ٿ����@�fP���3@.��Ə!?R�# <X�@�k�4��ٿY�j��@p\߫x�3@0�@�!?�$�	��@�k�4��ٿY�j��@p\߫x�3@0�@�!?�$�	��@�����ٿ�h�<J�@�����3@��dDK�!?o�O�@�����ٿ�h�<J�@�����3@��dDK�!?o�O�@�����ٿ�h�<J�@�����3@��dDK�!?o�O�@�����ٿ�h�<J�@�����3@��dDK�!?o�O�@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@��'���ٿS�{�0��@�I���3@�V��!?�$�/д@B��r�ٿ�17���@il=��3@�A��V�!?ʋB���@B��r�ٿ�17���@il=��3@�A��V�!?ʋB���@ Yk�"�ٿM�%��@d���?�3@t�}�_�!?�~�|!�@ Yk�"�ٿM�%��@d���?�3@t�}�_�!?�~�|!�@ Yk�"�ٿM�%��@d���?�3@t�}�_�!?�~�|!�@y�#��ٿ�Z�l,��@�U`��3@��q�!?�4�_�ߴ@y�#��ٿ�Z�l,��@�U`��3@��q�!?�4�_�ߴ@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@����D�ٿa2�Ȍ��@�6U-q�3@ynZ�V�!?ѳgB���@0��H�ٿ҉W�q��@ϫz	�3@P��f�!?�l�g��@0��H�ٿ҉W�q��@ϫz	�3@P��f�!?�l�g��@}I֑�ٿ�L��@P�j�l�3@_��K��!?�]©�մ@}I֑�ٿ�L��@P�j�l�3@_��K��!?�]©�մ@}I֑�ٿ�L��@P�j�l�3@_��K��!?�]©�մ@}I֑�ٿ�L��@P�j�l�3@_��K��!?�]©�մ@}I֑�ٿ�L��@P�j�l�3@_��K��!?�]©�մ@�g�Y�ٿ�A��@�\�v��3@I�K�A�!??�����@�g�Y�ٿ�A��@�\�v��3@I�K�A�!??�����@�g�Y�ٿ�A��@�\�v��3@I�K�A�!??�����@�g�Y�ٿ�A��@�\�v��3@I�K�A�!??�����@�g�Y�ٿ�A��@�\�v��3@I�K�A�!??�����@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�d���ٿ��ß�>�@��P�3@V�2�'�!?�,���@�].���ٿT���3�@���a��3@Av_�!?l=�g*ٵ@�0��ٿ�B{�U�@o���R�3@�m/N�!?��U�6�@�0��ٿ�B{�U�@o���R�3@�m/N�!?��U�6�@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@>��u�ٿ�k����@7�5n4@�qJl��!?R骅��@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��~�ٿ���a���@��]��3@*.;���!?�u��T�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@��a'�ٿ��گ�@��[U�3@]¥b�!?��N;�@_3:?�ٿ�(?��@�!D��3@"`e�!?�X��@_3:?�ٿ�(?��@�!D��3@"`e�!?�X��@_3:?�ٿ�(?��@�!D��3@"`e�!?�X��@_3:?�ٿ�(?��@�!D��3@"`e�!?�X��@Ă�-�ٿ�T��c�@��ěi�3@geكf�!?_z�o�@Ă�-�ٿ�T��c�@��ěi�3@geكf�!?_z�o�@Ă�-�ٿ�T��c�@��ěi�3@geكf�!?_z�o�@���p��ٿ��>ď�@3
�޽4@�<��!?�q���@���p��ٿ��>ď�@3
�޽4@�<��!?�q���@���p��ٿ��>ď�@3
�޽4@�<��!?�q���@���p��ٿ��>ď�@3
�޽4@�<��!?�q���@�'��ٿ����;�@��!{>�3@��X晐!?8/�sg�@�'��ٿ����;�@��!{>�3@��X晐!?8/�sg�@�'��ٿ����;�@��!{>�3@��X晐!?8/�sg�@�}�w�ٿ��i����@���3@��e!��!?Z�2z�۵@�}�w�ٿ��i����@���3@��e!��!?Z�2z�۵@�}�w�ٿ��i����@���3@��e!��!?Z�2z�۵@�}�w�ٿ��i����@���3@��e!��!?Z�2z�۵@�F<���ٿe<tc�>�@��K��3@�b6-�!?;�UP](�@�F<���ٿe<tc�>�@��K��3@�b6-�!?;�UP](�@�F<���ٿe<tc�>�@��K��3@�b6-�!?;�UP](�@�F<���ٿe<tc�>�@��K��3@�b6-�!?;�UP](�@�F<���ٿe<tc�>�@��K��3@�b6-�!?;�UP](�@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@��ղ��ٿ0�=}���@ʍ���3@�"����!?.�mJ��@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@������ٿ1&p�>^�@q��9��3@�-����!?g=�c�@��A,��ٿ^2re�@l�����3@m�͒�!?��/r�@4㛦g�ٿXW�q�@�f^���3@P5'�6�!?~�M���@�Bš�ٿQ�G8��@a�Mj��3@0.�X+�!?&����@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@f��S�ٿ���!�@��m@3�3@K!�!?�.��L;�@"�u��ٿ�b�� 2�@�$���3@!�[KF�!?�h �!�@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@aSUU��ٿ`��{���@ �(�F�3@��h�V�!?�zCrC��@�hp��ٿz��Du��@���f|�3@ͭ'�u�!?���3Kg�@�hp��ٿz��Du��@���f|�3@ͭ'�u�!?���3Kg�@]���ٿ]F�r�z�@i`,���3@�wG�!?EƋ�fB�@]���ٿ]F�r�z�@i`,���3@�wG�!?EƋ�fB�@��WW�ٿ͈����@��]���3@�U���!?H�Y��@��WW�ٿ͈����@��]���3@�U���!?H�Y��@��WW�ٿ͈����@��]���3@�U���!?H�Y��@��WW�ٿ͈����@��]���3@�U���!?H�Y��@��WW�ٿ͈����@��]���3@�U���!?H�Y��@^٭�k�ٿ���!�@�T����3@K���!?tq?ad�@^٭�k�ٿ���!�@�T����3@K���!?tq?ad�@^٭�k�ٿ���!�@�T����3@K���!?tq?ad�@^٭�k�ٿ���!�@�T����3@K���!?tq?ad�@�s�{�ٿ!��[��@>^�SF�3@�>�#�!?
��ɹ��@�s�{�ٿ!��[��@>^�SF�3@�>�#�!?
��ɹ��@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@������ٿ(��"o�@F����3@� �!? ]����@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@���ٿ��q����@>\?���3@�#�n+�!?�"��G�@����ٿ~̃(|��@�:mv�3@�x��!�!?]_4S���@����ٿ~̃(|��@�:mv�3@�x��!�!?]_4S���@����ٿ~̃(|��@�:mv�3@�x��!�!?]_4S���@����ٿ~̃(|��@�:mv�3@�x��!�!?]_4S���@�g�[��ٿ�[sן�@b�f 4@�?��!?���@�*��ٿ���z�@��&Ô4@�Q�T�!?�/*�P�@�*��ٿ���z�@��&Ô4@�Q�T�!?�/*�P�@��p��ٿ�5�=(�@���Q�3@Ǹ:Z^�!?Ml�Վ�@k1�.�ٿ�ZJp��@� ����3@S�5)�!?T���´@k1�.�ٿ�ZJp��@� ����3@S�5)�!?T���´@k1�.�ٿ�ZJp��@� ����3@S�5)�!?T���´@k1�.�ٿ�ZJp��@� ����3@S�5)�!?T���´@k1�.�ٿ�ZJp��@� ����3@S�5)�!?T���´@*��;��ٿY��}��@������3@6	�U3�!?�v���h�@�O��ٿ�-l=���@�;���3@QH,���!?�q����@�O��ٿ�-l=���@�;���3@QH,���!?�q����@�O��ٿ�-l=���@�;���3@QH,���!?�q����@�O��ٿ�-l=���@�;���3@QH,���!?�q����@�O��ٿ�-l=���@�;���3@QH,���!?�q����@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@+���ٿ�,��Ɵ�@�/�^�4@������!?7n=n�T�@��P���ٿ�T4v���@_KO�4�3@쑑4��!?9@���|�@��P���ٿ�T4v���@_KO�4�3@쑑4��!?9@���|�@��P���ٿ�T4v���@_KO�4�3@쑑4��!?9@���|�@��~�ӌٿ򦹳��@"G�A7�3@�N����!?�2ߴ�{�@	�=p�ٿC�����@���E�4@P��)/�!?�E��ޅ�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@�Ğ�ٿ|S��@���Y��3@����!?ȉ�,�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@ki�ܮ�ٿ�ꇞ���@#��ٛ�3@C�D�?�!?@�7��k�@�O�ٿ�)U�@n�,���3@�ӄ�Z�!?�%F�V�@�O�ٿ�)U�@n�,���3@�ӄ�Z�!?�%F�V�@^�L�5�ٿ4H�6���@�\�j��3@��d'Z�!?&~��7��@^�L�5�ٿ4H�6���@�\�j��3@��d'Z�!?&~��7��@^�L�5�ٿ4H�6���@�\�j��3@��d'Z�!?&~��7��@5�o�9�ٿy{!�I�@��� +�3@~��8�!?�����@5�o�9�ٿy{!�I�@��� +�3@~��8�!?�����@5�o�9�ٿy{!�I�@��� +�3@~��8�!?�����@5�o�9�ٿy{!�I�@��� +�3@~��8�!?�����@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@'ħr9�ٿ�23R��@�\J�3@�йx1�!?�N�D�B�@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@���mx�ٿ ����@��~B^�3@��q�P�!?�ps .��@����|�ٿ����@24|�3@ DӤ)�!?v`0�
�@����|�ٿ����@24|�3@ DӤ)�!?v`0�
�@����|�ٿ����@24|�3@ DӤ)�!?v`0�
�@����|�ٿ����@24|�3@ DӤ)�!?v`0�
�@����|�ٿ����@24|�3@ DӤ)�!?v`0�
�@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@���%M�ٿz�c��\�@Qc�^�3@�o�%1�!?�2����@{
��ٿԸ[� �@�ā�a�3@y���-�!?9ͭ2�@X�r���ٿ�i�m��@P ��Q�3@C�{zx�!?����@5�@X�r���ٿ�i�m��@P ��Q�3@C�{zx�!?����@5�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@�6آ�ٿy�TG�@ƶ���3@v0�W�!?��@��M�@
��p4�ٿ�مS���@���@d�3@��l�!?%h��^�@
��p4�ٿ�مS���@���@d�3@��l�!?%h��^�@��r�%�ٿ^T����@�C7�3@��P�0�!?���`)V�@��r�%�ٿ^T����@�C7�3@��P�0�!?���`)V�@��YÎٿ�����b�@aI���3@pT,�q�!?�ު�*�@��YÎٿ�����b�@aI���3@pT,�q�!?�ު�*�@��YÎٿ�����b�@aI���3@pT,�q�!?�ު�*�@��YÎٿ�����b�@aI���3@pT,�q�!?�ު�*�@�=�p�ٿ?���oq�@oR��3@ێ��<�!?���J�C�@�=�p�ٿ?���oq�@oR��3@ێ��<�!?���J�C�@�=�p�ٿ?���oq�@oR��3@ێ��<�!?���J�C�@�=�p�ٿ?���oq�@oR��3@ێ��<�!?���J�C�@�=�p�ٿ?���oq�@oR��3@ێ��<�!?���J�C�@�x�f�ٿ���)6��@C�z�3@	�_�W�!?�%ܴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@Y1�ʁ�ٿq��[X�@r��f0�3@�fo-ҏ!?a��+�ɴ@{�e�ٿ����c
�@}B�]4@#C?}��!?���W�0�@ni蜙ٿ����@�(��G�3@o�<I��!?�A|�@ni蜙ٿ����@�(��G�3@o�<I��!?�A|�@ni蜙ٿ����@�(��G�3@o�<I��!?�A|�@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@=���d�ٿ+�/v��@�v/���3@���na�!?�R6��@���B��ٿ�D>��@�v�
��3@76�؄�!?�1R(/U�@���B��ٿ�D>��@�v�
��3@76�؄�!?�1R(/U�@���B��ٿ�D>��@�v�
��3@76�؄�!?�1R(/U�@���B��ٿ�D>��@�v�
��3@76�؄�!?�1R(/U�@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@6XW��ٿ��9psz�@�@�L�3@�R��c�!?� (���@���2Ƙٿc�e��@�V�8��3@�1��!?I���@�+�J8�ٿE)Bv7q�@N�:�i�3@�<�B�!?�Y�>u�@�+�J8�ٿE)Bv7q�@N�:�i�3@�<�B�!?�Y�>u�@�+�J8�ٿE)Bv7q�@N�:�i�3@�<�B�!?�Y�>u�@�+�J8�ٿE)Bv7q�@N�:�i�3@�<�B�!?�Y�>u�@�+�J8�ٿE)Bv7q�@N�:�i�3@�<�B�!?�Y�>u�@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@�jE�[�ٿsw4�r��@�U��3@?&KM>�!?���G��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@���T�ٿ#�l\�K�@\N�Nz�3@.��3b�!?M	�#��@�/���ٿak�L���@~�p�3@�GL�S�!?�xZ�l�@����ٿ��bb�o�@��vj�3@�"���!?��z�@�cf��ٿ��L����@*�u�3@�o��!?�#�n�@�cf��ٿ��L����@*�u�3@�o��!?�#�n�@0{9A�ٿn�
��@f�`�3@ �fi��!?�Z�����@8#1"��ٿ$@�|�@H>V�K�3@�c��!?�Б$�@8#1"��ٿ$@�|�@H>V�K�3@�c��!?�Б$�@8#1"��ٿ$@�|�@H>V�K�3@�c��!?�Б$�@ڻ��n�ٿi� �\��@P�ԩu�3@n�T�U�!?g�Kj�@ڻ��n�ٿi� �\��@P�ԩu�3@n�T�U�!?g�Kj�@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@���I�ٿ�)�j��@@'׃��3@v�ҳ�!?-��WJ��@��a��ٿ9��ZH6�@������3@�Ǖ�!?��k�ҵ@d���ٿ�J=I��@1)	�a�3@Ac9�!?����ĵ@d���ٿ�J=I��@1)	�a�3@Ac9�!?����ĵ@d���ٿ�J=I��@1)	�a�3@Ac9�!?����ĵ@�B~�ٿ˝�)�@���ht�3@K�5�F�!?/2��@�@�B~�ٿ˝�)�@���ht�3@K�5�F�!?/2��@�@�ey�/�ٿ�������@�Q��W�3@c�G�~�!?؋���@�ey�/�ٿ�������@�Q��W�3@c�G�~�!?؋���@H,Q�ٿaH P��@�W���3@L��5{�!?d���b�@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@a����ٿ�v�a~.�@��Sj��3@l�;w��!?LJ[&+��@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@"(�֛ٿ��� ��@�O����3@���')�!?������@�Q�ږٿ�lT�b�@��;���3@0n�De�!?˾��ة�@�Q�ږٿ�lT�b�@��;���3@0n�De�!?˾��ة�@�Q�ږٿ�lT�b�@��;���3@0n�De�!?˾��ة�@�Q�ږٿ�lT�b�@��;���3@0n�De�!?˾��ة�@��[�ٿ����@^�3�� 4@�R��8�!?��jb�Z�@��[�ٿ����@^�3�� 4@�R��8�!?��jb�Z�@��[�ٿ����@^�3�� 4@�R��8�!?��jb�Z�@��[�ٿ����@^�3�� 4@�R��8�!?��jb�Z�@��[�ٿ����@^�3�� 4@�R��8�!?��jb�Z�@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@;>�W��ٿ�����@�Z�4@����?�!?�)���@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@�ԯ�ٿ�@�Y�@�-sm�3@��E�8�!?�ȏU��@���pF�ٿ��ы��@;FO@�3@W��H�!?`קN��@���pF�ٿ��ы��@;FO@�3@W��H�!?`קN��@���pF�ٿ��ы��@;FO@�3@W��H�!?`קN��@9Ez�9�ٿq��\8��@�u�\3�3@�2�r�!?Y�^<x�@¬,�9�ٿ`�&�Ɨ�@"?,��3@5��:�!?�.�담@o��x�ٿJ8y����@Ho_��3@��;&�!?c��寯�@�:��ٓٿ-��JO�@���MP�3@� w倐!?���h��@�:��ٓٿ-��JO�@���MP�3@� w倐!?���h��@E�	�v�ٿɜDM<$�@� ����3@+RRJ��!?=6��@=�J@P�ٿ$��0�T�@9�7���3@p��k�!?���>���@=�J@P�ٿ$��0�T�@9�7���3@p��k�!?���>���@=�J@P�ٿ$��0�T�@9�7���3@p��k�!?���>���@=�J@P�ٿ$��0�T�@9�7���3@p��k�!?���>���@�ݿ���ٿ�>ʗ��@�b�̵ 4@1@iO<�!?�Q+��2�@�ݿ���ٿ�>ʗ��@�b�̵ 4@1@iO<�!?�Q+��2�@e��UƑٿ=x�#�W�@}�g�P�3@�Dj(p�!?ڳ�D�@0�🝐ٿ�;:��?�@�n�lQ�3@s��)�!?v5�/8�@0�🝐ٿ�;:��?�@�n�lQ�3@s��)�!?v5�/8�@0�🝐ٿ�;:��?�@�n�lQ�3@s��)�!?v5�/8�@D����ٿ��A�%t�@?1��q�3@��Bm^�!?s�N�@D����ٿ��A�%t�@?1��q�3@��Bm^�!?s�N�@D����ٿ��A�%t�@?1��q�3@��Bm^�!?s�N�@[�<�܊ٿ�o����@Q�pd�3@;�)�F�!?\�[fI��@[�<�܊ٿ�o����@Q�pd�3@;�)�F�!?\�[fI��@[�<�܊ٿ�o����@Q�pd�3@;�)�F�!?\�[fI��@[�<�܊ٿ�o����@Q�pd�3@;�)�F�!?\�[fI��@����l�ٿ_�xL�.�@�!5�3@��ȍ1�!?��Ԕ�S�@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@#��l�ٿl��1dj�@��6_K�3@6��i�!?�5a���@����ٿ�|Ro�@�����3@{8,�!?_�u|��@����ٿ�|Ro�@�����3@{8,�!?_�u|��@����ٿ�|Ro�@�����3@{8,�!?_�u|��@����ٿ�|Ro�@�����3@{8,�!?_�u|��@����ٿ�|Ro�@�����3@{8,�!?_�u|��@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@�q32�ٿ�h�@��@ړ<�3@�j��D�!?�S�b�F�@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@8ƶ��ٿ��ַ�^�@/��_I�3@�{�H7�!?�P�<��@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@T��Y�ٿKh��-�@��� �3@��ӑg�!?�K^�@��w��ٿ=B4Za��@=�\�3@y0�F�!?;�u�nϴ@��w��ٿ=B4Za��@=�\�3@y0�F�!?;�u�nϴ@�x�u�ٿ���a��@/I<� 4@1y���!?_v��ʴ@�x�u�ٿ���a��@/I<� 4@1y���!?_v��ʴ@�x�u�ٿ���a��@/I<� 4@1y���!?_v��ʴ@�x�u�ٿ���a��@/I<� 4@1y���!?_v��ʴ@P�җٿ`߭Bx��@�ŭ�4@w�Q�c�!?sQ�#�@P�җٿ`߭Bx��@�ŭ�4@w�Q�c�!?sQ�#�@�*͠�ٿ��m��@c�O�w�3@�\�<�!?U���@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@!��X�ٿ�ٙ�e�@x��p�3@�u���!?�\.τߴ@�<N�ٿ�4���@�ìW_�3@0�|E�!?��6Ix.�@�<N�ٿ�4���@�ìW_�3@0�|E�!?��6Ix.�@�<N�ٿ�4���@�ìW_�3@0�|E�!?��6Ix.�@ jjx��ٿj�Ƃ"�@#�_:)�3@�(<xG�!?k��@ jjx��ٿj�Ƃ"�@#�_:)�3@�(<xG�!?k��@ܫ��[�ٿ��^�\��@ω���3@�M}�?�!?z�h����@ܫ��[�ٿ��^�\��@ω���3@�M}�?�!?z�h����@ܫ��[�ٿ��^�\��@ω���3@�M}�?�!?z�h����@F�p��ٿJ�M�@�jw3�3@�/��K�!?�bS��µ@F�p��ٿJ�M�@�jw3�3@�/��K�!?�bS��µ@aAR���ٿm/v1�r�@�����3@�q�tڏ!?����".�@�F����ٿ��/M�@��W,^�3@��}]ݏ!?��%�RL�@�F����ٿ��/M�@��W,^�3@��}]ݏ!?��%�RL�@�F����ٿ��/M�@��W,^�3@��}]ݏ!?��%�RL�@�F����ٿ��/M�@��W,^�3@��}]ݏ!?��%�RL�@�i7Dٿ�b����@qڐ��3@�UG��!?�թ�r��@{<M��ٿ"�5|���@�E��]�3@Nj��T�!?܄9#�@{<M��ٿ"�5|���@�E��]�3@Nj��T�!?܄9#�@{<M��ٿ"�5|���@�E��]�3@Nj��T�!?܄9#�@{<M��ٿ"�5|���@�E��]�3@Nj��T�!?܄9#�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�U~tn�ٿ���?N%�@��t|�3@��7�X�!?�s�1�@�/�9�ٿń��t��@�Sq��4@Źk�8�!?��%w��@�/�9�ٿń��t��@�Sq��4@Źk�8�!?��%w��@���_�ٿ�� _~��@q�0��3@�QqK�!?I�?��@���_�ٿ�� _~��@q�0��3@�QqK�!?I�?��@���_�ٿ�� _~��@q�0��3@�QqK�!?I�?��@���_�ٿ�� _~��@q�0��3@�QqK�!?I�?��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@#o�іٿbL
,��@ڀ���3@�)ތ��!?	}j��@��b�ٿ�H��@��C`�3@���Li�!?����$�@��b�ٿ�H��@��C`�3@���Li�!?����$�@��b�ٿ�H��@��C`�3@���Li�!?����$�@��b�ٿ�H��@��C`�3@���Li�!?����$�@3��t�ٿk:��]��@Q���4@s�8�!?��܊�@�멑ʎٿ�=�B��@DFƣ4@� זp�!?�As���@�멑ʎٿ�=�B��@DFƣ4@� זp�!?�As���@����ٿx�B�L��@�Ԕ�~4@�|{{�!?��ѹִ@\A#��ٿ�1b�*�@5��|�3@�F̟!�!?����N��@"��e��ٿu8eB�a�@��bR��3@�� �!?���^��@"��e��ٿu8eB�a�@��bR��3@�� �!?���^��@"��e��ٿu8eB�a�@��bR��3@�� �!?���^��@th��ٿݱ�����@6�>��3@q`�!?o�fQ�@th��ٿݱ�����@6�>��3@q`�!?o�fQ�@th��ٿݱ�����@6�>��3@q`�!?o�fQ�@���a��ٿ�k��ԃ�@���34@��*J�!?���>^�@���a��ٿ�k��ԃ�@���34@��*J�!?���>^�@���a��ٿ�k��ԃ�@���34@��*J�!?���>^�@���a��ٿ�k��ԃ�@���34@��*J�!?���>^�@�ۣ��ٿN���#�@?
4@74�W�!?��W��d�@�ۣ��ٿN���#�@?
4@74�W�!?��W��d�@��=I�ٿ��oK�p�@�:�c'�3@��6-�!?ng�B��@v��Hw�ٿ!OXT���@����t�3@�|�ZQ�!?[���Vٵ@v��Hw�ٿ!OXT���@����t�3@�|�ZQ�!?[���Vٵ@v��Hw�ٿ!OXT���@����t�3@�|�ZQ�!?[���Vٵ@v��Hw�ٿ!OXT���@����t�3@�|�ZQ�!?[���Vٵ@v��Hw�ٿ!OXT���@����t�3@�|�ZQ�!?[���Vٵ@
�js��ٿ�[�3���@fB���3@��C�W�!?�������@���ԏٿNQQ~��@P(L;��3@R�g$d�!?�~�5뎵@�%w%��ٿ"��;�[�@z�8�p4@���l�!?V��ly�@�m���ٿ�
����@�3���3@gݚ9��!?�R��v�@�m���ٿ�
����@�3���3@gݚ9��!?�R��v�@�m���ٿ�
����@�3���3@gݚ9��!?�R��v�@�m���ٿ�
����@�3���3@gݚ9��!?�R��v�@���q�ٿ�Y���C�@X�v��3@�>S��!?F�x��#�@���q�ٿ�Y���C�@X�v��3@�>S��!?F�x��#�@���q�ٿ�Y���C�@X�v��3@�>S��!?F�x��#�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@c0;5��ٿmDA��@z~@��3@w'S6�!?r�!n�@Ǯ��V�ٿY�:YH�@�0\��3@>�e�R�!?S+=�δ@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@z��-��ٿ������@^����3@�w�fW�!?������@��"�یٿ��4��@���,�3@��D1��!?M�Q�]�@F�x��ٿS�	s\��@�܋�4@��U���!?srG2�B�@C�C�ٿ�nv�f<�@��c4@�CME��!?��&P�O�@C�C�ٿ�nv�f<�@��c4@�CME��!?��&P�O�@C�C�ٿ�nv�f<�@��c4@�CME��!?��&P�O�@C�C�ٿ�nv�f<�@��c4@�CME��!?��&P�O�@C�C�ٿ�nv�f<�@��c4@�CME��!?��&P�O�@�g-�ؑٿBH�		�@q=&��3@7�Z��!?r�� $�@�g-�ؑٿBH�		�@q=&��3@7�Z��!?r�� $�@�g-�ؑٿBH�		�@q=&��3@7�Z��!?r�� $�@�g-�ؑٿBH�		�@q=&��3@7�Z��!?r�� $�@�����ٿo��w1�@mܖ}4@�L��F�!?�����I�@��"�l�ٿ#�a@"/�@WO�.��3@��;
�!?�`����@��"�l�ٿ#�a@"/�@WO�.��3@��;
�!?�`����@��"�l�ٿ#�a@"/�@WO�.��3@��;
�!?�`����@��"�l�ٿ#�a@"/�@WO�.��3@��;
�!?�`����@��~��ٿ_�.���@�X��.�3@��Η2�!?Ι*=z�@��~��ٿ_�.���@�X��.�3@��Η2�!?Ι*=z�@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@1
���ٿ��1�yh�@����1�3@����I�!?'������@�핊�ٿ�P�N���@�@T��3@�[��!?}�7�Ŵ@�핊�ٿ�P�N���@�@T��3@�[��!?}�7�Ŵ@�핊�ٿ�P�N���@�@T��3@�[��!?}�7�Ŵ@�핊�ٿ�P�N���@�@T��3@�[��!?}�7�Ŵ@�핊�ٿ�P�N���@�@T��3@�[��!?}�7�Ŵ@�n0�"�ٿ�42���@�����3@�ϯ �!?l%�@u�@8�+̏ٿ �"d�U�@#Pt�A�3@�ACKS�!?�ς�r�@8�+̏ٿ �"d�U�@#Pt�A�3@�ACKS�!?�ς�r�@8�+̏ٿ �"d�U�@#Pt�A�3@�ACKS�!?�ς�r�@�'�w�ٿ��t
���@Z���3@�Юy��!?�g��y�@�'�w�ٿ��t
���@Z���3@�Юy��!?�g��y�@�'�w�ٿ��t
���@Z���3@�Юy��!?�g��y�@��iߕٿI�-$��@x�H��3@vyf��!?2M>}!��@��iߕٿI�-$��@x�H��3@vyf��!?2M>}!��@Ps��ٿ���~f�@Qw魫�3@�c�m �!?}��K���@Ps��ٿ���~f�@Qw魫�3@�c�m �!?}��K���@Ps��ٿ���~f�@Qw魫�3@�c�m �!?}��K���@Ps��ٿ���~f�@Qw魫�3@�c�m �!?}��K���@ݛ�3��ٿؤ�E�@��M�3@��9N��!?k,y"�@ݛ�3��ٿؤ�E�@��M�3@��9N��!?k,y"�@ݛ�3��ٿؤ�E�@��M�3@��9N��!?k,y"�@^/��ٿ�|��@�2����3@f�>��!?��G�t �@^/��ٿ�|��@�2����3@f�>��!?��G�t �@^/��ٿ�|��@�2����3@f�>��!?��G�t �@r�u��ٿm���tL�@2���� 4@����$�!?��F䬴@r�u��ٿm���tL�@2���� 4@����$�!?��F䬴@r�u��ٿm���tL�@2���� 4@����$�!?��F䬴@r�u��ٿm���tL�@2���� 4@����$�!?��F䬴@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@*�Y�<�ٿ�Ԃ�3�@)�UW�4@�"1.�!?��e)+�@�t� �ٿ S]J]��@"��4@(P�[�!?�M=o�ٴ@�t� �ٿ S]J]��@"��4@(P�[�!?�M=o�ٴ@�t� �ٿ S]J]��@"��4@(P�[�!?�M=o�ٴ@�t� �ٿ S]J]��@"��4@(P�[�!?�M=o�ٴ@�t� �ٿ S]J]��@"��4@(P�[�!?�M=o�ٴ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@��I�^�ٿ����4r�@q���3@�AȜ+�!?��|��Ѵ@�䜨X�ٿ��}���@Te㖄�3@�M�3�!?����x�@�䜨X�ٿ��}���@Te㖄�3@�M�3�!?����x�@|��:�ٿ0��A���@��{F��3@��9Y1�!?�6�x6��@|��:�ٿ0��A���@��{F��3@��9Y1�!?�6�x6��@|��:�ٿ0��A���@��{F��3@��9Y1�!?�6�x6��@|��:�ٿ0��A���@��{F��3@��9Y1�!?�6�x6��@�ѭӸ�ٿZ�d`�f�@��DB�3@A ��!?і�[ȼ�@�ѭӸ�ٿZ�d`�f�@��DB�3@A ��!?і�[ȼ�@�ѭӸ�ٿZ�d`�f�@��DB�3@A ��!?і�[ȼ�@�ѭӸ�ٿZ�d`�f�@��DB�3@A ��!?і�[ȼ�@eͫ�ٿ�^E::�@'e���3@ay���!?�����@eͫ�ٿ�^E::�@'e���3@ay���!?�����@e���I�ٿ��]��#�@��{�3@�P�4�!?��~�r�@e���I�ٿ��]��#�@��{�3@�P�4�!?��~�r�@e���I�ٿ��]��#�@��{�3@�P�4�!?��~�r�@���ٿ�}��	��@�͠�3@mq���!?z7�+��@���ٿ�}��	��@�͠�3@mq���!?z7�+��@���ٿ�}��	��@�͠�3@mq���!?z7�+��@���ٿ�}��	��@�͠�3@mq���!?z7�+��@���ٿ�}��	��@�͠�3@mq���!?z7�+��@i"
nd�ٿ��)�i�@��\�3@���!?�̼,��@i"
nd�ٿ��)�i�@��\�3@���!?�̼,��@d|U�+�ٿj������@��L	�3@���!h�!?�
��@�s��ٿ�C �r�@�8��3@�)���!?Ky<�C��@�s��ٿ�C �r�@�8��3@�)���!?Ky<�C��@�s��ٿ�C �r�@�8��3@�)���!?Ky<�C��@�s��ٿ�C �r�@�8��3@�)���!?Ky<�C��@�s��ٿ�C �r�@�8��3@�)���!?Ky<�C��@�g�O��ٿ���>`�@��S��3@aqnH�!?�bWq���@�g�O��ٿ���>`�@��S��3@aqnH�!?�bWq���@�g�O��ٿ���>`�@��S��3@aqnH�!?�bWq���@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@Db#�[�ٿ��jv��@�Wfu�3@=ͯ`�!?�>sL�@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@+��[�ٿl�Ļ�@U�K��3@�3:I$�!?`��c��@M�逛�ٿ=������@tv_���3@����.�!?c�-x�@M�逛�ٿ=������@tv_���3@����.�!?c�-x�@M�逛�ٿ=������@tv_���3@����.�!?c�-x�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@��z�|�ٿ��P���@��m���3@!��F)�!?c�j>�1�@t2���ٿ��4W�@��Z�4@cخ6r�!?D��b3��@�ϋ:�ٿ(��B�@J�z�4@n���!?�|��_�@�ϋ:�ٿ(��B�@J�z�4@n���!?�|��_�@�ϋ:�ٿ(��B�@J�z�4@n���!?�|��_�@Tֆ���ٿ��t���@�O��3@�{���!?�,#�=�@Tֆ���ٿ��t���@�O��3@�{���!?�,#�=�@Tֆ���ٿ��t���@�O��3@�{���!?�,#�=�@Tֆ���ٿ��t���@�O��3@�{���!?�,#�=�@Tֆ���ٿ��t���@�O��3@�{���!?�,#�=�@����ٿ�`<���@ P6Q�3@ư>Q�!?�NGݢQ�@����ٿ�`<���@ P6Q�3@ư>Q�!?�NGݢQ�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@F�i���ٿ��q��@Ch�҂�3@��{�K�!?�ȁ�D1�@y�O�ٿ>#�`1�@C��N��3@�m]P�!?P����@y�O�ٿ>#�`1�@C��N��3@�m]P�!?P����@�Zt�ڞٿjFj�[�@��I��3@Q�2��!?��c�=�@�Zt�ڞٿjFj�[�@��I��3@Q�2��!?��c�=�@�Zt�ڞٿjFj�[�@��I��3@Q�2��!?��c�=�@�Zt�ڞٿjFj�[�@��I��3@Q�2��!?��c�=�@�hϞ��ٿ[h}��@5�&Q$�3@�B�!?�m�]��@�hϞ��ٿ[h}��@5�&Q$�3@�B�!?�m�]��@�hϞ��ٿ[h}��@5�&Q$�3@�B�!?�m�]��@�hϞ��ٿ[h}��@5�&Q$�3@�B�!?�m�]��@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@!<�;�ٿu�o��@]!�|�3@+_[2�!?,��h䴴@�Ԍԍ�ٿ�������@�*�-I�3@.��U�!? �q�a�@�Ԍԍ�ٿ�������@�*�-I�3@.��U�!? �q�a�@�Ԍԍ�ٿ�������@�*�-I�3@.��U�!? �q�a�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@���ٿ�{!���@/�	�|�3@�K���!?�JC-�@ӷ��+�ٿi�T��!�@4�н�3@��ؙ�!?yop�T5�@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@lV�ǀ�ٿ�d�y��@?z���3@�/�f�!?�m�8��@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@����Y�ٿ��`��@vm׽p�3@�3��M�!?viǊ�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@��Ü�ٿ�(�6<��@*�W�g�3@��!?H�'´s�@�d�R��ٿ��2����@!��VB�3@�m�%>�!?����@Xd�F�ٿY�%���@g����3@V�hnj�!?��N���@Xd�F�ٿY�%���@g����3@V�hnj�!?��N���@Xd�F�ٿY�%���@g����3@V�hnj�!?��N���@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@��M$�ٿ�K�#)��@t��
M�3@����^�!?�m��ڵ@9i2/��ٿDb�J�<�@J�	�:�3@ҁU]S�!?� �>µ@9i2/��ٿDb�J�<�@J�	�:�3@ҁU]S�!?� �>µ@�M��~�ٿ��H���@�[ȕR�3@����U�!?l�Бn �@4C����ٿ��m��@&�<��3@���2
�!?w�x+3�@req��ٿ������@~��H�3@sۢ�!?D���ģ�@s��CۚٿTm��f1�@Z�����3@��i>�!?�U󓎵@s��CۚٿTm��f1�@Z�����3@��i>�!?�U󓎵@s��CۚٿTm��f1�@Z�����3@��i>�!?�U󓎵@s��CۚٿTm��f1�@Z�����3@��i>�!?�U󓎵@s��CۚٿTm��f1�@Z�����3@��i>�!?�U󓎵@���ٿ�i�m3V�@�,�X��3@!�NLI�!?9�@q�@���ٿ�i�m3V�@�,�X��3@!�NLI�!?9�@q�@���ٿ�i�m3V�@�,�X��3@!�NLI�!?9�@q�@���ٿ�i�m3V�@�,�X��3@!�NLI�!?9�@q�@���ٿ�i�m3V�@�,�X��3@!�NLI�!?9�@q�@M!a�ٿ��yy_�@��G��3@'<��x�!?�S?z�@M!a�ٿ��yy_�@��G��3@'<��x�!?�S?z�@��D"�ٿ9�����@@9B��3@<�6z\�!? #�ct;�@��t'��ٿ���ݤ�@�.A4@�xQZ�!?˃���@��/ĕٿHP�q�@�@n2B���3@��/�!?u�JD���@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@��Pk��ٿ���S�@qgq�b�3@>�v �!?R���m��@�`�J<�ٿɾ�|��@8�����3@nÆ�	�!?DxKad��@�`�J<�ٿɾ�|��@8�����3@nÆ�	�!?DxKad��@����˒ٿ�>|i�@����4@�A�^l�!?����q۴@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@`A;���ٿ���st�@�Z��#�3@º����!?@11w�b�@�wv�ٿc~����@�q��	4@����Q�!?�l�:�@�wv�ٿc~����@�q��	4@����Q�!?�l�:�@�wv�ٿc~����@�q��	4@����Q�!?�l�:�@�wv�ٿc~����@�q��	4@����Q�!?�l�:�@��]\��ٿ ٘�e��@�u�r�4@.�d�b�!?� 
�-��@��]\��ٿ ٘�e��@�u�r�4@.�d�b�!?� 
�-��@s��Ēٿ}��jۜ�@�ʽ4@ESf�J�!?:a�F��@s��Ēٿ}��jۜ�@�ʽ4@ESf�J�!?:a�F��@s��Ēٿ}��jۜ�@�ʽ4@ESf�J�!?:a�F��@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@���D�ٿIdw���@��G�4@�,jO�!?�� Ԧ�@��\�b�ٿ��c��a�@��w�4@���`�!?sK�^���@�`IP��ٿ�e�w�@���4@Ş�@��!?~ddFv�@-RG���ٿ�����@��3;��3@�>ې!?��8�@-RG���ٿ�����@��3;��3@�>ې!?��8�@-RG���ٿ�����@��3;��3@�>ې!?��8�@-RG���ٿ�����@��3;��3@�>ې!?��8�@�3����ٿ�AF�(s�@Mbhv� 4@1�����!?LDzٴ.�@�3����ٿ�AF�(s�@Mbhv� 4@1�����!?LDzٴ.�@�3����ٿ�AF�(s�@Mbhv� 4@1�����!?LDzٴ.�@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�<� S�ٿ�W���@�WB>9 4@�Ӗِ!?�ic����@�X�՞ٿ�l�"�@R�2[4@�6>�Ɛ!?*}�پ��@[�Y�Ġٿ5}�A���@~�7v4@Mo�s!�!?%&�K7�@�M	�ٿf��aw��@��xy24@��w�e�!?8�JP���@�M	�ٿf��aw��@��xy24@��w�e�!?8�JP���@��W��ٿ��K��@�����3@��l'�!?�B�F��@��W��ٿ��K��@�����3@��l'�!?�B�F��@��W��ٿ��K��@�����3@��l'�!?�B�F��@GO	�h�ٿ>Ԯ�Mz�@Ԧ2�>�3@���z�!?I���l�@i1�l��ٿ�����@�(����3@}���!?a�݊:��@i1�l��ٿ�����@�(����3@}���!?a�݊:��@��:ض�ٿ6É�m��@S�A�t�3@����G�!?��/w�A�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@*`���ٿ������@�:5�3@������!?Q�i�H�@�W*�ܚٿ�J�*y�@���,��3@p�*/�!?�\t�;�@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@���ٿUa!H��@D��k*�3@D6�"�!?�e]̴@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@]E�w�ٿ3m9� �@!���;�3@��8�!?�:��@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@zA�F�ٿCm�M�k�@"s�c�3@�`Љ#�!?�8͚�7�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@�-��Ǔٿ$ΐ=˱�@�&9OH�3@�OKF�!?���s�@��oy�ٿ�L-B<i�@k�{nE�3@���hw�!?�K�u��@��oy�ٿ�L-B<i�@k�{nE�3@���hw�!?�K�u��@��oy�ٿ�L-B<i�@k�{nE�3@���hw�!?�K�u��@��oy�ٿ�L-B<i�@k�{nE�3@���hw�!?�K�u��@��oy�ٿ�L-B<i�@k�{nE�3@���hw�!?�K�u��@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@��y�ٿ A�k�@)z���3@����!?��esϴ@x��N��ٿXm5���@q�z�4@��ޑG�!?5XF
$�@x��N��ٿXm5���@q�z�4@��ޑG�!?5XF
$�@x��N��ٿXm5���@q�z�4@��ޑG�!?5XF
$�@x��N��ٿXm5���@q�z�4@��ޑG�!?5XF
$�@x��N��ٿXm5���@q�z�4@��ޑG�!?5XF
$�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@��r�#�ٿ��.߆��@lmqƨ4@߬�V�!?�G�%E�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@�����ٿ�J�?��@�GܲU�3@RI��!?�:
�@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@���P�ٿ��_��@�qOF�3@��}!�!?J���ꤴ@;Z訜�ٿ��y��@�*���3@��A�!?�@|.��@7�{x<�ٿ1υ���@�`\��4@
W��:�!?�M�y���@7�{x<�ٿ1υ���@�`\��4@
W��:�!?�M�y���@7�{x<�ٿ1υ���@�`\��4@
W��:�!?�M�y���@�U�8�ٿY���7�@W��WQ4@T?����!?��ӊ`�@�U�8�ٿY���7�@W��WQ4@T?����!?��ӊ`�@�ò*��ٿ0�@%t�@�8M��3@Ɯ^�t�!?�@��(��@�ò*��ٿ0�@%t�@�8M��3@Ɯ^�t�!?�@��(��@�ò*��ٿ0�@%t�@�8M��3@Ɯ^�t�!?�@��(��@�ò*��ٿ0�@%t�@�8M��3@Ɯ^�t�!?�@��(��@�ò*��ٿ0�@%t�@�8M��3@Ɯ^�t�!?�@��(��@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@!B<�ٿR �Q`n�@��\F�4@\g��}�!?�H���@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�6���ٿ�L�#��@���>4@���KP�!?0h�-�@�gI�=�ٿ��M�@B��{�3@-��7�!?�t+k��@�gI�=�ٿ��M�@B��{�3@-��7�!?�t+k��@��Ű�ٿ? ��5.�@�.���3@�-ET�!?\�:F�@��Ű�ٿ? ��5.�@�.���3@�-ET�!?\�:F�@w���טٿPk��e�@5���K�3@4�^�!?ᚃ#t3�@w���טٿPk��e�@5���K�3@4�^�!?ᚃ#t3�@�/]�ٿ�!h�t�@Z���3@yĶ�!?��JiSմ@Ox�yr�ٿޝNk��@�����3@����!?P���&�@Ox�yr�ٿޝNk��@�����3@����!?P���&�@�r8/r�ٿ������@ؐ��F�3@v>�֏!?�����@�r8/r�ٿ������@ؐ��F�3@v>�֏!?�����@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@r�7��ٿ��g�O��@^��^x�3@OB
�!?�v2��@����t�ٿ��9���@g�V8��3@��O�!?�Z�q b�@����t�ٿ��9���@g�V8��3@��O�!?�Z�q b�@����t�ٿ��9���@g�V8��3@��O�!?�Z�q b�@����t�ٿ��9���@g�V8��3@��O�!?�Z�q b�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@�v� �ٿ��1�"t�@�o=���3@(�i6O�!?�@Rt�T�@tpK��ٿ���H�3�@�J��#4@�����!?���`Z�@����Q�ٿ��J�[
�@%�T��4@ͷt~��!?C�f"۴@����Q�ٿ��J�[
�@%�T��4@ͷt~��!?C�f"۴@����Q�ٿ��J�[
�@%�T��4@ͷt~��!?C�f"۴@����Q�ٿ��J�[
�@%�T��4@ͷt~��!?C�f"۴@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@9��1�ٿ��cY��@#���4@ #�!?xq�=�@�3i��ٿ���hk%�@}�zM4@��j�!?0�݀��@�3i��ٿ���hk%�@}�zM4@��j�!?0�݀��@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@��w�	�ٿq���o�@�4@[IJ�!?��6-���@���#��ٿ3���p�@������3@"�R�!?��d�p�@���#��ٿ3���p�@������3@"�R�!?��d�p�@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@<?�7��ٿ|����`�@��|W��3@X3�7�!?�����@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@�����ٿ|��3Z�@V��(�3@���S�!?*���y�@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@��(��ٿ��V���@y{�V��3@����z�!?�e�Q,��@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@G�|n�ٿ�˥�?��@)(��3@���]R�!?q�D�> �@�cS�a�ٿ�3����@�HBA<�3@����i�!?��^�.�@�cS�a�ٿ�3����@�HBA<�3@����i�!?��^�.�@�&ά�ٿ{�7^��@h�'R�3@��9=D�!?�}�q2�@�&ά�ٿ{�7^��@h�'R�3@��9=D�!?�}�q2�@�&ά�ٿ{�7^��@h�'R�3@��9=D�!?�}�q2�@��f�ٿ��X�'�@�Ú˫�3@_@1���!?f��q��@��f�ٿ��X�'�@�Ú˫�3@_@1���!?f��q��@�c�J�ٿk��֥�@��:��3@�*�8�!?��ʔ�@�c�J�ٿk��֥�@��:��3@�*�8�!?��ʔ�@iwg��ٿ2Yd����@��|s�3@nSD���!?M�Nr2~�@iwg��ٿ2Yd����@��|s�3@nSD���!?M�Nr2~�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@�Y��Жٿ����@�i��m�3@������!?�Am�<-�@ݮV�T�ٿ����֥�@����4@7�u�!?qrݨ�G�@ݮV�T�ٿ����֥�@����4@7�u�!?qrݨ�G�@���{!�ٿ��C�D�@c ��44@ZsmR�!?h����ε@���{!�ٿ��C�D�@c ��44@ZsmR�!?h����ε@���{!�ٿ��C�D�@c ��44@ZsmR�!?h����ε@���{!�ٿ��C�D�@c ��44@ZsmR�!?h����ε@k^�~>�ٿl?B\�|�@�p���3@��z�k�!?\`,�J\�@k^�~>�ٿl?B\�|�@�p���3@��z�k�!?\`,�J\�@k^�~>�ٿl?B\�|�@�p���3@��z�k�!?\`,�J\�@22u0�ٿ�����$�@+��+4@�-��}�!?�E�Ҩ�@ˑx�r�ٿR�����@�'���4@)>�Ð!?_�R��@ˑx�r�ٿR�����@�'���4@)>�Ð!?_�R��@ˑx�r�ٿR�����@�'���4@)>�Ð!?_�R��@��C{�ٿ�Bg|5�@����3@���ξ�!?���NR�@��C{�ٿ�Bg|5�@����3@���ξ�!?���NR�@R�8�]�ٿ�7�8��@�s��4@xT慩�!?W-�Ǔ0�@R�8�]�ٿ�7�8��@�s��4@xT慩�!?W-�Ǔ0�@R�8�]�ٿ�7�8��@�s��4@xT慩�!?W-�Ǔ0�@R�8�]�ٿ�7�8��@�s��4@xT慩�!?W-�Ǔ0�@R�8�]�ٿ�7�8��@�s��4@xT慩�!?W-�Ǔ0�@�E&9S�ٿ+��V�@�W	U��3@r��ki�!?f����@�E&9S�ٿ+��V�@�W	U��3@r��ki�!?f����@Um��m�ٿ��$��v�@Qӫ�3@�.�J��!?������@Um��m�ٿ��$��v�@Qӫ�3@�.�J��!?������@���to�ٿ"K��K�@�JI)�3@�p�O�!?m��$v�@	�e�{�ٿ�r�P�@5�i
�3@'K����!?�o77�@	�e�{�ٿ�r�P�@5�i
�3@'K����!?�o77�@$U����ٿ}��ۑ�@{�_���3@�Ơ�e�!?Us��4�@g5�]�ٿ�1����@8�Q�F�3@%�M�L�!?~�Ktp��@�w��ٿxҳ�0��@�r�a4@Ky�FH�!?f���lδ@�w��ٿxҳ�0��@�r�a4@Ky�FH�!?f���lδ@�w��ٿxҳ�0��@�r�a4@Ky�FH�!?f���lδ@�w��ٿxҳ�0��@�r�a4@Ky�FH�!?f���lδ@�w��ٿxҳ�0��@�r�a4@Ky�FH�!?f���lδ@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@[��t�ٿ���4,�@�^���3@֮��1�!?[;qGvd�@+aÃ�ٿ�3�g���@w񡿧�3@[s�'�!?�E�X�@+aÃ�ٿ�3�g���@w񡿧�3@[s�'�!?�E�X�@z�v�ٿ�{�h5x�@�>C��3@�X��J�!?Ǯe���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@၏��ٿX����f�@��;��3@��`�O�!?:�A5���@��6O�ٿ���f[;�@�� �3@�6*��!?�]�ZH�@��6O�ٿ���f[;�@�� �3@�6*��!?�]�ZH�@��6O�ٿ���f[;�@�� �3@�6*��!?�]�ZH�@��A�ٿD�:ၣ�@�"YV�3@��e.�!?]� ��@��A�ٿD�:ၣ�@�"YV�3@��e.�!?]� ��@��A�ٿD�:ၣ�@�"YV�3@��e.�!?]� ��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@iF>���ٿmA&�k�@�!���3@����!?��tkU��@1LeՙٿBǬ6�@)�ZH�3@���V�!?���m�@1LeՙٿBǬ6�@)�ZH�3@���V�!?���m�@���<2�ٿ�t����@�����3@��GG�!?��q`���@���<2�ٿ�t����@�����3@��GG�!?��q`���@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@U�y�I�ٿ�j�QX�@��<�2�3@���!?���|��@��ۺ�ٿ�q�^��@���@��3@'_5=�!?���d���@��ۺ�ٿ�q�^��@���@��3@'_5=�!?���d���@��ۺ�ٿ�q�^��@���@��3@'_5=�!?���d���@��ۺ�ٿ�q�^��@���@��3@'_5=�!?���d���@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@v�(���ٿ��R���@R��$S�3@j�(�!?'<�9H�@��&J�ٿ8�&�|�@'���#�3@��_�b�!?e@�q���@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@��l+ٕٿ>����@�f9u� 4@䙿!�!?He��H��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@�Vd���ٿ/٤{�l�@�����	4@��"�!?9�g�Z��@:M����ٿ�-c�V�@E7�d�4@�4�6�!?�������@
�)]�ٿ߽	�4��@�M����3@�68�!?������@
�)]�ٿ߽	�4��@�M����3@�68�!?������@
�)]�ٿ߽	�4��@�M����3@�68�!?������@
�)]�ٿ߽	�4��@�M����3@�68�!?������@���a��ٿ�v�g2�@*����3@$(��)�!?x)�־�@���a��ٿ�v�g2�@*����3@$(��)�!?x)�־�@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@�S���ٿ\��!A��@p�_�3@����;�!?�!v_���@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@mp�ǉ�ٿ�1J�E�@���3@���|>�!?���;{�@���`3�ٿ�vS�3�@(�]�9�3@�W��}�!?�Q�7*��@���`3�ٿ�vS�3�@(�]�9�3@�W��}�!?�Q�7*��@���`3�ٿ�vS�3�@(�]�9�3@�W��}�!?�Q�7*��@���`3�ٿ�vS�3�@(�]�9�3@�W��}�!?�Q�7*��@�?�֗ٿ$��V�o�@3
@!�3@�2��1�!?L�j��m�@|-\��ٿ�Pm�@�¥,�3@W2�`�!?��	mn�@|-\��ٿ�Pm�@�¥,�3@W2�`�!?��	mn�@|-\��ٿ�Pm�@�¥,�3@W2�`�!?��	mn�@Sj�sp�ٿJĵ�8d�@��c�3@k��z�!?��lόw�@Sj�sp�ٿJĵ�8d�@��c�3@k��z�!?��lόw�@Sj�sp�ٿJĵ�8d�@��c�3@k��z�!?��lόw�@Sj�sp�ٿJĵ�8d�@��c�3@k��z�!?��lόw�@obלٿQW뾿��@��R�3@G.]W�!?�Q 5�@obלٿQW뾿��@��R�3@G.]W�!?�Q 5�@obלٿQW뾿��@��R�3@G.]W�!?�Q 5�@obלٿQW뾿��@��R�3@G.]W�!?�Q 5�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���b��ٿG�Û,+�@]<���3@����!?�{ L8�@���<P�ٿ�g(}
��@${^��3@0f��1�!?���C�y�@���<P�ٿ�g(}
��@${^��3@0f��1�!?���C�y�@���<P�ٿ�g(}
��@${^��3@0f��1�!?���C�y�@�J�'�ٿ/T-����@*��sY4@oq/���!?s��@�J�'�ٿ/T-����@*��sY4@oq/���!?s��@�J�'�ٿ/T-����@*��sY4@oq/���!?s��@�J�'�ٿ/T-����@*��sY4@oq/���!?s��@�J�'�ٿ/T-����@*��sY4@oq/���!?s��@�Gע�ٿ���oZ?�@�me�y�3@_"l� �!?���L��@�Gע�ٿ���oZ?�@�me�y�3@_"l� �!?���L��@�Gע�ٿ���oZ?�@�me�y�3@_"l� �!?���L��@�Gע�ٿ���oZ?�@�me�y�3@_"l� �!?���L��@��
��ٿg�����@-Eӫ��3@���'�!?n�q8G��@��
��ٿg�����@-Eӫ��3@���'�!?n�q8G��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@)ʚ�m�ٿ�*y�z
�@��섀�3@wK�`)�!?o�9�B��@��'	מٿ�]=�r�@W��T��3@ِ$�?�!?=�(R�@��'	מٿ�]=�r�@W��T��3@ِ$�?�!?=�(R�@��'	מٿ�]=�r�@W��T��3@ِ$�?�!?=�(R�@��'	מٿ�]=�r�@W��T��3@ِ$�?�!?=�(R�@�c뙻�ٿt�WE��@t�����3@�')�!?b��[ĵ@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@C��/�ٿ��J���@��s�q�3@�����!?���\6��@�t^���ٿ,��/��@�_p���3@=���!?�����@�t^���ٿ,��/��@�_p���3@=���!?�����@�t^���ٿ,��/��@�_p���3@=���!?�����@�t^���ٿ,��/��@�_p���3@=���!?�����@�t^���ٿ,��/��@�_p���3@=���!?�����@6�#5A�ٿ�"f���@b-��3@�8����!?���G�@6�#5A�ٿ�"f���@b-��3@�8����!?���G�@6�#5A�ٿ�"f���@b-��3@�8����!?���G�@6�#5A�ٿ�"f���@b-��3@�8����!?���G�@0>���ٿҘi��r�@�܊�:�3@�`�!?L��F�@0>���ٿҘi��r�@�܊�:�3@�`�!?L��F�@0>���ٿҘi��r�@�܊�:�3@�`�!?L��F�@0>���ٿҘi��r�@�܊�:�3@�`�!?L��F�@0>���ٿҘi��r�@�܊�:�3@�`�!?L��F�@O �%��ٿ���y�@�%�3@�<��,�!?l���@O �%��ٿ���y�@�%�3@�<��,�!?l���@O �%��ٿ���y�@�%�3@�<��,�!?l���@Ś?���ٿ��g_8��@�]+���3@�׺Q�!?q[>?�@Ś?���ٿ��g_8��@�]+���3@�׺Q�!?q[>?�@bN[`G�ٿ-5O��@�C�*g�3@���ro�!?d���
�@bN[`G�ٿ-5O��@�C�*g�3@���ro�!?d���
�@bN[`G�ٿ-5O��@�C�*g�3@���ro�!?d���
�@��>��ٿ���Q���@,�p�� 4@��3�H�!?�O��6-�@[&w	��ٿL@Q�J��@jR��04@�
�'[�!?��`�أ�@[&w	��ٿL@Q�J��@jR��04@�
�'[�!?��`�أ�@���T��ٿ�~Tڦ��@�TA�v�3@�_���!?�0I���@���T��ٿ�~Tڦ��@�TA�v�3@�_���!?�0I���@���T��ٿ�~Tڦ��@�TA�v�3@�_���!?�0I���@�0�L+�ٿ�84C���@-y�5o4@�!��M�!?�]���@��K���ٿ��,����@��ȨG4@/,�u�!?zc�>�=�@���x�ٿ�x���}�@f�����3@>���M�!?���(|J�@�w�>�ٿZ�Y�A��@�f���3@����2�!?�ˊ��@�w�>�ٿZ�Y�A��@�f���3@����2�!?�ˊ��@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@��"���ٿ5'[�0�@7�Z7��3@��A�!?nj��ɴ@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@[p�t�ٿ�`e9��@1��Y��3@��f��!?������@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@@�S�D�ٿ�tN=�@��_�[4@�^�B�!?�m�6��@�x��ǘٿ;(�ٛ�@�l����3@����!?��2�@�x��ǘٿ;(�ٛ�@�l����3@����!?��2�@~e�p��ٿڼ�\n��@5�8��3@��f�8�!?zʕ\Y�@��ы؟ٿ�[O����@`�>��3@&�,�!?��HnH�@��ы؟ٿ�[O����@`�>��3@&�,�!?��HnH�@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@�+��ėٿ]���O�@�e�3@��;���!?�/�ε@9��D�ٿm��IFk�@��*��3@��X�q�!?�t�ζ�@9��D�ٿm��IFk�@��*��3@��X�q�!?�t�ζ�@��fP�ٿ� �n��@w�|.�3@zsv�!?�S�s�S�@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@��s�ٿ�oj��@�����3@G�y�!?&�7��@;>R���ٿvO'��@ �.J�3@b&��7�!?�O���/�@	s��ٿ����/�@�7���3@С��W�!?�:o4�@	s��ٿ����/�@�7���3@С��W�!?�:o4�@	s��ٿ����/�@�7���3@С��W�!?�:o4�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@c��ٿ~��7���@4ܙpy4@߇�M�!?��3L�@���/�ٿ�_R]��@����4@�L��5�!?>8�Eִ@���/�ٿ�_R]��@����4@�L��5�!?>8�Eִ@�A�"<�ٿR�HZ�L�@t�u���3@f�WA��!?P(�����@�A�"<�ٿR�HZ�L�@t�u���3@f�WA��!?P(�����@�A�"<�ٿR�HZ�L�@t�u���3@f�WA��!?P(�����@�A�"<�ٿR�HZ�L�@t�u���3@f�WA��!?P(�����@�3�p�ٿiA��(�@�8p�-�3@���!?�G���@�3�p�ٿiA��(�@�8p�-�3@���!?�G���@�3�p�ٿiA��(�@�8p�-�3@���!?�G���@�3�p�ٿiA��(�@�8p�-�3@���!?�G���@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@=����ٿXd����@��1؈4@����%�!?��bBm�@���ٿ��O�'�@�vʦ�3@��l��!?�d�%��@���ٿ��O�'�@�vʦ�3@��l��!?�d�%��@���ٿ��O�'�@�vʦ�3@��l��!?�d�%��@���ٿ��O�'�@�vʦ�3@��l��!?�d�%��@�/��ٿF����@a����3@|͠-�!?.��%���@�/��ٿF����@a����3@|͠-�!?.��%���@�*=�ٿ"cDWs�@�{N�3@���7�!?=$�7?\�@�*=�ٿ"cDWs�@�{N�3@���7�!?=$�7?\�@�*=�ٿ"cDWs�@�{N�3@���7�!?=$�7?\�@zx<1�ٿ��B��@7�q���3@c{U�8�!?	Z�5��@zx<1�ٿ��B��@7�q���3@c{U�8�!?	Z�5��@zx<1�ٿ��B��@7�q���3@c{U�8�!?	Z�5��@zx<1�ٿ��B��@7�q���3@c{U�8�!?	Z�5��@zx<1�ٿ��B��@7�q���3@c{U�8�!?	Z�5��@�w�ޕٿ�����@d=��c�3@�yGL:�!?0������@�w�ޕٿ�����@d=��c�3@�yGL:�!?0������@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@U���ٿ�taO���@�B�l�4@���D��!?�� ��@�eD	��ٿ8�\��@��c�n�3@fdԢ��!?������@�eD	��ٿ8�\��@��c�n�3@fdԢ��!?������@�eD	��ٿ8�\��@��c�n�3@fdԢ��!?������@���3�ٿ7Z:����@�YX��3@����!?k՛���@�&��ٿ��<l�^�@	�����3@�΃�N�!?�K�,�c�@�&��ٿ��<l�^�@	�����3@�΃�N�!?�K�,�c�@�&��ٿ��<l�^�@	�����3@�΃�N�!?�K�,�c�@�&��ٿ��<l�^�@	�����3@�΃�N�!?�K�,�c�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@d�����ٿ�0���@s2<��3@��z0ݏ!?����(�@�*;�I�ٿ]g��֞�@>� t�3@aI%�!?=����ٴ@�:��r�ٿ::u#mh�@��9 4@0�ABW�!?��o��@��`�e�ٿv������@|��ۑ�3@��*s�!?c�����@̠���ٿT�I�L�@T�B< �3@���	�!?`�r{�@̠���ٿT�I�L�@T�B< �3@���	�!?`�r{�@̠���ٿT�I�L�@T�B< �3@���	�!?`�r{�@��X]��ٿ�J�e�y�@�:���3@��7�.�!?o^�.e�@��X]��ٿ�J�e�y�@�:���3@��7�.�!?o^�.e�@��X]��ٿ�J�e�y�@�:���3@��7�.�!?o^�.e�@ro<U�ٿ�|�>q��@������3@�AD�K�!?g�gP�G�@�yaV�ٿİ����@1�4�R�3@��q/�!?	���4��@�yaV�ٿİ����@1�4�R�3@��q/�!?	���4��@�yaV�ٿİ����@1�4�R�3@��q/�!?	���4��@�5���ٿ?k-�j��@ �S��3@L��Z�!?S�Nı�@�5���ٿ?k-�j��@ �S��3@L��Z�!?S�Nı�@�c���ٿ�0}�Y!�@VAO��3@�8\�V�!?�I.�m�@�c���ٿ�0}�Y!�@VAO��3@�8\�V�!?�I.�m�@�c���ٿ�0}�Y!�@VAO��3@�8\�V�!?�I.�m�@�c���ٿ�0}�Y!�@VAO��3@�8\�V�!?�I.�m�@�c���ٿ�0}�Y!�@VAO��3@�8\�V�!?�I.�m�@o3�P֝ٿ�cG<$�@�z)���3@2b)[�!?�D��=�@o3�P֝ٿ�cG<$�@�z)���3@2b)[�!?�D��=�@o3�P֝ٿ�cG<$�@�z)���3@2b)[�!?�D��=�@o3�P֝ٿ�cG<$�@�z)���3@2b)[�!?�D��=�@�2	���ٿ~�����@Uo�u�3@:ûQ�!?[�����@�2	���ٿ~�����@Uo�u�3@:ûQ�!?[�����@�2	���ٿ~�����@Uo�u�3@:ûQ�!?[�����@�2	���ٿ~�����@Uo�u�3@:ûQ�!?[�����@>�D��ٿ�4����@�&/x4@�~H$D�!?Ap�!:B�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@����c�ٿ�hK�a�@��]B(�3@�x(��!?��?P�*�@� �I�ٿB�[��k�@a3a@�3@���?�!?���W�@K�W�ٿh�n%��@|s֝J�3@M��F�!?��;E�~�@K�W�ٿh�n%��@|s֝J�3@M��F�!?��;E�~�@K�W�ٿh�n%��@|s֝J�3@M��F�!?��;E�~�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@h!�BF�ٿ���;�@@`�ί�3@��d�T�!?P��46I�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@d�	ٻ�ٿ裎9��@�>��3@Bа�_�!?�sr�?u�@��H`�ٿ��C�z�@���[4@�4UV�!?�L-,д@��H`�ٿ��C�z�@���[4@�4UV�!?�L-,д@��H`�ٿ��C�z�@���[4@�4UV�!?�L-,д@�CcP/�ٿ�m�ݜ]�@Yp�A�4@z�&��!?�咯��@�CcP/�ٿ�m�ݜ]�@Yp�A�4@z�&��!?�咯��@�CcP/�ٿ�m�ݜ]�@Yp�A�4@z�&��!?�咯��@�CcP/�ٿ�m�ݜ]�@Yp�A�4@z�&��!?�咯��@�CcP/�ٿ�m�ݜ]�@Yp�A�4@z�&��!?�咯��@�@���ٿ����87�@=	D�|�3@�����!?SN���Ӵ@j�6Ԓٿ�{�P*��@�ͥ^��3@�.H��!?ъ.~b�@j�6Ԓٿ�{�P*��@�ͥ^��3@�.H��!?ъ.~b�@j�6Ԓٿ�{�P*��@�ͥ^��3@�.H��!?ъ.~b�@j�6Ԓٿ�{�P*��@�ͥ^��3@�.H��!?ъ.~b�@)��q�ٿ��.2�B�@�<����3@�W�'�!?�t|a�Դ@)��q�ٿ��.2�B�@�<����3@�W�'�!?�t|a�Դ@)��q�ٿ��.2�B�@�<����3@�W�'�!?�t|a�Դ@�����ٿ�������@���΋4@p6q�X�!??���|m�@�����ٿ�������@���΋4@p6q�X�!??���|m�@D���J�ٿ�5��@�C���3@,ڤe�!?i��-�@D���J�ٿ�5��@�C���3@,ڤe�!?i��-�@	4�K��ٿ�.�Œ��@��y�U�3@����!?RS�Or;�@�G���ٿ��	���@�(C���3@�뾍�!?r�E#�@�G���ٿ��	���@�(C���3@�뾍�!?r�E#�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@���:�ٿ�\��C��@2����3@�:�j�!?n��ܛ�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@&��W]�ٿJ�,;���@#�3@��=�!?�?T��m�@z��67�ٿ�����@r"���4@�����!?����)�@z��67�ٿ�����@r"���4@�����!?����)�@n�^��ٿ+w
����@�X?;Y�3@;�vH�!?x��R|�@n�^��ٿ+w
����@�X?;Y�3@;�vH�!?x��R|�@ʁՂb�ٿ�P9��@��b 4�3@���$�!?�eHX
�@ʁՂb�ٿ�P9��@��b 4�3@���$�!?�eHX
�@3�R�	�ٿ��$���@7��P�3@������!?�^��f��@3�R�	�ٿ��$���@7��P�3@������!?�^��f��@�bٿ�B��
e�@��I��3@;vQ��!?|?�ݵ@�&i��ٿ�]ٛ�@��m�s�3@R*U��!?���28�@,��M��ٿ����@��9
��3@�ķY��!?��f��`�@,��M��ٿ����@��9
��3@�ķY��!?��f��`�@,��M��ٿ����@��9
��3@�ķY��!?��f��`�@*o�Z��ٿ�R-g'��@��@d�3@\sOJ�!?2�j�C��@�9�w�ٿ�uf��@��1�3@��d�;�!?�k�3���@�9�w�ٿ�uf��@��1�3@��d�;�!?�k�3���@�"@
�ٿ>�?�:l�@�j>nx	4@RD%��!?MC�A_�@�"@
�ٿ>�?�:l�@�j>nx	4@RD%��!?MC�A_�@O�.�ٿ=�Vy'|�@�?��v�3@�"���!?��o��@O�.�ٿ=�Vy'|�@�?��v�3@�"���!?��o��@?j`�ٿr��1�W�@�����3@0#�bh�!?z'�<_�@?j`�ٿr��1�W�@�����3@0#�bh�!?z'�<_�@?j`�ٿr��1�W�@�����3@0#�bh�!?z'�<_�@?j`�ٿr��1�W�@�����3@0#�bh�!?z'�<_�@?j`�ٿr��1�W�@�����3@0#�bh�!?z'�<_�@������ٿ�7]�En�@�ƙ�L�3@�H�g��!?).�塵@�Ŷ���ٿ����w�@�:~3�3@:k����!?*�ҋG�@�Ŷ���ٿ����w�@�:~3�3@:k����!?*�ҋG�@T��ٿ�Q�,�{�@�wH�6�3@�r�!?2V!Ϗ4�@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@�X���ٿ[�v��y�@��9B�3@���yl�!?E�I�g��@.T�@�ٿ�Ș���@�����3@.��sS�!?|�AT��@.T�@�ٿ�Ș���@�����3@.��sS�!?|�AT��@.T�@�ٿ�Ș���@�����3@.��sS�!?|�AT��@.T�@�ٿ�Ș���@�����3@.��sS�!?|�AT��@.T�@�ٿ�Ș���@�����3@.��sS�!?|�AT��@~RAŞٿ�H�;�4�@�Ì�4@P�])n�!?��"xf�@���K{�ٿ�����-�@4Hm4@��-X�!?cse�zд@���K{�ٿ�����-�@4Hm4@��-X�!?cse�zд@��Y�ٿ8#� ��@���7�4@�[t��!?M�����@��Y�ٿ8#� ��@���7�4@�[t��!?M�����@ڠ;;סٿ	�mJ���@� �l��3@^aÙ�!?��n��@ڠ;;סٿ	�mJ���@� �l��3@^aÙ�!?��n��@ڠ;;סٿ	�mJ���@� �l��3@^aÙ�!?��n��@ڠ;;סٿ	�mJ���@� �l��3@^aÙ�!?��n��@ڠ;;סٿ	�mJ���@� �l��3@^aÙ�!?��n��@����,�ٿ�R�0�@�J±��3@�I�#�!?�I�*�/�@�7e�q�ٿ�)�sw/�@�r�x�4@KK�+�!?jl���Ŵ@�7e�q�ٿ�)�sw/�@�r�x�4@KK�+�!?jl���Ŵ@���I{�ٿ��չ�@��4,��3@jV�5�!?���_{�@���I{�ٿ��չ�@��4,��3@jV�5�!?���_{�@���I{�ٿ��չ�@��4,��3@jV�5�!?���_{�@���I{�ٿ��չ�@��4,��3@jV�5�!?���_{�@���I{�ٿ��չ�@��4,��3@jV�5�!?���_{�@
�B�N�ٿ�>� �@E��M�4@����U�!?���LU�@
�B�N�ٿ�>� �@E��M�4@����U�!?���LU�@��N�ٿ�TDv��@�=WM�	4@:�WM�!?O�Z�j	�@��N�ٿ�TDv��@�=WM�	4@:�WM�!?O�Z�j	�@��N�ٿ�TDv��@�=WM�	4@:�WM�!?O�Z�j	�@�٨K+�ٿ�4Dt4�@�eB+4@��*P��!?Zj\�>��@~u�+2�ٿ�g�Г�@s�e�5�3@�4?�!?��L�ĵ@�\���ٿpqKM��@6�gRV4@1���Ǐ!?� �"�@�\���ٿpqKM��@6�gRV4@1���Ǐ!?� �"�@1 �}�ٿ�*�-D��@l�^��3@j��뢐!?:��	'�@1 �}�ٿ�*�-D��@l�^��3@j��뢐!?:��	'�@1 �}�ٿ�*�-D��@l�^��3@j��뢐!?:��	'�@��V �ٿ��6A�@������3@+�}]�!?���f�@��V �ٿ��6A�@������3@+�}]�!?���f�@��V �ٿ��6A�@������3@+�}]�!?���f�@��V �ٿ��6A�@������3@+�}]�!?���f�@�
記ٿ��g���@tx�t�3@��3�g�!?3ʣ��@�
記ٿ��g���@tx�t�3@��3�g�!?3ʣ��@�
記ٿ��g���@tx�t�3@��3�g�!?3ʣ��@�
記ٿ��g���@tx�t�3@��3�g�!?3ʣ��@gF�
H�ٿk����@R�4�3@���F�!?���b��@gF�
H�ٿk����@R�4�3@���F�!?���b��@h#Gܙٿ�t�_�d�@�աT�3@�)��i�!?�i �@h#Gܙٿ�t�_�d�@�աT�3@�)��i�!?�i �@h#Gܙٿ�t�_�d�@�աT�3@�)��i�!?�i �@�\W�n�ٿ?>7��@��W�3@~y+|�!?;�=P���@�\W�n�ٿ?>7��@��W�3@~y+|�!?;�=P���@�\W�n�ٿ?>7��@��W�3@~y+|�!?;�=P���@�\W�n�ٿ?>7��@��W�3@~y+|�!?;�=P���@݉4��ٿj������@e��� 4@p�)�J�!?�آ��@���H��ٿ�^�'�+�@�C���3@X��~�!?�3� g�@���H��ٿ�^�'�+�@�C���3@X��~�!?�3� g�@���H��ٿ�^�'�+�@�C���3@X��~�!?�3� g�@���H��ٿ�^�'�+�@�C���3@X��~�!?�3� g�@���H��ٿ�^�'�+�@�C���3@X��~�!?�3� g�@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@oQ(�ٿ�Ԩ'��@�p���4@�4m�l�!?����@�p�i��ٿ�E`�:��@���h4@B(%��!?�%%����@�p�i��ٿ�E`�:��@���h4@B(%��!?�%%����@�p�i��ٿ�E`�:��@���h4@B(%��!?�%%����@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@-ឝ��ٿ��M��@t=A��3@�&/�!?�� �ߵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@���f�ٿ��A��U�@��.�3@�2"=�!?��Q�ĵ@~��q��ٿӗ���@0~B�3@}�b��!?��ߙ]�@��Ԑ�ٿ�[(ws��@���3@��!?���֝{�@��Ԑ�ٿ�[(ws��@���3@��!?���֝{�@��Ԑ�ٿ�[(ws��@���3@��!?���֝{�@��Ԑ�ٿ�[(ws��@���3@��!?���֝{�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@���\~�ٿ*e���@�7Q�d�3@���騐!?f����4�@N��h7�ٿ5M\�@�"K��4@�ϐ�!?�J���@N��h7�ٿ5M\�@�"K��4@�ϐ�!?�J���@N��h7�ٿ5M\�@�"K��4@�ϐ�!?�J���@N��h7�ٿ5M\�@�"K��4@�ϐ�!?�J���@�\��0�ٿ��:eC��@@G�i�3@�0@�j�!?K���@�\��0�ٿ��:eC��@@G�i�3@�0@�j�!?K���@�\��0�ٿ��:eC��@@G�i�3@�0@�j�!?K���@�\��0�ٿ��:eC��@@G�i�3@�0@�j�!?K���@�\��0�ٿ��:eC��@@G�i�3@�0@�j�!?K���@c�?@�ٿ�N<\Vz�@��� 4@�u53Đ!?�L~I��@�7�ᐚٿ9������@�;��3@b��*�!?E��gX�@����җٿӯwP={�@��<�3@\\�:�!?(m|DQ��@����җٿӯwP={�@��<�3@\\�:�!?(m|DQ��@����җٿӯwP={�@��<�3@\\�:�!?(m|DQ��@�oA0�ٿ0ə$f^�@�W���3@=�`�'�!?��}2�@�oA0�ٿ0ə$f^�@�W���3@=�`�'�!?��}2�@�oA0�ٿ0ə$f^�@�W���3@=�`�'�!?��}2�@�oA0�ٿ0ə$f^�@�W���3@=�`�'�!?��}2�@�oA0�ٿ0ə$f^�@�W���3@=�`�'�!?��}2�@���'�ٿ,w����@HB�R��3@��As�!?���É�@���'�ٿ,w����@HB�R��3@��As�!?���É�@���'�ٿ,w����@HB�R��3@��As�!?���É�@���'�ٿ,w����@HB�R��3@��As�!?���É�@���'�ٿ,w����@HB�R��3@��As�!?���É�@+R^���ٿ��4BI��@��(d��3@��w��!?TFa��8�@of�{C�ٿt��Y��@���� 4@-�*V�!?�H�S-i�@�E.?,�ٿ�|�mu`�@GL�f�3@�dLe�!?����@�E.?,�ٿ�|�mu`�@GL�f�3@�dLe�!?����@�	�.�ٿ�Z�Y�@�^�u�3@;���k�!?[�TH�@F,u�ٿ�k�:�8�@�(d:0�3@�-��,�!?���(�1�@F,u�ٿ�k�:�8�@�(d:0�3@�-��,�!?���(�1�@F,u�ٿ�k�:�8�@�(d:0�3@�-��,�!?���(�1�@���ϒٿQ-D@���@yO�U��3@��V�3�!?A���d��@���ϒٿQ-D@���@yO�U��3@��V�3�!?A���d��@���ϒٿQ-D@���@yO�U��3@��V�3�!?A���d��@���ϒٿQ-D@���@yO�U��3@��V�3�!?A���d��@xw���ٿ����v�@nK���3@p�5��!?|;��ә�@xw���ٿ����v�@nK���3@p�5��!?|;��ә�@xw���ٿ����v�@nK���3@p�5��!?|;��ә�@xw���ٿ����v�@nK���3@p�5��!?|;��ә�@xw���ٿ����v�@nK���3@p�5��!?|;��ә�@%O�䭙ٿ���)�b�@-��4@*�E�!?�o�h�@%O�䭙ٿ���)�b�@-��4@*�E�!?�o�h�@%�J�@�ٿ�̳��@���4@�Z�!?�I��:�@%�J�@�ٿ�̳��@���4@�Z�!?�I��:�@%�J�@�ٿ�̳��@���4@�Z�!?�I��:�@>MD���ٿr�@_)�@���m�4@n.ͮ+�!?�l
�0�@>MD���ٿr�@_)�@���m�4@n.ͮ+�!?�l
�0�@>MD���ٿr�@_)�@���m�4@n.ͮ+�!?�l
�0�@��l��ٿ�r1���@���@4@4�Q�K�!?�pS�U�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@��x���ٿh,n���@ڴ��@�3@��G��!?�y|B&;�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�T-��ٿ7�R���@����3@��L�P�!?�F���j�@�r�!�ٿ��*/��@B̝��3@Jŏ,�!?PͲO�+�@���P��ٿ�ؓ��@+i���3@nE�xۏ!?K����@���P��ٿ�ؓ��@+i���3@nE�xۏ!?K����@���P��ٿ�ؓ��@+i���3@nE�xۏ!?K����@�Ǟ;*�ٿ��on#�@���:H�3@���X�!?���'���@�Ǟ;*�ٿ��on#�@���:H�3@���X�!?���'���@��D���ٿ������@/g��3@��:4�!?[�µ@��D���ٿ������@/g��3@��:4�!?[�µ@�x��G�ٿ�� ��@�i���3@��aCL�!?@��L7�@�x��G�ٿ�� ��@�i���3@��aCL�!?@��L7�@�x��G�ٿ�� ��@�i���3@��aCL�!?@��L7�@�x��G�ٿ�� ��@�i���3@��aCL�!?@��L7�@�|`�u�ٿ��Y�a�@����}�3@�����!?D���Ƞ�@�|`�u�ٿ��Y�a�@����}�3@�����!?D���Ƞ�@�|`�u�ٿ��Y�a�@����}�3@�����!?D���Ƞ�@8�[��ٿC�4�(~�@C�?��3@ ����!?0� ��@8�[��ٿC�4�(~�@C�?��3@ ����!?0� ��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@���ƍٿ�"���@���}��3@���D�!?R�.��@�Г�-�ٿO1jA��@[ӟm�3@x�p.�!?ԖE�~�@�Г�-�ٿO1jA��@[ӟm�3@x�p.�!?ԖE�~�@�Г�-�ٿO1jA��@[ӟm�3@x�p.�!?ԖE�~�@�So�8�ٿ�2���@׮&�/�3@|��#�!?+!$Vk�@�So�8�ٿ�2���@׮&�/�3@|��#�!?+!$Vk�@�So�8�ٿ�2���@׮&�/�3@|��#�!?+!$Vk�@��H=�ٿs�M |��@{�p�3@�`��3�!?��&U���@��H=�ٿs�M |��@{�p�3@�`��3�!?��&U���@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@C��	Y�ٿ��q�~U�@dv�2��3@P�Si�!?�5B}\�@g��э�ٿD��Xd�@�9>�#�3@	���u�!?�Z����@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@��L���ٿ�?˧��@"�:�3@���p�!?-Ѝ/��@�$LǛٿ��B8���@z5�\;�3@@rϡ��!?K�T�@S�@�$LǛٿ��B8���@z5�\;�3@@rϡ��!?K�T�@S�@�$LǛٿ��B8���@z5�\;�3@@rϡ��!?K�T�@S�@�$LǛٿ��B8���@z5�\;�3@@rϡ��!?K�T�@S�@�$LǛٿ��B8���@z5�\;�3@@rϡ��!?K�T�@S�@�F�)�ٿHUY~M��@���D 4@���e�!?j���@�F�)�ٿHUY~M��@���D 4@���e�!?j���@�F�)�ٿHUY~M��@���D 4@���e�!?j���@R�H��ٿ�zG��@�_�d�4@�%U�!?��H��@R�H��ٿ�zG��@�_�d�4@�%U�!?��H��@R�H��ٿ�zG��@�_�d�4@�%U�!?��H��@R�H��ٿ�zG��@�_�d�4@�%U�!?��H��@R�H��ٿ�zG��@�_�d�4@�%U�!?��H��@��~�ٿ�$�;�,�@8E��V�3@�OX�e�!?�����:�@��~�ٿ�$�;�,�@8E��V�3@�OX�e�!?�����:�@��~�ٿ�$�;�,�@8E��V�3@�OX�e�!?�����:�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@�l�<1�ٿ�b��JQ�@>*�:��3@�H(s��!?-�1o�;�@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@v֥�ٿ���V�@��OzM4@�s�4�!?�9�����@���o�ٿ��z����@
��4"�3@q�8t�!?��fXM�@���o�ٿ��z����@
��4"�3@q�8t�!?��fXM�@V�~�ٿ$]��jo�@�A����3@��ʾD�!?����/�@��F��ٿ�)�ɷ�@�m�J�4@H�"R��!?ܤ�����@�0�#ԕٿuɡe��@�Φ84@s �5{�!?�T��&�@�0�#ԕٿuɡe��@�Φ84@s �5{�!?�T��&�@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�6c�ٿ��!��@-a�Oe�3@�͝��!?WO�Ց��@�&�ٿ��<5�<�@�;����3@����z�!?�-eY��@[�ÇёٿQ��.��@A5���3@�*p��!?hL@kŵ@[�ÇёٿQ��.��@A5���3@�*p��!?hL@kŵ@[�ÇёٿQ��.��@A5���3@�*p��!?hL@kŵ@[�ÇёٿQ��.��@A5���3@�*p��!?hL@kŵ@[�ÇёٿQ��.��@A5���3@�*p��!?hL@kŵ@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@��D`�ٿ1������@��[%r�3@{O* �!?$�����@aC����ٿ[�2Ln�@�!�!�3@��oҏ!?� �]��@aC����ٿ[�2Ln�@�!�!�3@��oҏ!?� �]��@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@A�@#�ٿ�vi�"��@������3@䧮b�!?9���N�@�[��ٿ� SO"�@bڅV��3@,��`��!?]�C�͇�@�[��ٿ� SO"�@bڅV��3@,��`��!?]�C�͇�@�[��ٿ� SO"�@bڅV��3@,��`��!?]�C�͇�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@�����ٿqN���B�@�%!8��3@����|�!?�z�t�(�@��T�ٿiP�=�@�Rٷ4@�$� ��!?�ʠ(���@��T�ٿiP�=�@�Rٷ4@�$� ��!?�ʠ(���@��T�ٿiP�=�@�Rٷ4@�$� ��!?�ʠ(���@�8فH�ٿ;CZ���@�^�4�4@��w|�!?���( w�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@�!�>�ٿ��C�9�@�xE��3@�Y-Vt�!?Jh��b�@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@¢�K�ٿc��}��@ڐ|y�3@�J�D�!?V}��;��@e���ٿ��w�%�@:VK���3@��C� �!?,v*����@e���ٿ��w�%�@:VK���3@��C� �!?,v*����@e���ٿ��w�%�@:VK���3@��C� �!?,v*����@�6$p�ٿGfk$��@�X����3@����<�!?8��Y<2�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@st�o8�ٿry�����@��os�3@�^�_�!?	i���+�@��I/�ٿ��I��o�@�y�-�4@�;m���!?>r�X[��@��I/�ٿ��I��o�@�y�-�4@�;m���!?>r�X[��@i7-��ٿ��e4&�@
U��0�3@2SQ��!?ր���@i7-��ٿ��e4&�@
U��0�3@2SQ��!?ր���@�;:��ٿ�oc��@x���D�3@�2���!?4ю���@�;:��ٿ�oc��@x���D�3@�2���!?4ю���@�;:��ٿ�oc��@x���D�3@�2���!?4ю���@�;:��ٿ�oc��@x���D�3@�2���!?4ю���@�;:��ٿ�oc��@x���D�3@�2���!?4ю���@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@�y�v�ٿ��U�4��@(X���3@�s�b�!?���iSv�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@��T*Z�ٿ��=�q*�@Aӣ��3@1��3.�!?jA�@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@e��<�ٿ����N�@X7�2�3@�=.*�!?V��׵@嵢�ϐٿ\|2�2��@k���Z�3@��Is�!?V��ܵ@�iX�ٿ?�w��@���^�3@h�>rd�!?�N�;*�@(˄\e�ٿ�����L�@�4��3@�O�)l�!?�A�)p~�@(˄\e�ٿ�����L�@�4��3@�O�)l�!?�A�)p~�@���W�ٿ(��b�@�=�g�3@>�%��!?E�&�]�@���W�ٿ(��b�@�=�g�3@>�%��!?E�&�]�@���W�ٿ(��b�@�=�g�3@>�%��!?E�&�]�@O��ӕٿ�.+ms�@R�k�3@��ׯ�!?����E�@O��ӕٿ�.+ms�@R�k�3@��ׯ�!?����E�@O��ӕٿ�.+ms�@R�k�3@��ׯ�!?����E�@O��ӕٿ�.+ms�@R�k�3@��ׯ�!?����E�@Ϝ�}�ٿ�m���@_X�L:�3@f��x�!?�RT����@Ϝ�}�ٿ�m���@_X�L:�3@f��x�!?�RT����@��X�u�ٿ��-<�@���L��3@t5|���!?��"Z}̵@��X�u�ٿ��-<�@���L��3@t5|���!?��"Z}̵@��X�u�ٿ��-<�@���L��3@t5|���!?��"Z}̵@��X�u�ٿ��-<�@���L��3@t5|���!?��"Z}̵@��X�u�ٿ��-<�@���L��3@t5|���!?��"Z}̵@����ڕٿF
@�;��@�Vk�3@y%s���!?�zX�"õ@����ڕٿF
@�;��@�Vk�3@y%s���!?�zX�"õ@!S'8��ٿiz�ڧ��@y{qT��3@�LGʐ!?F��;���@]�~)�ٿx����@�����3@��q�ؐ!?�aEq��@]�~)�ٿx����@�����3@��q�ؐ!?�aEq��@f��'F�ٿѷ����@33,Օ�3@�i�?�!?��2�Xδ@f��'F�ٿѷ����@33,Օ�3@�i�?�!?��2�Xδ@f��'F�ٿѷ����@33,Օ�3@�i�?�!?��2�Xδ@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@ʾ��h�ٿEƄ+�m�@��l��3@��s�!?R�Gl1�@��'52�ٿ�2Us���@��q�.�3@d�D=_�!?dۇ���@��'52�ٿ�2Us���@��q�.�3@d�D=_�!?dۇ���@Ȫw�o�ٿ c~f�@-,��3@b��I,�!?G��� �@Ȫw�o�ٿ c~f�@-,��3@b��I,�!?G��� �@Ȫw�o�ٿ c~f�@-,��3@b��I,�!?G��� �@Ȫw�o�ٿ c~f�@-,��3@b��I,�!?G��� �@Ȫw�o�ٿ c~f�@-,��3@b��I,�!?G��� �@P�[�X�ٿn�q(��@_��pS�3@ɻ\D�!?��ָ���@P�[�X�ٿn�q(��@_��pS�3@ɻ\D�!?��ָ���@P�[�X�ٿn�q(��@_��pS�3@ɻ\D�!?��ָ���@L���ۗٿ�����@�cs4@f�D-�!?�TI
ӵ@�Rx[�ٿve�b��@��}��3@����+�!?�WX���@�Rx[�ٿve�b��@��}��3@����+�!?�WX���@�Rx[�ٿve�b��@��}��3@����+�!?�WX���@P4
z�ٿ�D�Y�^�@�vk���3@��E�!?�K�-9�@P4
z�ٿ�D�Y�^�@�vk���3@��E�!?�K�-9�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@C$���ٿ��QX
�@;-F���3@D��N��!?q��� "�@E�Qv��ٿ��+���@/�ynn�3@!�I�!?��+��)�@E�Qv��ٿ��+���@/�ynn�3@!�I�!?��+��)�@E�Qv��ٿ��+���@/�ynn�3@!�I�!?��+��)�@E�Qv��ٿ��+���@/�ynn�3@!�I�!?��+��)�@E�Qv��ٿ��+���@/�ynn�3@!�I�!?��+��)�@}���ٿl�~���@U$�3@q�!�_�!?�h .&�@��WBd�ٿ&g}p[��@P6[��3@���.��!?���ꮉ�@��WBd�ٿ&g}p[��@P6[��3@���.��!?���ꮉ�@��WBd�ٿ&g}p[��@P6[��3@���.��!?���ꮉ�@��WBd�ٿ&g}p[��@P6[��3@���.��!?���ꮉ�@��WBd�ٿ&g}p[��@P6[��3@���.��!?���ꮉ�@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@��Lc�ٿ�ٷ�i��@;�$�4@!�_�S�!?i �G��@(⎴�ٿZ �����@Y��ދ4@�m��!?Q�pPl�@>]*)��ٿS�3����@z�-�4@G�ar��!?����b�@{�'��ٿ�u���@��ّ��3@k�����!?�D���@{�'��ٿ�u���@��ّ��3@k�����!?�D���@{�'��ٿ�u���@��ّ��3@k�����!?�D���@{�'��ٿ�u���@��ّ��3@k�����!?�D���@����ٿWD%��@���J_�3@���B�!?�R~��@����ٿWD%��@���J_�3@���B�!?�R~��@����ٿWD%��@���J_�3@���B�!?�R~��@����ٿWD%��@���J_�3@���B�!?�R~��@����ٿWD%��@���J_�3@���B�!?�R~��@�NX��ٿ']QW���@"�W���3@9���)�!?M�����@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@i>'�ݞٿ�.Ҁ��@\]	Mf�3@��E�M�!?\B�r�@��-A{�ٿ�e�AY�@����3@���U�!?mt�|8�@��-A{�ٿ�e�AY�@����3@���U�!?mt�|8�@��-A{�ٿ�e�AY�@����3@���U�!?mt�|8�@1QY���ٿG��Τ�@l}k�3@�)�u�!?sp��@1QY���ٿG��Τ�@l}k�3@�)�u�!?sp��@1QY���ٿG��Τ�@l}k�3@�)�u�!?sp��@1QY���ٿG��Τ�@l}k�3@�)�u�!?sp��@�M��/�ٿ��ǯv�@�����3@=���Y�!?$i4,��@�M��/�ٿ��ǯv�@�����3@=���Y�!?$i4,��@�M��/�ٿ��ǯv�@�����3@=���Y�!?$i4,��@�M��/�ٿ��ǯv�@�����3@=���Y�!?$i4,��@��0�j�ٿY�G3���@��V�3@�2���!?Ť���R�@��5�ٿ�����@��^�*�3@4�u0�!?^������@��5�ٿ�����@��^�*�3@4�u0�!?^������@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@z0�h̔ٿ��]��@ .4���3@�S\q/�!?���|�@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@l��\^�ٿS�.��[�@hb9,��3@�/�u_�!?}�rO��@	�Oˏ�ٿ�#�U�@B����3@i�ג��!?3�E$Q�@	�Oˏ�ٿ�#�U�@B����3@i�ג��!?3�E$Q�@	�Oˏ�ٿ�#�U�@B����3@i�ג��!?3�E$Q�@	�Oˏ�ٿ�#�U�@B����3@i�ג��!?3�E$Q�@	�Oˏ�ٿ�#�U�@B����3@i�ג��!?3�E$Q�@8�r�ٿ��z6�z�@=����3@u}���!?��i���@8�r�ٿ��z6�z�@=����3@u}���!?��i���@8�r�ٿ��z6�z�@=����3@u}���!?��i���@8�r�ٿ��z6�z�@=����3@u}���!?��i���@�R�G��ٿ}�g@8�@9D���3@����!?����rB�@���W��ٿA.��w�@\K*ؘ�3@���ӏ!?�s3G�@���W��ٿA.��w�@\K*ؘ�3@���ӏ!?�s3G�@����ٿ*]�~z��@s�3yS�3@��ycӏ!?��C��@����ٿ���E��@qAJ1��3@����<�!?�'��@����ٿ���E��@qAJ1��3@����<�!?�'��@9q?�Ïٿ,��AE��@�Y^�4@��5}~�!?���6�@9q?�Ïٿ,��AE��@�Y^�4@��5}~�!?���6�@8P���ٿh��x���@GA�Z��3@�f����!?U���M�@8P���ٿh��x���@GA�Z��3@�f����!?U���M�@8P���ٿh��x���@GA�Z��3@�f����!?U���M�@9n���ٿĥ�E7f�@4^��|�3@lAx�!?�h�G�1�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@�#�ٿG�Iͷ�@��EH��3@F�A�p�!?H�t�03�@	n�Ôٿd�jP�@㣒���3@ޱ!'��!?�_�"r��@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@�=)=�ٿ��?���@����8�3@2�F�!?��=H7�@XM㹗ٿ9�3(V��@;$�3@���Q\�!?M<ݖCn�@�b?l��ٿ��{���@�|F���3@�.��
�!?w_�%���@�b?l��ٿ��{���@�|F���3@�.��
�!?w_�%���@�b?l��ٿ��{���@�|F���3@�.��
�!?w_�%���@�b?l��ٿ��{���@�|F���3@�.��
�!?w_�%���@�b?l��ٿ��{���@�|F���3@�.��
�!?w_�%���@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@�E�ɛٿ���v���@t�η��3@�ʺF�!?
\����@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@$p(ꓑٿc�7����@-r�e�3@�J�:�!?C#��<�@��x'F�ٿ�/}�2�@+*h[�4@�Y�X�!?!�$c��@1_^��ٿ
�-1��@ �����3@,�k�!?PZ()�ڴ@1_^��ٿ
�-1��@ �����3@,�k�!?PZ()�ڴ@1_^��ٿ
�-1��@ �����3@,�k�!?PZ()�ڴ@1_^��ٿ
�-1��@ �����3@,�k�!?PZ()�ڴ@1_^��ٿ
�-1��@ �����3@,�k�!?PZ()�ڴ@� �U��ٿm쿹�$�@I�0���3@��K��!?A�#��w�@� �U��ٿm쿹�$�@I�0���3@��K��!?A�#��w�@����ٿ����l��@��j��3@��I�!?�Z�E0��@����ٿ����l��@��j��3@��I�!?�Z�E0��@����ٿ����l��@��j��3@��I�!?�Z�E0��@����ٿ����l��@��j��3@��I�!?�Z�E0��@����ٿ����l��@��j��3@��I�!?�Z�E0��@�5���ٿ���2�@�L�<�4@����	�!?Dŭj�ϴ@�5���ٿ���2�@�L�<�4@����	�!?Dŭj�ϴ@�5���ٿ���2�@�L�<�4@����	�!?Dŭj�ϴ@�ӄ.9�ٿ�gZM�w�@��+�34@�����!?8�}Y&��@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@{�&�+�ٿ6\�@��@$�I�/4@����1�!?�U�0�@/&�� �ٿ�N�?�@��g%�4@�D,�Z�!?.��Q��@/&�� �ٿ�N�?�@��g%�4@�D,�Z�!?.��Q��@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@)7|'�ٿE��`���@��$���3@2�?�!?�-�gF�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@߇���ٿ��.�;��@In��`�3@�\Ni�!?b0.P$)�@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@V�7	�ٿ[��~'�@Eaj��3@E��_��!?�z�8��@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@LЕ$�ٿ�Hl�u�@��1��3@E�f�b�!?�w�o�@��_�ٿ�yK%��@b?����3@������!?����L�@��_�ٿ�yK%��@b?����3@������!?����L�@��_�ٿ�yK%��@b?����3@������!?����L�@��_�ٿ�yK%��@b?����3@������!?����L�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@��п�ٿ�d�Ecp�@ �W�1�3@�\�u�!?���#�8�@����ٿ���ŭW�@ڶn��3@��u<��!?������@����ٿ���ŭW�@ڶn��3@��u<��!?������@����ٿ���ŭW�@ڶn��3@��u<��!?������@����ٿ���ŭW�@ڶn��3@��u<��!?������@]6Ke�ٿ)��9���@������3@�O�ŏ�!?R�Q��@]6Ke�ٿ)��9���@������3@�O�ŏ�!?R�Q��@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@<Z 0�ٿ���P>��@ʹ���3@2�Q���!?���`|�@�1��ٿ�@��,�@�+
���3@&���!?�?8b��@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@x<�A��ٿBţ����@ y����3@�
hݼ�!?-,ml8�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@����ٿ�vdv���@|X���3@jb�ס�!?���-b�@���]�ٿS��3!��@��C��3@L�*M.�!?�^�����@���]�ٿS��3!��@��C��3@L�*M.�!?�^�����@���]�ٿS��3!��@��C��3@L�*M.�!?�^�����@���]�ٿS��3!��@��C��3@L�*M.�!?�^�����@���]�ٿS��3!��@��C��3@L�*M.�!?�^�����@�iO���ٿއo�G�@������3@w/-]��!?{2{�1�@�iO���ٿއo�G�@������3@w/-]��!?{2{�1�@�
�\�ٿ%F�xƿ@{�D�3@��x��!?��(�{�@�-�Ŕٿ��5A,
�@D/q��3@ѝYѾ�!?�g���ݴ@:�N��ٿ���|�f�@�6��%�3@��5ɐ!?��ә��@:�N��ٿ���|�f�@�6��%�3@��5ɐ!?��ә��@:�N��ٿ���|�f�@�6��%�3@��5ɐ!?��ә��@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@ʀt�ǜٿ���(�J�@'Z���3@RD8�U�!?H�� �@����ٿxy����@�v���3@{�]�!?|P[%���@����ٿxy����@�v���3@{�]�!?|P[%���@����ٿxy����@�v���3@{�]�!?|P[%���@{�$�ٿv�N ���@`,U�-�3@���vx�!?^:�7�?�@{�$�ٿv�N ���@`,U�-�3@���vx�!?^:�7�?�@{�$�ٿv�N ���@`,U�-�3@���vx�!?^:�7�?�@{�$�ٿv�N ���@`,U�-�3@���vx�!?^:�7�?�@%�G�ٿq�hG�@0N"j44@��?c�!?�;d�?��@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�ë=�ٿY�z�@ۖή+4@�8�!?���u�F�@�+�d��ٿ���%���@<�sS�4@�)�i�!?{Z���@�+�d��ٿ���%���@<�sS�4@�)�i�!?{Z���@�+�d��ٿ���%���@<�sS�4@�)�i�!?{Z���@�+�d��ٿ���%���@<�sS�4@�)�i�!?{Z���@�+�d��ٿ���%���@<�sS�4@�)�i�!?{Z���@�'��j�ٿ3�J��@M$`�4@��Ł�!?뭓�R��@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@,�oݖ�ٿ�G�@�x�T��3@�nzh�!?��~WC�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@W����ٿV�[�+��@H��JP�3@��H:�!?-��i�@����ٿݩ�i���@����3@������!?�%��Ŵ@����ٿݩ�i���@����3@������!?�%��Ŵ@� �D�ٿ�`\ݡ�@��M��3@.���i�!?.&>�瘵@� �D�ٿ�`\ݡ�@��M��3@.���i�!?.&>�瘵@� �D�ٿ�`\ݡ�@��M��3@.���i�!?.&>�瘵@� �D�ٿ�`\ݡ�@��M��3@.���i�!?.&>�瘵@� �D�ٿ�`\ݡ�@��M��3@.���i�!?.&>�瘵@��_3��ٿٲ�@2��@��hy7�3@x�.��!?�x&2��@��_3��ٿٲ�@2��@��hy7�3@x�.��!?�x&2��@��_3��ٿٲ�@2��@��hy7�3@x�.��!?�x&2��@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@��i6ڜٿrXF*q�@�XAQ+�3@��R(S�!?�H�Ҵ@hf(��ٿ�c��N�@�s(��3@���I��!?d�P�(��@hf(��ٿ�c��N�@�s(��3@���I��!?d�P�(��@hf(��ٿ�c��N�@�s(��3@���I��!?d�P�(��@hf(��ٿ�c��N�@�s(��3@���I��!?d�P�(��@�.��t�ٿ���Y�@��%\�3@�o�z@�!?�a]4<�@�.��t�ٿ���Y�@��%\�3@�o�z@�!?�a]4<�@#��
N�ٿ�;L9�]�@ʈ���3@`��Ə!?��M��Y�@#��
N�ٿ�;L9�]�@ʈ���3@`��Ə!?��M��Y�@#��
N�ٿ�;L9�]�@ʈ���3@`��Ə!?��M��Y�@#��
N�ٿ�;L9�]�@ʈ���3@`��Ə!?��M��Y�@#��
N�ٿ�;L9�]�@ʈ���3@`��Ə!?��M��Y�@����5�ٿ�����m�@?�1Sb�3@�d^H-�!?�����@����5�ٿ�����m�@?�1Sb�3@�d^H-�!?�����@����5�ٿ�����m�@?�1Sb�3@�d^H-�!?�����@����5�ٿ�����m�@?�1Sb�3@�d^H-�!?�����@����5�ٿ�����m�@?�1Sb�3@�d^H-�!?�����@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@���g��ٿ*b�)�@�&
v�3@�H�-�!?���Ӵ@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ſY4�ٿnm��@��D�3@�y&dc�!?�	^U���@ꢸB�ٿjJu�/��@�4d���3@�Gz�B�!?o|��-�@ꢸB�ٿjJu�/��@�4d���3@�Gz�B�!?o|��-�@ꢸB�ٿjJu�/��@�4d���3@�Gz�B�!?o|��-�@ꢸB�ٿjJu�/��@�4d���3@�Gz�B�!?o|��-�@ꢸB�ٿjJu�/��@�4d���3@�Gz�B�!?o|��-�@ �%Xk�ٿ3�{"�e�@��U��3@ �1�5�!?�r6c7�@ �%Xk�ٿ3�{"�e�@��U��3@ �1�5�!?�r6c7�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@P �z{�ٿ�7�M��@�ғ��4@�y�h�!?��(x4�@��e(�ٿ	���t��@��s#<�3@�^!?�!�-m��@��e(�ٿ	���t��@��s#<�3@�^!?�!�-m��@�	*OB�ٿ<ձ,��@X��_X�3@�d�)O�!?��q��ȴ@�	*OB�ٿ<ձ,��@X��_X�3@�d�)O�!?��q��ȴ@�	*OB�ٿ<ձ,��@X��_X�3@�d�)O�!?��q��ȴ@�	*OB�ٿ<ձ,��@X��_X�3@�d�)O�!?��q��ȴ@�	*OB�ٿ<ձ,��@X��_X�3@�d�)O�!?��q��ȴ@�����ٿ� ʿM�@���%�3@�$md�!?+3�_�@�����ٿ� ʿM�@���%�3@�$md�!?+3�_�@�����ٿ� ʿM�@���%�3@�$md�!?+3�_�@�����ٿ� ʿM�@���%�3@�$md�!?+3�_�@rV���ٿ�\L�Z��@;����3@�U��W�!?��Y���@rV���ٿ�\L�Z��@;����3@�U��W�!?��Y���@rV���ٿ�\L�Z��@;����3@�U��W�!?��Y���@�MO�I�ٿ8 ����@-�oł�3@��V0��!?��S���@�MO�I�ٿ8 ����@-�oł�3@��V0��!?��S���@�MO�I�ٿ8 ����@-�oł�3@��V0��!?��S���@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@7j��ٿ;'��Y��@4�C���3@��>���!?U��'7�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�w�ѕٿ�\O �@�1ʅ�3@ѥ�R��!?�x��6*�@�*.��ٿx���l��@%��BH�3@����{�!?��8�k�@�*.��ٿx���l��@%��BH�3@����{�!?��8�k�@�*.��ٿx���l��@%��BH�3@����{�!?��8�k�@�5�+�ٿ:@1���@��\<��3@<���f�!?	�D����@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@� ��
�ٿ#������@ŭf]� 4@{:W��!?����ɴ@�	3���ٿZ�+���@�z��\�3@m*�;�!?}c����@��6��ٿo���A�@��u�3@Y�k+b�!?Ǔ�p�ǵ@�!��ٿRs�p���@CX�I�3@(���V�!?;�����@�!��ٿRs�p���@CX�I�3@(���V�!?;�����@�!��ٿRs�p���@CX�I�3@(���V�!?;�����@~A����ٿ�Ka8n�@� m��3@��*�!?��|df�@~A����ٿ�Ka8n�@� m��3@��*�!?��|df�@v���;�ٿ�4�S4�@��ZI�3@�x!?����
�@v���;�ٿ�4�S4�@��ZI�3@�x!?����
�@v���;�ٿ�4�S4�@��ZI�3@�x!?����
�@v���;�ٿ�4�S4�@��ZI�3@�x!?����
�@���Z�ٿ�y~]g��@��T�3@z|�S�!?ze8����@���Z�ٿ�y~]g��@��T�3@z|�S�!?ze8����@CyS Ûٿ��=���@�����3@��J��!?�>�@CyS Ûٿ��=���@�����3@��J��!?�>�@CyS Ûٿ��=���@�����3@��J��!?�>�@O�����ٿ�4"-�)�@��tC�3@ ��!?��iQ��@O�����ٿ�4"-�)�@��tC�3@ ��!?��iQ��@O�����ٿ�4"-�)�@��tC�3@ ��!?��iQ��@,�ű�ٿ��Z����@�;p;��3@�ӑ*-�!?�A��¸�@�i� ��ٿNa��Dj�@!�5�3@��A�!?�i⎵@��x`R�ٿ���
���@[`�o��3@�눇�!?0P���]�@Gt�N	�ٿ��7���@�k��3@A�)h�!?�#ed��@Gt�N	�ٿ��7���@�k��3@A�)h�!?�#ed��@DV�Ͳ�ٿ�O���[�@��f(�4@~i�p�!?�Zӻd;�@���m�ٿ�^K ���@����4@HM�V��!?�RVC�@���m�ٿ�^K ���@����4@HM�V��!?�RVC�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��W���ٿ=ī����@����4@�7,K��!?�Qnyk�@��B��ٿ���@�R��Q4@�	��z�!?ԄU)�մ@��B��ٿ���@�R��Q4@�	��z�!?ԄU)�մ@��B��ٿ���@�R��Q4@�	��z�!?ԄU)�մ@%��p�ٿ����O�@�+���4@�ߌYC�!?�N	�P^�@8:yl�ٿ8���wI�@d��<�4@6+HDH�!?ޕ����@8:yl�ٿ8���wI�@d��<�4@6+HDH�!?ޕ����@8:yl�ٿ8���wI�@d��<�4@6+HDH�!?ޕ����@7?��V�ٿrW��g�@S9`��4@��rC��!?͠�yF�@7?��V�ٿrW��g�@S9`��4@��rC��!?͠�yF�@���L�ٿ���0x��@�e���4@��A���!?������@���L�ٿ���0x��@�e���4@��A���!?������@����U�ٿ?��/mE�@F��D4@1:����!?2$L�@5�8���ٿ��9dM��@�=�E;4@au�2
�!?�b��δ@5�8���ٿ��9dM��@�=�E;4@au�2
�!?�b��δ@5�8���ٿ��9dM��@�=�E;4@au�2
�!?�b��δ@�2[��ٿ�u��a�@�47y�3@��$}�!?i1z���@�2[��ٿ�u��a�@�47y�3@��$}�!?i1z���@�2[��ٿ�u��a�@�47y�3@��$}�!?i1z���@�2[��ٿ�u��a�@�47y�3@��$}�!?i1z���@�2[��ٿ�u��a�@�47y�3@��$}�!?i1z���@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@�cNT�ٿ7Ɩ;(�@Y�w��4@�`��!?��Њ$K�@4܊tq�ٿ( Ā2�@�44@k��)V�!?�X�S�@4܊tq�ٿ( Ā2�@�44@k��)V�!?�X�S�@±L=��ٿ���AC�@h�<�4@�f|Z]�!?ǳ�{`�@±L=��ٿ���AC�@h�<�4@�f|Z]�!?ǳ�{`�@�\�1Зٿ�����@0B}r�4@#]pN�!?��@���@'��ǎ�ٿ=<�y`l�@�_ӟ��3@��IPz�!?ӓI�Z+�@'��ǎ�ٿ=<�y`l�@�_ӟ��3@��IPz�!?ӓI�Z+�@�L&�9�ٿ�=���@�k�	4@ �GJ�!?�]a
�@E,�彘ٿ#�b��@#��zX�3@���W�!?�{���˴@E,�彘ٿ#�b��@#��zX�3@���W�!?�{���˴@E,�彘ٿ#�b��@#��zX�3@���W�!?�{���˴@E,�彘ٿ#�b��@#��zX�3@���W�!?�{���˴@E,�彘ٿ#�b��@#��zX�3@���W�!?�{���˴@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@�ؤ
�ٿ'�����@#ij�
�3@&���z�!?�]���	�@ڭ�毚ٿ�}��-��@�jRvz4@Z��)�!?)6:��S�@�\�ٿ#�x�)4�@UX;v�3@�f��!?�8�y�@�\�ٿ#�x�)4�@UX;v�3@�f��!?�8�y�@�\�ٿ#�x�)4�@UX;v�3@�f��!?�8�y�@�\�ٿ#�x�)4�@UX;v�3@�f��!?�8�y�@�\�ٿ#�x�)4�@UX;v�3@�f��!?�8�y�@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@X��d�ٿ<r
�f�@ ����3@�h�^�!?������@C�+��ٿ���E\_�@M��a��3@LH��7�!?� �ҏ��@C�+��ٿ���E\_�@M��a��3@LH��7�!?� �ҏ��@C�+��ٿ���E\_�@M��a��3@LH��7�!?� �ҏ��@C�+��ٿ���E\_�@M��a��3@LH��7�!?� �ҏ��@C�+��ٿ���E\_�@M��a��3@LH��7�!?� �ҏ��@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@J�I�ٿt1�lp��@ jY��3@g���!?��]G���@Q�Jo#�ٿ
V�N_e�@���_��3@ԃ=
ُ!?Q�h��@�2�0s�ٿ�_�n�@�g��3@�)#�/�!?2΋Ҵ@�2�0s�ٿ�_�n�@�g��3@�)#�/�!?2΋Ҵ@�2�0s�ٿ�_�n�@�g��3@�)#�/�!?2΋Ҵ@�2�0s�ٿ�_�n�@�g��3@�)#�/�!?2΋Ҵ@�2�0s�ٿ�_�n�@�g��3@�)#�/�!?2΋Ҵ@A��)�ٿm�~۟��@]��:? 4@C#��]�!?w�ǎa��@A��)�ٿm�~۟��@]��:? 4@C#��]�!?w�ǎa��@A��)�ٿm�~۟��@]��:? 4@C#��]�!?w�ǎa��@A��)�ٿm�~۟��@]��:? 4@C#��]�!?w�ǎa��@��e睒ٿ�X�����@4��f�4@�=����!?��f4���@��e睒ٿ�X�����@4��f�4@�=����!?��f4���@e�D\%�ٿ!�v���@R�q�� 4@�v�98�!?���,(��@�j��ٿü��E��@]���4@��q-�!?���8E/�@�j��ٿü��E��@]���4@��q-�!?���8E/�@�j��ٿü��E��@]���4@��q-�!?���8E/�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@�9���ٿa�����@_T .�4@��원!?���\s$�@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@��KĞٿJ�����@��^��3@WIw�0�!?�8�~޴@Mt�<�ٿE�aY�(�@�ߟ��3@��8-N�!?�
��翴@Mt�<�ٿE�aY�(�@�ߟ��3@��8-N�!?�
��翴@�(SJ{�ٿ v���@I$G�<�3@�c����!?=�i�i�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@����o�ٿ0 ��@o�W|�3@F:�Gr�!?=�S�9"�@8v�'n�ٿlJ���@.�(J�3@s(h�!?�]��ȴ@8v�'n�ٿlJ���@.�(J�3@s(h�!?�]��ȴ@8v�'n�ٿlJ���@.�(J�3@s(h�!?�]��ȴ@8v�'n�ٿlJ���@.�(J�3@s(h�!?�]��ȴ@8v�'n�ٿlJ���@.�(J�3@s(h�!?�]��ȴ@`N-Hn�ٿ�qD�|��@29PY�3@9����!?�������@`N-Hn�ٿ�qD�|��@29PY�3@9����!?�������@`N-Hn�ٿ�qD�|��@29PY�3@9����!?�������@�y�W�ٿ��e��M�@�YC��3@ A\uD�!?B��u�Y�@�y�W�ٿ��e��M�@�YC��3@ A\uD�!?B��u�Y�@�y�W�ٿ��e��M�@�YC��3@ A\uD�!?B��u�Y�@�y�W�ٿ��e��M�@�YC��3@ A\uD�!?B��u�Y�@V����ٿ����c��@��A/�3@UU7�M�!?0���D�@���g�ٿS��`�@Y#ť��3@=*1bq�!?��jߊf�@���g�ٿS��`�@Y#ť��3@=*1bq�!?��jߊf�@���g�ٿS��`�@Y#ť��3@=*1bq�!?��jߊf�@���g�ٿS��`�@Y#ť��3@=*1bq�!?��jߊf�@���g�ٿS��`�@Y#ť��3@=*1bq�!?��jߊf�@�]�6�ٿF��.<X�@u!��z�3@��Zg�!?{�c�@�]�6�ٿF��.<X�@u!��z�3@��Zg�!?{�c�@�]�6�ٿF��.<X�@u!��z�3@��Zg�!?{�c�@�]�6�ٿF��.<X�@u!��z�3@��Zg�!?{�c�@�]�6�ٿF��.<X�@u!��z�3@��Zg�!?{�c�@#C�2#�ٿR�`�@�S�u�3@���D�!?�в���@#C�2#�ٿR�`�@�S�u�3@���D�!?�в���@#C�2#�ٿR�`�@�S�u�3@���D�!?�в���@#C�2#�ٿR�`�@�S�u�3@���D�!?�в���@#C�2#�ٿR�`�@�S�u�3@���D�!?�в���@��d�7�ٿ]Kܶ��@�߂���3@	�98�!?���~V�@��d�7�ٿ]Kܶ��@�߂���3@	�98�!?���~V�@��d�7�ٿ]Kܶ��@�߂���3@	�98�!?���~V�@��d�7�ٿ]Kܶ��@�߂���3@	�98�!?���~V�@���K �ٿ�qx��@�]��3@U��*\�!?��2��@���K �ٿ�qx��@�]��3@U��*\�!?��2��@���K �ٿ�qx��@�]��3@U��*\�!?��2��@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@�C�|F�ٿ.�����@[�g��3@�V��A�!?!X��櫵@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@'
'z��ٿ�c�o�z�@N.~n��3@���B�!?�	ش@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@V�)�ٿ*a��H�@�a�	��3@A��S��!?���oL��@JC����ٿ�&S���@WG⼜�3@���|j�!?��
X��@JC����ٿ�&S���@WG⼜�3@���|j�!?��
X��@JC����ٿ�&S���@WG⼜�3@���|j�!?��
X��@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@G?1ےٿJ6I��1�@�=�4�3@���$��!?��ݨ7x�@�����ٿQ�%ͻk�@ژ�RE�3@L���y�!?w������@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@=8��^�ٿ>�_��@E�[:��3@`UMW�!?��o8��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@���q�ٿXJ�҈S�@��wm��3@Ԃ[�o�!?h/-
��@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@�/�Κٿ��bk��@��^a�4@2;�e`�!?�/C0>�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@��?M�ٿٟ�3���@� �E&�3@�y�k�!?���c�I�@F-]Jٛٿ�9;g���@<��7��3@�^�m�!?���n��@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��Tl��ٿ:w����@�B��3@���4c�!?���oʹ@��B# �ٿ�7����@6&3|�3@w���!?�	ߍǴ@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@v�R�u�ٿڄ���0�@���3@��4��!?j�9�5E�@��	�ٿ�ɣX;��@�"DZ��3@�4�-�!?f���ҵ@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@�h�.2�ٿ\���wN�@�Pj�f�3@!���!?�%��;�@p�M��ٿTR��@I.l�3@�y�C_�!?��CIA �@p�M��ٿTR��@I.l�3@�y�C_�!?��CIA �@p�M��ٿTR��@I.l�3@�y�C_�!?��CIA �@^n@�4�ٿ]��d��@oZ����3@�s�c�!?'z���Ƶ@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�Zn�ٿ5�!���@K����3@�<�d�!?��gKo�@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@�� ���ٿq�p���@�L�5�3@|�7<g�!?{��<���@m���ٿ��I|�@�º^}�3@�P��!??ɤj���@m���ٿ��I|�@�º^}�3@�P��!??ɤj���@�$�іٿ] 3��@U.�?��3@~����!?�8p!��@�$�іٿ] 3��@U.�?��3@~����!?�8p!��@�$�іٿ] 3��@U.�?��3@~����!?�8p!��@@^uYݙٿ�9�|	�@zZ5�G�3@��ٷ�!?�]E�?��@@^uYݙٿ�9�|	�@zZ5�G�3@��ٷ�!?�]E�?��@�����ٿݙD�	��@sN�,�3@k��a�!?3�k���@�����ٿݙD�	��@sN�,�3@k��a�!?3�k���@�����ٿݙD�	��@sN�,�3@k��a�!?3�k���@��U�ٿ�Ii���@)�:���3@W�lb�!?D�  �j�@��U�ٿ�Ii���@)�:���3@W�lb�!?D�  �j�@��U�ٿ�Ii���@)�:���3@W�lb�!?D�  �j�@p��!�ٿ�9��x��@���k�3@oEX�!?6,�7��@>�F���ٿ����@wF�B�3@UB>Z�!?0�0m�
�@�ې��ٿ�Qr�
��@2�@P��3@xѷ�f�!?:g	-�z�@�ې��ٿ�Qr�
��@2�@P��3@xѷ�f�!?:g	-�z�@�ې��ٿ�Qr�
��@2�@P��3@xѷ�f�!?:g	-�z�@�ې��ٿ�Qr�
��@2�@P��3@xѷ�f�!?:g	-�z�@�ې��ٿ�Qr�
��@2�@P��3@xѷ�f�!?:g	-�z�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@:�ֵ��ٿ���jt'�@��bf:�3@�8�Zg�!?t72(�@�-�m�ٿ������@�b���3@��zq�!?5����ڴ@�-�m�ٿ������@�b���3@��zq�!?5����ڴ@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@7�c̕�ٿ�~�m��@���9�3@K��;[�!?W<�hkd�@��0�ٿ�xo[E��@�}��t�3@����B�!?7�/B�i�@��0�ٿ�xo[E��@�}��t�3@����B�!?7�/B�i�@��0�ٿ�xo[E��@�}��t�3@����B�!?7�/B�i�@��0�ٿ�xo[E��@�}��t�3@����B�!?7�/B�i�@��0�ٿ�xo[E��@�}��t�3@����B�!?7�/B�i�@�b��"�ٿ�`��g�@WIC��3@�c�X�!?���I|�@�b��"�ٿ�`��g�@WIC��3@�c�X�!?���I|�@�b��"�ٿ�`��g�@WIC��3@�c�X�!?���I|�@�b��"�ٿ�`��g�@WIC��3@�c�X�!?���I|�@�b��"�ٿ�`��g�@WIC��3@�c�X�!?���I|�@�z����ٿ�q�8���@���s�3@	�Ŀ��!?]w����@�z����ٿ�q�8���@���s�3@	�Ŀ��!?]w����@������ٿ%}�����@�[��P�3@=e񴂐!?
L5���@�^B��ٿh����@�u���3@-�-橐!?ّ}iLO�@�^B��ٿh����@�u���3@-�-橐!?ّ}iLO�@x�/d��ٿ����X�@��+�3@�hN!��!?�Q��@x�/d��ٿ����X�@��+�3@�hN!��!?�Q��@x�/d��ٿ����X�@��+�3@�hN!��!?�Q��@x�/d��ٿ����X�@��+�3@�hN!��!?�Q��@���vٿ�C��@�0����3@�?dM�!??Uy�G�@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@[#c�d�ٿ��M����@�n\R�3@ ���U�!?���@z�)��ٿ��x>��@��{q��3@Ɂl<�!?��yC~B�@z�)��ٿ��x>��@��{q��3@Ɂl<�!?��yC~B�@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�D�i��ٿ�r}��@Un����3@��5� �!?�h�?��@�R����ٿ�ҀghY�@wL�3@կn�^�!?�)�#�@�R����ٿ�ҀghY�@wL�3@կn�^�!?�)�#�@�~W��ٿ�n����@����^�3@b�{p�!?%��O홵@�~W��ٿ�n����@����^�3@b�{p�!?%��O홵@�~W��ٿ�n����@����^�3@b�{p�!?%��O홵@�A,E��ٿ��})))�@�^����3@p'Ѐ��!?�m���W�@ ��㯚ٿ3�_�O��@S�'���3@"jw��!?k�Ys��@���˯�ٿj�Aڡ�@�)��Y�3@������!?1�SS%4�@���˯�ٿj�Aڡ�@�)��Y�3@������!?1�SS%4�@���˯�ٿj�Aڡ�@�)��Y�3@������!?1�SS%4�@���˯�ٿj�Aڡ�@�)��Y�3@������!?1�SS%4�@���˯�ٿj�Aڡ�@�)��Y�3@������!?1�SS%4�@:tG�M�ٿ�2n��U�@j�֒5�3@w����!?;B:4���@:tG�M�ٿ�2n��U�@j�֒5�3@w����!?;B:4���@:tG�M�ٿ�2n��U�@j�֒5�3@w����!?;B:4���@:tG�M�ٿ�2n��U�@j�֒5�3@w����!?;B:4���@���K�ٿDl��l�@q[�:�3@���En�!?�Kܴ@���K�ٿDl��l�@q[�:�3@���En�!?�Kܴ@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�#m�ٿLN^�x�@h�@��3@�;pQ�!?�!�����@�~�	'�ٿS�2	,�@�C�3�3@,�O�i�!?ɾT���@���,��ٿ��_GI�@I��2��3@��a]��!?�*~���@���,��ٿ��_GI�@I��2��3@��a]��!?�*~���@���,��ٿ��_GI�@I��2��3@��a]��!?�*~���@'�ٶz�ٿt�!ŉ�@�m���3@tR�{��!?a���=�@�aYwo�ٿ���fv9�@�7-��3@~̭>�!?���UY׳@�%@�$�ٿ��mO��@�~�`��3@�tڅ�!?p(��	�@�%@�$�ٿ��mO��@�~�`��3@�tڅ�!?p(��	�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@��ozp�ٿ��u����@��ˇ4@v���A�!?���[�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@�Λ�֒ٿ�(�Ŋ�@V9pR��3@��;�7�!?I@�svS�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@]{W�u�ٿN(���@�~�o��3@E�b:�!?qG�Lz8�@s�;�g�ٿ�/���@���aB�3@>���!?�\��F��@s�;�g�ٿ�/���@���aB�3@>���!?�\��F��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@����ٿ1��4���@k���g�3@��h�!?�uo�=��@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@
B��ޖٿ��8��_�@q����3@	LY�!?���-o�@A��/�ٿIٳm��@r=q��3@S� ď!?�Q�Y3�@A��/�ٿIٳm��@r=q��3@S� ď!?�Q�Y3�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@x0r=B�ٿ��G�۵�@ୈ�+�3@��!)�!?���Q�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@�P0�]�ٿ����@�k0(R�3@2��f�!?1�PR�)�@��p���ٿcWx���@��q��3@´yF�!?����@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@o",蜗ٿ�#~�@��&��3@�ǒ�!?�9[$k�@���d�ٿ�����@�.�b��3@���o�!?9\R@���d�ٿ�����@�.�b��3@���o�!?9\R@���d�ٿ�����@�.�b��3@���o�!?9\R@���d�ٿ�����@�.�b��3@���o�!?9\R@���d�ٿ�����@�.�b��3@���o�!?9\R@���d�ٿ�����@�.�b��3@���o�!?9\R@M�����ٿ���w߲�@�+3j+�3@���y�!?��� ��@�a<W��ٿ��!�n��@Z��F�3@��ц�!?,���@�a<W��ٿ��!�n��@Z��F�3@��ц�!?,���@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@l����ٿ5K�z�@+���v�3@<M�P��!?O���#�@�9�,J�ٿ�ؗ~j��@a_����3@�6P3q�!?��7!�@�9�,J�ٿ�ؗ~j��@a_����3@�6P3q�!?��7!�@�9�,J�ٿ�ؗ~j��@a_����3@�6P3q�!?��7!�@�9�,J�ٿ�ؗ~j��@a_����3@�6P3q�!?��7!�@䲓���ٿ]���J�@e���3@s�[�!?K��JdE�@䲓���ٿ]���J�@e���3@s�[�!?K��JdE�@�u�ٿDGg�j��@#��8i�3@�٪��!?��Põ@�u�ٿDGg�j��@#��8i�3@�٪��!?��Põ@���n�ٿH�ƙ1�@�C��W�3@^�1b��!?.A��Nݵ@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@�ʭ��ٿY����@X}���3@f���K�!?�;b�@֎�ٿv�&K�@�u�B��3@��L�!?�Ӵ�:�@֎�ٿv�&K�@�u�B��3@��L�!?�Ӵ�:�@@=+ܐٿ*<v��X�@[����3@چ�B�!?A��b��@@=+ܐٿ*<v��X�@[����3@چ�B�!?A��b��@@=+ܐٿ*<v��X�@[����3@چ�B�!?A��b��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�����ٿMLbhxU�@T��vw�3@�M�w��!?.�~3��@�
����ٿY�&�	�@ ����3@�]�`̐!?a���@�
����ٿY�&�	�@ ����3@�]�`̐!?a���@�
����ٿY�&�	�@ ����3@�]�`̐!?a���@�
����ٿY�&�	�@ ����3@�]�`̐!?a���@�Ry'�ٿ�u"ڿ@V�����3@y�!(��!?���`e�@�Ry'�ٿ�u"ڿ@V�����3@y�!(��!?���`e�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@��,м�ٿ�]����@�q,m�3@�=�Gq�!?�߫9Q�@D�>-�ٿ��s�rο@>l~B�3@��)�!?g�h��@D�>-�ٿ��s�rο@>l~B�3@��)�!?g�h��@D�>-�ٿ��s�rο@>l~B�3@��)�!?g�h��@D�>-�ٿ��s�rο@>l~B�3@��)�!?g�h��@|�b��ٿG��M���@e����3@𝿧)�!?8��;\�@>m4�1�ٿ�0���@K_7�B�3@cET�>�!?0#$Um�@>m4�1�ٿ�0���@K_7�B�3@cET�>�!?0#$Um�@>m4�1�ٿ�0���@K_7�B�3@cET�>�!?0#$Um�@>m4�1�ٿ�0���@K_7�B�3@cET�>�!?0#$Um�@6�LL�ٿG��$�@�����3@B��=�!?���an	�@6�LL�ٿG��$�@�����3@B��=�!?���an	�@6�LL�ٿG��$�@�����3@B��=�!?���an	�@�-��q�ٿ� =&I��@���n��3@���1�!?m�Ǽ�@E��3��ٿ��`����@q��ԥ�3@U`Dڏ!?��=J�ʹ@
2�E"�ٿ�)��@{��`�3@�T`�L�!?��K��Z�@
2�E"�ٿ�)��@{��`�3@�T`�L�!?��K��Z�@
2�E"�ٿ�)��@{��`�3@�T`�L�!?��K��Z�@����I�ٿ�f�(���@&�m��4@���!?�J���N�@����I�ٿ�f�(���@&�m��4@���!?�J���N�@����I�ٿ�f�(���@&�m��4@���!?�J���N�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@j�¶=�ٿ��P-��@��<_�3@w����!?M��ج�@��nZ��ٿ1����@/Y�L4@^1념!?��hk��@F�bL�ٿ�^�?�?�@|�4�4@�8-r�!?L���e�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@����A�ٿS`�5���@u�)�
4@�6��i�!?�b+�=v�@�WP]�ٿ�X���@�CD�<�3@-�DU�!?\鑪�m�@�WP]�ٿ�X���@�CD�<�3@-�DU�!?\鑪�m�@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@;�U<5�ٿ'NK��@�W�K�3@B�|�!?Q$���δ@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@	�n,��ٿ�	TV��@���˾�3@�����!?r��-�@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@�/�b×ٿl�)�c��@����� 4@0n>f��!?�Ɵ�wڴ@����]�ٿ���]�@&��3@�V+:�!?�w�ߔ�@����]�ٿ���]�@&��3@�V+:�!?�w�ߔ�@����]�ٿ���]�@&��3@�V+:�!?�w�ߔ�@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@���V3�ٿu�,S�@�pt�'�3@��U�-�!?*U��y��@\�����ٿJ洬`�@Kd�j�3@	9�	E�!?�d(b���@\�����ٿJ洬`�@Kd�j�3@	9�	E�!?�d(b���@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@F'�+I�ٿ�"���@�6��3@7�󐀐!?El ��õ@`�D��ٿ��4����@�+|N��3@u�����!?��f�e�@`�D��ٿ��4����@�+|N��3@u�����!?��f�e�@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@��lX8�ٿ�T�nE�@�z
���3@�@H�!?��')��@M��ٿ6X��9��@��ՖS�3@|ã���!?H����<�@M��ٿ6X��9��@��ՖS�3@|ã���!?H����<�@M��ٿ6X��9��@��ՖS�3@|ã���!?H����<�@M��ٿ6X��9��@��ՖS�3@|ã���!?H����<�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@i{B���ٿe�6�Kl�@�h�JU�3@N��CB�!?BH���W�@���5`�ٿ�"� ��@�K��t�3@x��X�!?�N��ĵ@9b'�a�ٿ/@��U-�@��T e�3@��@;�!?'�y���@9b'�a�ٿ/@��U-�@��T e�3@��@;�!?'�y���@