�NUMPY v {'descr': '<f8', 'fortran_order': False, 'shape': (3, 10000, 5), }                                                   
������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@B�8�|�ٿ�)T4 ��@���S��3@o,��!? �'�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@8[l�s�ٿ\�����@��+� 4@�|�ޠ�!? Qn@�+�@:N��}�ٿ�{Ǳ���@4;F 4@����!?��$K�+�@:N��}�ٿ�{Ǳ���@4;F 4@����!?��$K�+�@:N��}�ٿ�{Ǳ���@4;F 4@����!?��$K�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@{��K��ٿ�������@��� 4@�+w���!?�Q�X�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@�{]Nٿ#�d����@�`C� 4@ή�CĐ!?(��\�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@��"'��ٿ�]:����@�ǃ 4@�%]0��!?�?�Z�+�@+#�f��ٿ<f)����@q32 4@���!?C��j�+�@+#�f��ٿ<f)����@q32 4@���!?C��j�+�@�nnm��ٿm7Q����@^��9 4@S�j>��!?��$j�+�@�nnm��ٿm7Q����@^��9 4@S�j>��!?��$j�+�@�nnm��ٿm7Q����@^��9 4@S�j>��!?��$j�+�@�nnm��ٿm7Q����@^��9 4@S�j>��!?��$j�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@G�����ٿ��-����@
�� 4@eHf�ΐ!?��3n�+�@�%���ٿ�\�����@��z, 4@)8A��!?'i�+�@���ѯ�ٿ�K�����@փ�Z 4@�Q}ꢐ!?���m�+�@�w���ٿ�������@ 
' 4@�X�&{�!?�O�p�+�@�w���ٿ�������@ 
' 4@�X�&{�!?�O�p�+�@�w���ٿ�������@ 
' 4@�X�&{�!?�O�p�+�@ї0a��ٿ��%����@�cl 4@��ݼ�!?vzq�+�@(Z܁��ٿ/�����@�jij 4@#݃��!?��`s�+�@(Z܁��ٿ/�����@�jij 4@#݃��!?��`s�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@o81U��ٿ�x����@5��; 4@�l��!?&�<i�+�@ȧp��ٿ�@�����@��4 4@>��ѐ!?��e�+�@|ģ�ٿ�������@��H 4@�$���!?�U$_�+�@,��৙ٿ�&����@�y� 4@wy��!?��\�+�@,��৙ٿ�&����@�y� 4@wy��!?��\�+�@��w��ٿb�����@K�T 4@l[ɓ}�!?S�oc�+�@�D���ٿ'�����@]~�, 4@�/�&̐!?�9�Z�+�@vYx��ٿb/����@��"� 4@���!?�\n\�+�@vYx��ٿb/����@��"� 4@���!?�\n\�+�@��h]��ٿĔ����@=#-� 4@l>�:��!?��\S�+�@��h]��ٿĔ����@=#-� 4@l>�:��!?��\S�+�@
o����ٿ+�t ��@Y?� 4@��\ϐ!?Iz�R�+�@9c>��ٿ��: ��@k�)�  4@�G%�ݐ!?�3�U�+�@9c>��ٿ��: ��@k�)�  4@�G%�ݐ!?�3�U�+�@0��c��ٿ=y	 ��@#��= 4@!����!?3	�O�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@���g��ٿJS! ��@g ��  4@߄���!?���G�+�@�Ҥ�ٿ�3" ��@�.8�  4@�r�~l�!?Zs�>�+�@�J�ՠ�ٿv� ��@HC��  4@6��x�!?��;�+�@�lb��ٿ��Z ��@��8�  4@s�B��!?�T�=�+�@�lb��ٿ��Z ��@��8�  4@s�B��!?�T�=�+�@r�*��ٿD ��@�5tk  4@��[��!?���?�+�@���מ�ٿA�9����@�.O  4@Ve���!?�&K�+�@���מ�ٿA�9����@�.O  4@Ve���!?�&K�+�@]*6��ٿ�96  ��@���=  4@�A�$��!? ��G�+�@?�$���ٿ�	*����@a?�~  4@	�1��!?� �C�+�@?�$���ٿ�	*����@a?�~  4@	�1��!?� �C�+�@?�$���ٿ�	*����@a?�~  4@	�1��!?� �C�+�@-~�W��ٿSb����@��a�  4@����{�!?:mF�+�@�;ޟ�ٿ}1Q����@#}��  4@v�`ΐ!?�@
G�+�@�;ޟ�ٿ}1Q����@#}��  4@v�`ΐ!?�@
G�+�@��z���ٿܢ3����@])�^  4@����!?ü�J�+�@��z���ٿܢ3����@])�^  4@����!?ü�J�+�@��z���ٿܢ3����@])�^  4@����!?ü�J�+�@�ͭn��ٿ������@�w�x  4@ъ$2�!?�<M�+�@0�rj��ٿ�1����@��R�  4@я��(�!?:ɏQ�+�@�	��ٿr7�����@:�h	 4@��~��!?qYQ�+�@j{���ٿ>4����@�'= 4@#�c.?�!?@��N�+�@�n���ٿ�˗����@O$Y 4@:�z���!?p��S�+�@�K���ٿ������@zA�o 4@S?&��!?1t�R�+�@�K���ٿ������@zA�o 4@S?&��!?1t�R�+�@������ٿɓ�����@ΑBW 4@}�A��!?d�V�+�@�����ٿ؈X����@��H� 4@ �5g�!?��9T�+�@�����ٿ؈X����@��H� 4@ �5g�!?��9T�+�@�ҠR��ٿ�f3����@���* 4@oZ���!?�S�I�+�@�&�ߡ�ٿ�/s ��@��Q�  4@��>�&�!?(1F�+�@�IpH��ٿBY� ��@ڟ�A 4@���~Ր!?�F�+�@����ٿ��  ��@�\�  4@m�����!?�s�?�+�@$%�ݛ�ٿ�u�	 ��@�+u!  4@c|��q�!?�HQ=�+�@$%�ݛ�ٿ�u�	 ��@�+u!  4@c|��q�!?�HQ=�+�@$%�ݛ�ٿ�u�	 ��@�+u!  4@c|��q�!?�HQ=�+�@^ᤜ�ٿQv�	 ��@T��g  4@eUGc��!?VVmA�+�@��u���ٿ_�� ��@6E�k  4@Nk��!?N�7<�+�@��u���ٿ_�� ��@6E�k  4@Nk��!?N�7<�+�@�[����ٿ��� ��@]��h  4@�Gg��!?DA�+�@:�럙ٿ/� ��@�rv�  4@�]ŝ��!?N{B�+�@:�럙ٿ/� ��@�rv�  4@�]ŝ��!?N{B�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@�.�Ӡ�ٿ��� ��@�q��  4@���i�!?��>�+�@}�K���ٿ�@�	 ��@#�ݶ  4@b4��|�!? e�>�+�@��?,��ٿC�� ��@�'fm  4@��N���!?��<�+�@b/���ٿ�"� ��@!�  4@��uᐐ!?���>�+�@b/���ٿ�"� ��@!�  4@��uᐐ!?���>�+�@��[���ٿ��� ��@~��  4@ƽ͹�!?��B�+�@�T[X��ٿ	�A ��@Z�B�  4@���VÐ!?	�jB�+�@�PG1��ٿB~F ��@^��  4@
u:g�!?�X�<�+�@&��Ǟ�ٿ�~d ��@���  4@�M�b�!?�V�7�+�@&��Ǟ�ٿ�~d ��@���  4@�M�b�!?�V�7�+�@&��Ǟ�ٿ�~d ��@���  4@�M�b�!?�V�7�+�@l�(��ٿ�C4 ��@�,�  4@��q�u�!?�+H:�+�@+�<䝙ٿ	�� ��@f�  4@Գd���!?"F�=�+�@��Bќ�ٿ��� ��@p��r  4@�~�Ǻ�!?ކ�B�+�@�>ޞ�ٿZ� ��@�d�  4@ڶ�ԝ�!?h��@�+�@9�#e��ٿ�µ ��@\�w�  4@=�ĝ�!?�3�>�+�@9�׍��ٿm�I  ��@����  4@��h���!?�~>�+�@*>XH��ٿ������@)[ 9 4@��뎿�!?���@�+�@�O�`��ٿ,{P����@ݼ
V 4@����!?-�@�+�@�O�`��ٿ,{P����@ݼ
V 4@����!?-�@�+�@�����ٿη�����@)�% 4@�j��O�!?�̛>�+�@�����ٿη�����@)�% 4@�j��O�!?�̛>�+�@M���ٿ������@��$ 4@E_W�/�!?��=�+�@�	��ٿ8�� ��@����  4@$�3�!?x#�:�+�@�	��ٿ8�� ��@����  4@$�3�!?x#�:�+�@�	��ٿ8�� ��@����  4@$�3�!?x#�:�+�@����ٿ��� ��@����  4@d�=�G�!?I�2�+�@p����ٿ�J� ��@�CZ�  4@Q��M�!?681�+�@��l��ٿ�� ��@����  4@���\�!?��R4�+�@��l��ٿ�� ��@����  4@���\�!?��R4�+�@��l��ٿ�� ��@����  4@���\�!?��R4�+�@�C���ٿ\4� ��@ཌ�  4@*�=��!?�1�2�+�@�h�à�ٿ�u� ��@�C��  4@%�!? 3�4�+�@fH,���ٿb� ��@��Ĳ  4@�����!?hC:�+�@ �H���ٿ�r ��@��  4@�d7sƐ!?��4?�+�@�`lӠ�ٿ5Zr  ��@^rx�  4@:��H��!?�>�+�@QB���ٿ8�T ��@���  4@��~�Ɛ!?Vsy?�+�@Nbۤ��ٿ�_�����@`�t�  4@O����!?�߳F�+�@�S����ٿ442����@}k  4@j�ƍ��!?��rF�+�@'+����ٿZYp����@�! 4@R+�ѐ!?�?E�+�@͡IV��ٿ@d�����@��8�  4@��P��!?W>XH�+�@͡IV��ٿ@d�����@��8�  4@��P��!?W>XH�+�@P�����ٿ�������@���  4@D��E��!?��I�+�@�]>��ٿ�� ��@n�<�  4@�ϟ��!?�A/I�+�@m�o���ٿ��"����@I%:
 4@[.���!?1K�+�@m�o���ٿ��"����@I%:
 4@[.���!?1K�+�@��j���ٿx� ��@�jW 4@��7&��!?)]>E�+�@��j���ٿx� ��@�jW 4@��7&��!?)]>E�+�@��j���ٿx� ��@�jW 4@��7&��!?)]>E�+�@���휙ٿV�o ��@����  4@�eo��!?���?�+�@��>ܛ�ٿف�  ��@9�� 4@k��9��!?g�I�+�@=4�x��ٿ�$o  ��@"� 4@�~���!?2uF�+�@�����ٿͩ�����@�7z�  4@�5��!?���E�+�@��֠�ٿy.�����@�?A�  4@�S�U��!?��H�+�@���q��ٿ�u�����@&�4�  4@�Ӹ��!?�4SO�+�@Vƙ��ٿ�W�����@zRN�  4@�\��!?�}LR�+�@������ٿ�,�����@2���  4@�1����!?b�RV�+�@;.����ٿ������@����  4@���!?�i^Y�+�@�)fՙ�ٿ�3�����@�e�  4@�r���!?4އ[�+�@�H��ٿ������@is`�  4@��Vwm�!?�RbY�+�@�H��ٿ������@is`�  4@��Vwm�!?�RbY�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@5뽛��ٿ^B����@q��  4@8{ch�!?���P�+�@\�7�ٿS��  ��@���  4@�w�<T�!?hP�+�@ 
��ٿ��� ��@pS��  4@&$��r�!?6>:H�+�@�x���ٿ�"7 ��@�:k�  4@I����!?=�zH�+�@e2���ٿɇ� ��@xt8�  4@��8��!?���H�+�@9��ٿ�Qe ��@��u�  4@]���!?G��I�+�@9����ٿ+�� ��@��  4@��Z���!?��yU�+�@�Ʈ���ٿ�a� ��@�vi�  4@1㶐!?��=W�+�@:%�8��ٿ���  ��@O�T
 4@8����!?5M�Z�+�@��rc��ٿ� ����@� 4@�R��!?*�X�+�@<�9ԟ�ٿm�4 ��@�*��  4@1��ސ!?7^�Q�+�@�f�⠙ٿX� ��@jR<�  4@Ȍ���!?��WJ�+�@E�c���ٿ!� ��@�a�  4@|��P+�!?c�WL�+�@E�c���ٿ!� ��@�a�  4@|��P+�!?c�WL�+�@����ٿ��H ��@��s�  4@�iD��!?��J�+�@��?��ٿ�� ��@��R  4@!��gB�!?�VF�+�@����ٿu�� ��@l�W 4@pqd&O�!?�9@�+�@����ٿu�� ��@l�W 4@pqd&O�!?�9@�+�@��Ȯ��ٿ�C` ��@VX 4@,W5�Q�!?�R[A�+�@��Ȯ��ٿ�C` ��@VX 4@,W5�Q�!?�R[A�+�@��Y'��ٿ��O ��@��a# 4@��l�k�!?�C�+�@��Y'��ٿ��O ��@��a# 4@��l�k�!?�C�+�@��Y'��ٿ��O ��@��a# 4@��l�k�!?�C�+�@��Mr��ٿ�P� ��@�y�/ 4@:�vK�!?�{J�+�@gbt��ٿ06  ��@s�2 4@A,�/J�!?���I�+�@gbt��ٿ06  ��@s�2 4@A,�/J�!?���I�+�@gbt��ٿ06  ��@s�2 4@A,�/J�!?���I�+�@p-�ܟ�ٿ�[ ��@bZ��  4@��+'�!?o!B�+�@p-�ܟ�ٿ�[ ��@bZ��  4@��+'�!?o!B�+�@��͠�ٿ���
 ��@���  4@*{�r�!?]5;�+�@�cp��ٿ"t ��@<��  4@Қ���!?ppKC�+�@�cp��ٿ"t ��@<��  4@Қ���!?ppKC�+�@�%���ٿ}N�
 ��@{<�  4@�7C�!?�޼A�+�@��=E��ٿ�� ��@E	}�  4@�.)��!??̓A�+�@��1��ٿ#T�	 ��@+��  4@�% �!?��C�+�@� j��ٿr�� ��@�w�  4@$����!?��:�+�@_j�ã�ٿ��\ ��@	H  4@�l��ܐ!?r/�=�+�@��IΣ�ٿ�. ��@�W�  4@;b�֐!?os�:�+�@��IΣ�ٿ�. ��@�W�  4@;b�֐!?os�:�+�@��IΣ�ٿ�. ��@�W�  4@;b�֐!?os�:�+�@��5���ٿgf9 ��@������3@���k��!?�f6�+�@opٿp� ��@!}����3@NlU��!?��0�+�@�8Ue��ٿoi� ��@v�9���3@V��ې!?��V5�+�@?����ٿ�2 ��@��֫��3@����!?0��=�+�@:��̩�ٿnb� ��@ġ���3@���n%�!?Qo�9�+�@:��̩�ٿnb� ��@ġ���3@���n%�!?Qo�9�+�@f�87��ٿU�� ��@�����3@�0�1��!?��+9�+�@f�87��ٿU�� ��@�����3@�0�1��!?��+9�+�@f�87��ٿU�� ��@�����3@�0�1��!?��+9�+�@_����ٿ
�! ��@yn���3@���!?�)�2�+�@���ͯ�ٿ���$ ��@��JW��3@��4��!?Y�-�+�@���ͯ�ٿ���$ ��@��JW��3@��4��!?Y�-�+�@���ͯ�ٿ���$ ��@��JW��3@��4��!?Y�-�+�@���ͯ�ٿ���$ ��@��JW��3@��4��!?Y�-�+�@���ͯ�ٿ���$ ��@��JW��3@��4��!?Y�-�+�@�(�׭�ٿ��~ ��@������3@�}���!?��&�+�@<yO��ٿ�l�% ��@Tz����3@�#O��!?�� �+�@<yO��ٿ�l�% ��@Tz����3@�#O��!?�� �+�@<yO��ٿ�l�% ��@Tz����3@�#O��!?�� �+�@<yO��ٿ�l�% ��@Tz����3@�#O��!?�� �+�@a?���ٿb�( ��@G�JM��3@��V��!?��/!�+�@�����ٿ� �  ��@Z���3@R��7��!?���-�+�@�����ٿ�5 ��@1�3k��3@ڵh0Ð!?;��-�+�@T�x���ٿ���  ��@ɘԹ��3@��Տ`�!?�͚4�+�@T�x���ٿ���  ��@ɘԹ��3@��Տ`�!?�͚4�+�@�/3j��ٿ��� ��@'�����3@}��[�!?�k.@�+�@t�H��ٿZ�  ��@�o4���3@�� ��!?�_w<�+�@t�H��ٿZ�  ��@�o4���3@�� ��!?�_w<�+�@t�H��ٿZ�  ��@�o4���3@�� ��!?�_w<�+�@t�H��ٿZ�  ��@�o4���3@�� ��!?�_w<�+�@��7u��ٿ���) ��@͒�,��3@Z[�D��!?�Y�'�+�@�����ٿ�</ ��@�#���3@'\Ǖn�!?��(�+�@�����ٿ�</ ��@�#���3@'\Ǖn�!?��(�+�@���|��ٿ��� ��@Ǻ���3@���(��!?t�I7�+�@�wQP��ٿ���' ��@_v���3@��`�!?v�
&�+�@ ���ٿ��K ��@�9���3@/6`���!?��/3�+�@r|bǥ�ٿ⬧ ��@���_  4@�֑�>�!?�dI�+�@���ٿ�c ��@|����3@A�AF8�!?��?�+�@<h�]��ٿ��� ��@� �X  4@ZeA�9�!?�8�F�+�@<h�]��ٿ��� ��@� �X  4@ZeA�9�!?�8�F�+�@��1��ٿ�)� ��@�RԾ��3@{Tøǐ!?/22�+�@��1��ٿ�)� ��@�RԾ��3@{Tøǐ!?/22�+�@�F����ٿ���	 ��@'H��  4@+2�Ɛ!?9
IB�+�@�F����ٿ���	 ��@'H��  4@+2�Ɛ!?9
IB�+�@&sE���ٿ{�+ ��@~��J  4@!oO��!?�v@�+�@�ۥ�ٿҁ� ��@&o(���3@t����!?Ru�7�+�@nĘ���ٿ8/� ��@��IT  4@��C�Ӑ!?|�@�+�@���*��ٿ?q� ��@F�=p��3@�IƮ�!?{��.�+�@��B��ٿ�E ��@_F6  4@�H�6��!?���H�+�@��B��ٿ�E ��@_F6  4@�H�6��!?���H�+�@�
����ٿ������@�>�- 4@ v�# �!?��b�+�@�
����ٿ������@�>�- 4@ v�# �!?��b�+�@�
����ٿ������@�>�- 4@ v�# �!?��b�+�@�
����ٿ������@�>�- 4@ v�# �!?��b�+�@����ٿ�Ӄ ��@9�$  4@�_�oƐ!?�a�+�@��L��ٿMz}	 ��@V����3@'�傐!?>I�^�+�@�M���ٿ�Y� ��@���a  4@��!?���S�+�@���:��ٿ�t% ��@�H�E  4@�y�#Ő!?��@�+�@��#��ٿ�{ ��@`�(&  4@�Ajǐ!?��OG�+�@D��ϛ�ٿ�"�  ��@\D�d 4@ǎ]3��!?l^0J�+�@��a֓�ٿ�9;����@Е�L 4@��.��!?�cWP�+�@��a֓�ٿ�9;����@Е�L 4@��.��!?�cWP�+�@Û.���ٿ�n$����@��p 4@nN��!?�{�W�+�@�q��ٿ[�c����@��R� 4@�,*ʐ!?s�I�+�@��a��ٿK�-����@O�� 4@a�D���!?�6F�+�@5�"~�ٿ�9p����@�� 4@]c����!?8��U�+�@5�"~�ٿ�9p����@�� 4@]c����!?8��U�+�@�a�ޓ�ٿ� �����@x�0 4@�@��А!?�^H�+�@�a�ޓ�ٿ� �����@x�0 4@�@��А!?�^H�+�@^�N$��ٿ�%8����@Wx� 4@��>q��!?j�Y�+�@^�N$��ٿ�%8����@Wx� 4@��>q��!?j�Y�+�@�~�s��ٿY�����@{�� 4@z�dɐ!?��eK�+�@.�x��ٿd�` ��@ǋl0��3@��UGʐ!?37�+�@.�x��ٿd�` ��@ǋl0��3@��UGʐ!?37�+�@.�x��ٿd�` ��@ǋl0��3@��UGʐ!?37�+�@�^����ٿ%3�	 ��@��ۜ��3@F1ԧ��!?Q{'<�+�@�^����ٿ%3�	 ��@��ۜ��3@F1ԧ��!?Q{'<�+�@Z�ڊ��ٿ��U����@؝	[ 4@X`?i��!?�\�:�+�@Z�ڊ��ٿ��U����@؝	[ 4@X`?i��!?�\�:�+�@����ٿ�������@���	 4@7�w�!?�u84�+�@����ٿ�������@���	 4@7�w�!?�u84�+�@���˃�ٿ�������@�	�N 4@Q��!?�A�-�+�@����ٿ.������@�d�s 4@(�����!?���'�+�@�_�ٿ6T ��@����3@ˆ���!?���+�@�_�ٿ6T ��@����3@ˆ���!?���+�@f��ٿBfP ��@���]��3@������!?BЄ�+�@N����ٿ&�� ��@ғ  4@�#�y��!?�w��+�@P4�ٿ"Ҳ����@���v 4@r�'�!?�5���+�@��ӎ��ٿ߂+����@M��P 4@�s��!?q���+�@��ӎ��ٿ߂+����@M��P 4@�s��!?q���+�@� t�ٿ#�+����@�L� 4@+bF ��!?�	��+�@�x�ٿ�������@�t� 4@�B���!?�J �+�@�m7r�ٿ��|����@�P 4@��r�!?�Q�+�@�!=��ٿ�WJ����@�^.@ 4@��u(��!?�6cT�+�@�S���ٿF������@&�l 4@�o^ǋ�!?D��c�+�@)�v�ٿ�����@�� 4@l'S��!?!�b�+�@)�v�ٿ�����@�� 4@l'S��!?!�b�+�@�|����ٿy�����@�8�� 4@����!?�4��+�@��4�p�ٿɒƶ���@�ܟ� 4@�侷��!?0���+�@����k�ٿ�ʭ���@P>�	 4@��<���!?�W�t�+�@����k�ٿ�ʭ���@P>�	 4@��<���!?�W�t�+�@��5z�ٿ43����@�f]� 4@�e���!?C����+�@��X��ٿ�I����@ػL 4@Z���Ր!?�����+�@��X��ٿ�I����@ػL 4@Z���Ր!?�����+�@��jfr�ٿ�3/����@/�� 4@C�E��!?�nρ�+�@�5]\�ٿp�����@="-U 4@��u��!?����+�@�5]\�ٿp�����@="-U 4@��u��!?����+�@�5]\�ٿp�����@="-U 4@��u��!?����+�@m�r�ٿ������@%wɩ 4@o1���!?����+�@m�r�ٿ������@%wɩ 4@o1���!?����+�@m�r�ٿ������@%wɩ 4@o1���!?����+�@�j8y�ٿ]�����@�G�@ 4@�y��ː!?��Oo�+�@��CT��ٿ�������@��U� 4@�/���!?���+�@�GIٿ��Q����@0g�� 4@�7֓�!?9	-��+�@4X#{��ٿ�����@�CE 4@X�z-�!?�"L�+�@7�bh��ٿ�E����@M��� 4@�Ƴ�!?��D�+�@7�bh��ٿ�E����@M��� 4@�Ƴ�!?��D�+�@7�bh��ٿ�E����@M��� 4@�Ƴ�!?��D�+�@S�O_��ٿP������@�R 4@�����!?���+�@S�O_��ٿP������@�R 4@�����!?���+�@S�O_��ٿP������@�R 4@�����!?���+�@���X��ٿ�Ѷ ��@�B�  4@-!qސ!?��Pu�+�@R��A��ٿM) ��@) cH��3@F� +�!?��=�+�@R��A��ٿM) ��@) cH��3@F� +�!?��=�+�@�g�=��ٿ�����@ن�r 4@S��r��!?J�=�+�@�C���ٿG*b ��@����  4@ƪ�3�!?EF��+�@ǃ��ٿŗ�  ��@@d�� 4@�7�o�!?�6��+�@f:��z�ٿ.;|����@��2> 4@Dk���!?g�Z.�+�@aUS���ٿQ�����@�C< 4@�.N�֐!?���+�@��)悙ٿ
�����@��E 4@�]��ϐ!?dC� �+�@��)悙ٿ
�����@��E 4@�]��ϐ!?dC� �+�@��Y���ٿ�P����@�F� 4@�����!?��0X�+�@��Y���ٿ�P����@�F� 4@�����!?��0X�+�@��Y���ٿ�P����@�F� 4@�����!?��0X�+�@��ֈ~�ٿw�v����@��M0 4@�)Kː!?5q��+�@�����ٿI]#����@�@x� 4@̵Pڐ!?����+�@�*c�ٿ������@�m�
 4@Pv�~�!?.�"�+�@����k�ٿ̤����@[1� 4@��Տ��!?�x���+�@Û7�]�ٿ�E�����@6�!E	 4@�Qz�Ȑ!?V�3��+�@tYT�M�ٿ���]���@�r=L 4@�j��!?6� ��+�@�FYE�ٿ|�e���@0W� 4@!"��!?��F��+�@�FYE�ٿ|�e���@0W� 4@!"��!?��F��+�@SX�ٿ�m�����@�G�� 4@��BrJ�!?���+�@�vmd#�ٿ��H*���@lM̢ 4@��:-�!?�Q��+�@>r+G�ٿ޿.P���@�BV� 4@��c��!??����+�@_so瑙ٿ�o� ��@��G� 4@��W���!?�/���+�@_so瑙ٿ�o� ��@��G� 4@��W���!?�/���+�@��z3~�ٿUs ��@ȍ� 4@1�}�D�!?�W�+�@��z3~�ٿUs ��@ȍ� 4@1�}�D�!?�W�+�@��z3~�ٿUs ��@ȍ� 4@1�}�D�!?�W�+�@I:&P�ٿzӉ����@�b{ 4@m?v�!?��tj�+�@.�G莙ٿ�`�����@<%v� 4@f����!? gIC�+�@�F��ٿ�ܖ���@?� 4@����!?��Mx�+�@�F��ٿ�ܖ���@?� 4@����!?��Mx�+�@�F��ٿ�ܖ���@?� 4@����!?��Mx�+�@�b	ϙٿ�u�����@��]R��3@���t�!?F�|��+�@���\��ٿY�W5���@��z 4@�5XHݐ!?:Z��+�@��)-��ٿjR�����@���'  4@g8�a�!?��
�+�@��)-��ٿjR�����@���'  4@g8�a�!?��
�+�@��)-��ٿjR�����@���'  4@g8�a�!?��
�+�@�m�ܙٿre�����@ d}��3@�De�Ӑ!?�v�d�+�@�m�ܙٿre�����@ d}��3@�De�Ӑ!?�v�d�+�@���8ݙٿ\EQ ��@fR��3@���ѐ!?/���+�@�`����ٿ���" ��@�q�u��3@O섓�!?b/�Z�+�@Fc:��ٿ�������@<�����3@/�b�!?M�w��+�@?�gpq�ٿ\Pj���@��	 4@W��4�!?�h5��+�@?�gpq�ٿ\Pj���@��	 4@W��4�!?�h5��+�@?�gpq�ٿ\Pj���@��	 4@W��4�!?�h5��+�@?�gpq�ٿ\Pj���@��	 4@W��4�!?�h5��+�@��!F��ٿ�i�E���@���% 4@�}^�!?F�)��+�@	�A��ٿ�(<���@����	 4@�,�߈�!?ȨF��+�@	�A��ٿ�(<���@����	 4@�,�߈�!?ȨF��+�@|�\�F�ٿ�������@�� 4@ �(u�!?ޤ��+�@?"b�a�ٿj|�����@�ò 4@t�����!?]����+�@?"b�a�ٿj|�����@�ò 4@t�����!?]����+�@v ���ٿ؟|����@yS�� 4@幌�!?6Xk��+�@v ���ٿ؟|����@yS�� 4@幌�!?6Xk��+�@v ���ٿ؟|����@yS�� 4@幌�!?6Xk��+�@�v�<ęٿ)��T���@\ʦ� 4@�y��!?<f|y�+�@K��ϙٿA��F���@Q�	 4@�"�ԯ�!?!m���+�@K��ϙٿA��F���@Q�	 4@�"�ԯ�!?!m���+�@a$�/ۙٿ$gY����@�� 4@D�VĐ!?y��\�+�@a$�/ۙٿ$gY����@�� 4@D�VĐ!?y��\�+�@a$�/ۙٿ$gY����@�� 4@D�VĐ!?y��\�+�@=/�Aۙٿ���y���@��� 4@ F��Ӑ!?���+�@=/�Aۙٿ���y���@��� 4@ F��Ӑ!?���+�@���ٿ�����@\�� 4@�"���!?��ad�+�@���ٿ�����@\�� 4@�"���!?��ad�+�@���ٿ�����@\�� 4@�"���!?��ad�+�@���ٿ�����@\�� 4@�"���!?��ad�+�@���ٿ�����@\�� 4@�"���!?��ad�+�@��řٿ�eD���@�]��3@p�ː!?��H	�+�@��řٿ�eD���@�]��3@p�ː!?��H	�+�@��řٿ�eD���@�]��3@p�ː!?��H	�+�@`���p�ٿH����@��F��3@����!?1l�_�+�@I��׆�ٿǟ� ��@7���3@Jҥ�g�!?��`5�+�@Q�$~�ٿ8k����@���U��3@��y�u�!?杞�+�@Q�$~�ٿ8k����@���U��3@��y�u�!?杞�+�@���ٿ<Z�k ��@*���3@�8Cٽ�!?qw�+�@� �S��ٿo�P���@Z�	��3@���i��!?Q*{��+�@� �S��ٿo�P���@Z�	��3@���i��!?Q*{��+�@T�n?�ٿ��7� ��@�����3@B��H�!?n�o��+�@��
���ٿ��O/��@gkx͎�3@S�l�x�!?�)���+�@��
���ٿ��O/��@gkx͎�3@S�l�x�!?�)���+�@��
���ٿ��O/��@gkx͎�3@S�l�x�!?�)���+�@��
���ٿ��O/��@gkx͎�3@S�l�x�!?�)���+�@o�V��ٿ�����@ͽ�9��3@��|zu�!?Jk:��+�@P���P�ٿ~~���@��CX�3@��N4K�!?y:���+�@P���P�ٿ~~���@��CX�3@��N4K�!?y:���+�@P���P�ٿ~~���@��CX�3@��N4K�!?y:���+�@��u>B�ٿ
j�����@�O� 4@�3:ΐ!?���M�+�@��ٿ߿n��@G%�4��3@�2-j!?p���+�@��ٿ߿n��@G%�4��3@�2-j!?p���+�@��ٿ߿n��@G%�4��3@�2-j!?p���+�@���̾�ٿ$\�����@rB��P 4@��%!��!?�����+�@���̾�ٿ$\�����@rB��P 4@��%!��!?�����+�@���̾�ٿ$\�����@rB��P 4@��%!��!?�����+�@�}��!�ٿ��;���@~�_�� 4@�Qq�!?����+�@�}��!�ٿ��;���@~�_�� 4@�Qq�!?����+�@�}��!�ٿ��;���@~�_�� 4@�Qq�!?����+�@�}��!�ٿ��;���@~�_�� 4@�Qq�!?����+�@�}��!�ٿ��;���@~�_�� 4@�Qq�!?����+�@��ژٿ.]����@����g 4@P�&:��!?��^��+�@Mg�B�ٿA��� ��@^<+��3@������!?˹X��+�@Mg�B�ٿA��� ��@^<+��3@������!?˹X��+�@Mg�B�ٿA��� ��@^<+��3@������!?˹X��+�@���?ܙٿ4�����@x�m���3@��Rڏ�!?�C���+�@���?ܙٿ4�����@x�m���3@��Rڏ�!?�C���+�@���?ܙٿ4�����@x�m���3@��Rڏ�!?�C���+�@�k��ٿ��9���@I��w� 4@!���!?��5�+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@G�<��ٿ��K����@{&�ʮ 4@:3X��!? {9��+�@@�ܫ��ٿ�0���@<�FjN4@hi��!?'����+�@���1��ٿsc(��@f j��4@�ﯭ�!?#_^�+�@���1��ٿsc(��@f j��4@�ﯭ�!?#_^�+�@���1��ٿsc(��@f j��4@�ﯭ�!?#_^�+�@ì>Ƶ�ٿ���B���@Y�x4@�p��.�!?'��+�@ì>Ƶ�ٿ���B���@Y�x4@�p��.�!?'��+�@��S��ٿ:sc��@��8��4@�DZ�K�!?4�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��%w�ٿۢ����@�:\��4@3yV&K�!?��9�+�@��!v��ٿq8i���@TG@54@�Fbzѐ!?�����+�@��!v��ٿq8i���@TG@54@�Fbzѐ!?�����+�@��!v��ٿq8i���@TG@54@�Fbzѐ!?�����+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@=Y�ȥ�ٿU\IZ͇�@
"dع4@��r�!?�V��+�@�u�S+�ٿ^�}���@��3=�4@,�߳!?M�L�+�@�u�S+�ٿ^�}���@��3=�4@,�߳!?M�L�+�@;TQ�ȇٿ��Ǚɇ�@! �4@�����!?�P�,�@;TQ�ȇٿ��Ǚɇ�@! �4@�����!?�P�,�@;TQ�ȇٿ��Ǚɇ�@! �4@�����!?�P�,�@;TQ�ȇٿ��Ǚɇ�@! �4@�����!?�P�,�@;TQ�ȇٿ��Ǚɇ�@! �4@�����!?�P�,�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@L�Oi��ٿ��͇�@/��?4@�)?ؐ!?�����+�@m:\��ٿt��Q͇�@�
���4@��.��!?���+�@�:?�݈ٿ;`��·�@��!w4@���Ȑ!?6�Y��+�@�:?�݈ٿ;`��·�@��!w4@���Ȑ!?6�Y��+�@�:?�݈ٿ;`��·�@��!w4@���Ȑ!?6�Y��+�@�:?�݈ٿ;`��·�@��!w4@���Ȑ!?6�Y��+�@;�鹅ٿ�Y*NÇ�@q��	4@�A��!?:�6�,�@;�鹅ٿ�Y*NÇ�@q��	4@�A��!?:�6�,�@?K����ٿ��0�Ç�@��]�=	4@7֎���!?k�q�,�@?K����ٿ��0�Ç�@��]�=	4@7֎���!?k�q�,�@?K����ٿ��0�Ç�@��]�=	4@7֎���!?k�q�,�@?K����ٿ��0�Ç�@��]�=	4@7֎���!?k�q�,�@?K����ٿ��0�Ç�@��]�=	4@7֎���!?k�q�,�@P���Q�ٿ�0����@���s4@�� ��!?�x�+�@P���Q�ٿ�0����@���s4@�� ��!?�x�+�@P���Q�ٿ�0����@���s4@�� ��!?�x�+�@P���Q�ٿ�0����@���s4@�� ��!?�x�+�@P���Q�ٿ�0����@���s4@�� ��!?�x�+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@�T�3�ٿ�C����@�
y�D4@s���!?�����+�@��tu�ٿ�����@S���4@jeu3��!?��%*�+�@{}|�o�ٿ�K�W߇�@F*ǪP4@.�!��!?)���+�@{}|�o�ٿ�K�W߇�@F*ǪP4@.�!��!?)���+�@}o(ڌٿ����ه�@�P��4@�/^%ؐ!?��eI�+�@}o(ڌٿ����ه�@�P��4@�/^%ؐ!?��eI�+�@}o(ڌٿ����ه�@�P��4@�/^%ؐ!?��eI�+�@�إ���ٿ�B�ȇ�@5&�N4@�f᧐!?�>\�,�@�إ���ٿ�B�ȇ�@5&�N4@�f᧐!?�>\�,�@�إ���ٿ�B�ȇ�@5&�N4@�f᧐!?�>\�,�@�إ���ٿ�B�ȇ�@5&�N4@�f᧐!?�>\�,�@�@�Y�ٿ;�����@�L{��	4@tn���!?�JJ!,�@�@�Y�ٿ;�����@�L{��	4@tn���!?�JJ!,�@�@�Y�ٿ;�����@�L{��	4@tn���!?�JJ!,�@�@�Y�ٿ;�����@�L{��	4@tn���!?�JJ!,�@�@�Y�ٿ;�����@�L{��	4@tn���!?�JJ!,�@�Q,1�{ٿH���@��Q\4@�|�!?Q�&�,�@�Q,1�{ٿH���@��Q\4@�|�!?Q�&�,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@m3���ٿ+z�hƇ�@ٿ��4@[�&��!?��$,�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@0q��L�ٿ�|��ׇ�@����4@�9ؿ�!?x��F�+�@
ǧ�-�ٿ�J���@iA~94@f�%�!?�s���+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@&<s�b�ٿ&��U��@��r�c4@�0�ʐ!?���_�+�@�=�{��ٿ��K���@��μ	4@&S&}!?�T#,�@�=�{��ٿ��K���@��μ	4@&S&}!?�T#,�@�=�{��ٿ��K���@��μ	4@&S&}!?�T#,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@����ٿs��ʇ�@�`Xf�4@z��{o�!?>�,,�@M)ȯ�ٿ�Rn~���@�N���	4@����!?�.�2!,�@M)ȯ�ٿ�Rn~���@�N���	4@����!?�.�2!,�@l��ٿA ��ˇ�@6,�J4@9�/�\�!?�ϔI,�@꼟��ٿO�{�Ƈ�@>�?�4@L�5q�!?�2X�%,�@꼟��ٿO�{�Ƈ�@>�?�4@L�5q�!?�2X�%,�@��L�ٿ�{�鱇�@pg#�>
4@3�)ɰ�!?f�0�/,�@��L�ٿ�{�鱇�@pg#�>
4@3�)ɰ�!?f�0�/,�@�S�f��ٿ8߬�ɇ�@�/�:4@]��g��!?m��S",�@�S�f��ٿ8߬�ɇ�@�/�:4@]��g��!?m��S",�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@͵��ٿ6-Ok��@�.4@�ۿDѐ!?Fpl}�+�@:�OT"�ٿ��$��@x䣱�4@�4�վ�!?;���+�@:�OT"�ٿ��$��@x䣱�4@�4�վ�!?;���+�@:�OT"�ٿ��$��@x䣱�4@�4�վ�!?;���+�@:�OT"�ٿ��$��@x䣱�4@�4�վ�!?;���+�@:�OT"�ٿ��$��@x䣱�4@�4�վ�!?;���+�@U\犅ٿ`m����@���C4@Y�����!?�l��+�@U\犅ٿ`m����@���C4@Y�����!?�l��+�@U\犅ٿ`m����@���C4@Y�����!?�l��+�@U\犅ٿ`m����@���C4@Y�����!?�l��+�@U\犅ٿ`m����@���C4@Y�����!?�l��+�@�`�0�ٿ�y��ۇ�@���)F4@*�Jǐ!?=��+�@�`�0�ٿ�y��ۇ�@���)F4@*�Jǐ!?=��+�@�`�0�ٿ�y��ۇ�@���)F4@*�Jǐ!?=��+�@��:?��ٿ>���@-�Q��4@yN��!?ù#��+�@��u�ٿG`,ه�@IT�9�4@2j�M��!? ���+�@��u�ٿG`,ه�@IT�9�4@2j�M��!? ���+�@��u�ٿG`,ه�@IT�9�4@2j�M��!? ���+�@:����ٿ�{bއ�@~bv/�4@E�W���!?i��+�@8!�Ɲ�ٿ�rW��@_��IX4@m�"�N�!?�W9��+�@�g�y�ٿX}���@bH���4@�xWt�!?S]�Gp+�@�g�y�ٿX}���@bH���4@�xWt�!?S]�Gp+�@�g�y�ٿX}���@bH���4@�xWt�!?S]�Gp+�@�R�q&�ٿ������@$��}�4@}���!?���8�+�@�R�q&�ٿ������@$��}�4@}���!?���8�+�@�R�q&�ٿ������@$��}�4@}���!?���8�+�@�R�q&�ٿ������@$��}�4@}���!?���8�+�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@��F��ٿ�DrF��@��  4@��-��!?MJ�M�*�@N��:�ٿ=�J���@�[9�4@M��j�!?��֓+�@N��:�ٿ=�J���@�[9�4@M��j�!?��֓+�@N��:�ٿ=�J���@�[9�4@M��j�!?��֓+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@��`rt�ٿ[:����@i���4@��KӨ�!?$Z/l+�@�����ٿ����@]SuSc4@�nGM��!?�9B��+�@�����ٿ����@]SuSc4@�nGM��!?�9B��+�@�����ٿ����@]SuSc4@�nGM��!?�9B��+�@�����ٿ����@]SuSc4@�nGM��!?�9B��+�@�����ٿ����@]SuSc4@�nGM��!?�9B��+�@{
K��ٿ������@�gh��4@�<�G��!?����+�@{
K��ٿ������@�gh��4@�<�G��!?����+�@)��M$�ٿ�eѾ��@�֝z�4@Aa+ 7�!?x$�0,�@?�n���ٿ�7Ň�@��x4@��E� �!?�0'�&,�@?�n���ٿ�7Ň�@��x4@��E� �!?�0'�&,�@?�n���ٿ�7Ň�@��x4@��E� �!?�0'�&,�@$u���ٿ��{���@��0 4@B����!?�i��+�@$u���ٿ��{���@��0 4@B����!?�i��+�@$u���ٿ��{���@��0 4@B����!?�i��+�@�p��ٿ�؏|���@j5�[�	4@
�tK�!?`�7^�,�@�p��ٿ�؏|���@j5�[�	4@
�tK�!?`�7^�,�@�p��ٿ�؏|���@j5�[�	4@
�tK�!?`�7^�,�@�p��ٿ�؏|���@j5�[�	4@
�tK�!?`�7^�,�@�p��ٿ�؏|���@j5�[�	4@
�tK�!?`�7^�,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@y�J�ٿ�\phχ�@p*��?4@B��.P�!?�ӴE
,�@K10g�ٿ�ړ��@D�g9�
4@ΣAf��!?�%��o,�@K10g�ٿ�ړ��@D�g9�
4@ΣAf��!?�%��o,�@���ϐٿ-S�|��@�0)4@Ѕ��!?����,�@���ϐٿ-S�|��@�0)4@Ѕ��!?����,�@���ϐٿ-S�|��@�0)4@Ѕ��!?����,�@���ϐٿ-S�|��@�0)4@Ѕ��!?����,�@�q@�ٿ�p�}��@���vU4@%{��!?M�!��+�@�q@�ٿ�p�}��@���vU4@%{��!?M�!��+�@�q@�ٿ�p�}��@���vU4@%{��!?M�!��+�@��s��ٿ��鸈�@���*�4@h^6ΐ!?"8�y)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@,�����ٿ��̈�@�/��� 4@	��\�!?���e)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@��(��ٿ��<����@���$4@e��ې!?���)�@�W��͊ٿ]S�y��@�e` � 4@�f����!?�[B\*�@�W��͊ٿ]S�y��@�e` � 4@�f����!?�[B\*�@�0�ٿ�f'��@�y|��3@�	=Ð!?#�@js(�@�0�ٿ�f'��@�y|��3@�	=Ð!?#�@js(�@�=x쀓ٿbG����@�q�}[4@��Ґ!?���U�+�@�=x쀓ٿbG����@�q�}[4@��Ґ!?���U�+�@�=x쀓ٿbG����@�q�}[4@��Ґ!?���U�+�@�=x쀓ٿbG����@�q�}[4@��Ґ!?���U�+�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@���\�ٿ�Ժ��@�4@��Dc�!?���RQ,�@O:^�܍ٿ�ts+��@���	4@϶D�C�!?  ��-�@_��F�ٿ���IІ�@�Wgծ
4@�ᑭ �!?��
`.�@:R�㛁ٿ&�h�L��@�
�^
4@'Y*�R�!?��8�,�@l�	��ٿ�Qzb��@���v4@d�*�W�!?lM��,�@l�	��ٿ�Qzb��@���v4@d�*�W�!?lM��,�@l�	��ٿ�Qzb��@���v4@d�*�W�!?lM��,�@l�	��ٿ�Qzb��@���v4@d�*�W�!?lM��,�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@|��Ds�ٿ1�2����@��il(4@bO ې!?@���)�@�1����ٿ�nB����@-��4@�� �!?zj��A,�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�N��>�ٿ�FU��@��F�[4@Q��㔐!?�x���*�@�:�)�ٿ�/�:��@���{�4@Wd���!?ӋN��(�@��&�ٿV�h0K��@�u�0A 4@��j��!?�m���%�@'DQ3�~ٿ)c�:��@����4@�JO�!?0�)&�@'DQ3�~ٿ)c�:��@����4@�JO�!?0�)&�@'DQ3�~ٿ)c�:��@����4@�JO�!?0�)&�@'DQ3�~ٿ)c�:��@����4@�JO�!?0�)&�@'DQ3�~ٿ)c�:��@����4@�JO�!?0�)&�@��|ÁٿN�/����@�9F�N
4@��uI��!?�
(�@��|ÁٿN�/����@�9F�N
4@��uI��!?�
(�@��|ÁٿN�/����@�9F�N
4@��uI��!?�
(�@���Ezٿ]��J���@����4@��q�!?_��!#�@���Ezٿ]��J���@����4@��q�!?_��!#�@���Ezٿ]��J���@����4@��q�!?_��!#�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@j{�^6�ٿ�X.1ϊ�@�5a��	4@� ?���!?�\�b[%�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@E�R�N�ٿY�Ň�@���&�4@&�i�!?]m{�,�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@A�9���ٿ�xf9���@�^�A4@S��\N�!?����*�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@�wY��ٿ՞bN���@��]�\4@7:�0�!?v(�w'�@."u{�~ٿ8�D)���@g�Ϗ�4@�t��|�!?�x�C�&�@."u{�~ٿ8�D)���@g�Ϗ�4@�t��|�!?�x�C�&�@."u{�~ٿ8�D)���@g�Ϗ�4@�t��|�!?�x�C�&�@�~n%�ٿc�Fˌ�@7)��4@�mlW��!?L�~�� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@fđ�B�ٿ��+���@�ʧ�i	4@Զ����!?��^� �@$��ٿG�k>���@'"Xe�4@�E�ᯐ!?�P��9!�@$��ٿG�k>���@'"Xe�4@�E�ᯐ!?�P��9!�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@�D��w�ٿEp�0V��@}hc�4@-�����!?]Nz�1�@x9E�ٿe�~x��@B���d4@��>��!?����K�@x9E�ٿe�~x��@B���d4@��>��!?����K�@a��5�{ٿ[5�.#��@l4@
ٶꀐ!?�f�,�@9���)|ٿ�������@�&D� 4@��&m�!?�<B�	�@K,����ٿ*-`D��@"7���4@a�!?;����@K,����ٿ*-`D��@"7���4@a�!?;����@K,����ٿ*-`D��@"7���4@a�!?;����@K,����ٿ*-`D��@"7���4@a�!?;����@����xٿ1���>��@<W�4@Z��ݐ!?�0[��@����xٿ1���>��@<W�4@Z��ݐ!?�0[��@����xٿ1���>��@<W�4@Z��ݐ!?�0[��@����xٿ1���>��@<W�4@Z��ݐ!?�0[��@����xٿ1���>��@<W�4@Z��ݐ!?�0[��@aϝ(��ٿ:���ˋ�@ܗ�4@��2�!?Ho1��#�@aϝ(��ٿ:���ˋ�@ܗ�4@��2�!?Ho1��#�@aϝ(��ٿ:���ˋ�@ܗ�4@��2�!?Ho1��#�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@�S�`��ٿ�v��͌�@��p�4@[����!?�Ĳ�!�@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@��}�xٿy�e�֢�@�_���4@}ڊא!?��?i��@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@,Rl�,�ٿ�<��@�4#P�4@���K�!?S'�I���@���-w�ٿ��9���@�����
4@[^���!?�u���@���-w�ٿ��9���@�����
4@[^���!?�u���@q!��M�ٿ��no��@|
���4@ef�H�!?�c)s��@q!��M�ٿ��no��@|
���4@ef�H�!?�c)s��@q!��M�ٿ��no��@|
���4@ef�H�!?�c)s��@���\�|ٿ�<f���@ �
t�4@p�xА!?{s�E��@���\�|ٿ�<f���@ �
t�4@p�xА!?{s�E��@���\�|ٿ�<f���@ �
t�4@p�xА!?{s�E��@���\�|ٿ�<f���@ �
t�4@p�xА!?{s�E��@Z� ��ٿa Q��@���4@��+�H�!?l�AL��@Z� ��ٿa Q��@���4@��+�H�!?l�AL��@Z� ��ٿa Q��@���4@��+�H�!?l�AL��@ѡvI�ٿI�'V���@ȗh�%4@��qyŐ!?��;��	�@ѡvI�ٿI�'V���@ȗh�%4@��qyŐ!?��;��	�@ѡvI�ٿI�'V���@ȗh�%4@��qyŐ!?��;��	�@�)�$��ٿ�fe���@*:�\T4@���:�!?��Zz���@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@E=l�Ɍٿq`xʕ�@��Խ4@ۻa��!?Q՚�@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�p#!b�ٿ�D���@�r#�#4@���!?�L7����@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@�e�뇋ٿ'�di���@�(�C4@�~t�/�!?���(�@��r1=�ٿ9���O��@L�x<4@�I��M�!?��sѠ�@��r1=�ٿ9���O��@L�x<4@�I��M�!?��sѠ�@4U�O-�ٿN/��m��@Qj��4@	}�"�!? _�����@�� �ٿ�E�&���@�_��� 4@ݒ�ҟ�!?����1�@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@R[ۄ܏ٿDFϔ��@����4@\�ܔ�!?�ռ��@OK]N1{ٿ�����@���c(4@���i��!?�b�����@OK]N1{ٿ�����@���c(4@���i��!?�b�����@ X,PU{ٿΙŏ��@�	�4@�W�Zِ!?hM����@ X,PU{ٿΙŏ��@�	�4@�W�Zِ!?hM����@ X,PU{ٿΙŏ��@�	�4@�W�Zِ!?hM����@ X,PU{ٿΙŏ��@�	�4@�W�Zِ!?hM����@�T��ٿ/_�zǩ�@m�z84@�K�~&�!?
MJ��@�T��ٿ/_�zǩ�@m�z84@�K�~&�!?
MJ��@�T��ٿ/_�zǩ�@m�z84@�K�~&�!?
MJ��@�T��ٿ/_�zǩ�@m�z84@�K�~&�!?
MJ��@~��{~ٿ���L]��@
v��4@7�O�Ր!?��x���@�.f�ٿi'J���@����4@ƍ���!?�?�u��@�.f�ٿi'J���@����4@ƍ���!?�?�u��@��76�ٿ���@�?a4@�wŐ!?�"C��@��76�ٿ���@�?a4@�wŐ!?�"C��@��76�ٿ���@�?a4@�wŐ!?�"C��@��76�ٿ���@�?a4@�wŐ!?�"C��@��76�ٿ���@�?a4@�wŐ!?�"C��@"�5v�~ٿ{��,���@�s�NH4@%��zܐ!?F�0�/��@"�5v�~ٿ{��,���@�s�NH4@%��zܐ!?F�0�/��@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@x�<�ٿɾ��1��@�g��k4@~x͙�!?G�)!���@�Y����ٿN?�0��@/�Ś�4@�'���!?S(o��@�Y����ٿN?�0��@/�Ś�4@�'���!?S(o��@�Y����ٿN?�0��@/�Ś�4@�'���!?S(o��@|G�)�ٿ�pm%��@B�/ 4@���!?�Q:���@|G�)�ٿ�pm%��@B�/ 4@���!?�Q:���@l�Ɖٿ+�<m��@}nFP�4@�\���!?*�+���@l�Ɖٿ+�<m��@}nFP�4@�\���!?*�+���@l�Ɖٿ+�<m��@}nFP�4@�\���!?*�+���@�QZ8\�ٿv�ē��@���94@VT[�D�!?����@����ٿ���e¨�@p��4@�:F~�!?�)����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@`\d��ٿ�*�1���@�+���4@����!?��n����@�Ȭ�[�ٿ�ٛ7��@�$�ȗ4@�K��!?�S},���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@�X�ٿ(U|��@�m�O�4@�ЮH�!?4;�J���@��Ғ�zٿ9����@��
��4@*�_���!?�8)�]�@k���_�ٿ�\R���@]��n�4@߫2���!?xvlG]P�@k���_�ٿ�\R���@]��n�4@߫2���!?xvlG]P�@�X��ٿa�@Q��@�w�j!4@����!?��U��z�@�X��ٿa�@Q��@�w�j!4@����!?��U��z�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@�S�_z�ٿ07�((��@��ngH4@'�uː!?es<X�`�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@����}ٿǡ�ɬ��@�*Ai94@;�O���!?����^�@1�N�
�ٿ���i���@G��`4@��ڒ�!?E9���c�@1�N�
�ٿ���i���@G��`4@��ڒ�!?E9���c�@1�N�
�ٿ���i���@G��`4@��ڒ�!?E9���c�@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@!���E~ٿ٧�aD�@M���y4@��Ő!?�C�l��@�#癄ٿp����@�T��4@�2�>Ґ!?�8b��a�@�#癄ٿp����@�T��4@�2�>Ґ!?�8b��a�@�#癄ٿp����@�T��4@�2�>Ґ!?�8b��a�@�#癄ٿp����@�T��4@�2�>Ґ!?�8b��a�@y=���ٿ+����?�@�G�c�4@�B�Đ!??�΂d��@��௅ٿ�!n,A!�@@~�Y�4@0����!?=��Ά��@��௅ٿ�!n,A!�@@~�Y�4@0����!?=��Ά��@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@N�i��ٿIi�)���@��6k�
4@f��А!?^�CU�9�@(| ���ٿ4��e�@a̙!�4@	-�8�!?}c!�[�@(| ���ٿ4��e�@a̙!�4@	-�8�!?}c!�[�@(| ���ٿ4��e�@a̙!�4@	-�8�!?}c!�[�@(| ���ٿ4��e�@a̙!�4@	-�8�!?}c!�[�@(| ���ٿ4��e�@a̙!�4@	-�8�!?}c!�[�@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@[]��~ٿ�^9�q�@QVEE4@[6���!?BfB�.��@Ϙ�>��ٿm�D���@FB�h4@y���!?7����@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@4�Р.�ٿ,����@�oA�[4@V16S �!?���j���@��gbZ�ٿ�{�N�@di�v	4@R��+�!?~E$���@��gbZ�ٿ�{�N�@di�v	4@R��+�!?~E$���@��0�zٿ�MV�A�@��[6�4@R8���!?�#GK��@��0�zٿ�MV�A�@��[6�4@R8���!?�#GK��@��0�zٿ�MV�A�@��[6�4@R8���!?�#GK��@��0�zٿ�MV�A�@��[6�4@R8���!?�#GK��@��0�zٿ�MV�A�@��[6�4@R8���!?�#GK��@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@�ugT{ٿ6%xL�@��Д4@�9�¹�!?��G]���@p%!Ńٿ�<�46��@��_�4@5h���!?�)��u�@�(,l-vٿ�-O�@E���x4@�&�ӹ�!?�^�Z�@�(,l-vٿ�-O�@E���x4@�&�ӹ�!?�^�Z�@�(,l-vٿ�-O�@E���x4@�&�ӹ�!?�^�Z�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@t�-�yٿ��x2�g�@V�Nt�4@���!?���#�B�@E��qvٿ�1'˵7�@�7���4@(u~ΐ!?�?��
��@E��qvٿ�1'˵7�@�7���4@(u~ΐ!?�?��
��@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@}��!Mٿ~�;)G��@Q��x�
4@���t�!?�r��+�@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�en��ٿo��,��@[>�Q�4@1s�9�!?�}3-���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@�c03+�ٿ�v�����@ut�O�4@,��/�!?�u�q���@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@%k�ٿj��D���@�kaO	4@�HO��!?j���؞�@!�ö��ٿ��1z��@��[b4@�ZY��!?��K_�Q�@�w�ٿy\�T���@�G=1�4@���ᵐ!?�Ņ��@�w�ٿy\�T���@�G=1�4@���ᵐ!?�Ņ��@�w�ٿy\�T���@�G=1�4@���ᵐ!?�Ņ��@N.Y��ٿ|MՁ��@���9�4@0�Z��!?��T�b��@N.Y��ٿ|MՁ��@���9�4@0�Z��!?��T�b��@�-9 �ٿ�]�΄@�@��bc/
4@��!��!?[D�����@�-9 �ٿ�]�΄@�@��bc/
4@��!��!?[D�����@�)��ٿE��m��@��-4@^k-�ː!?W�{�7�@�)��ٿE��m��@��-4@^k-�ː!?W�{�7�@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��gw��ٿGR�u%;�@k��4@F\\pא!?�#�d>��@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@��S�Ѕٿ��J}}\�@����d4@�n�XƐ!?�7�Z�@:�=O�ٿah��[\�@�'��a4@g	mː!?̅�,Z�@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@���)�ٿ�3�*�@/{
7p4@�Ŏ��!?/�cH ��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@��T(֎ٿ�{�t�-�@9�"��4@�´�!?�"R��@v_��4�ٿ�O�� ��@lq٢74@�r�X��!?A��S]�@v_��4�ٿ�O�� ��@lq٢74@�r�X��!?A��S]�@v_��4�ٿ�O�� ��@lq٢74@�r�X��!?A��S]�@v_��4�ٿ�O�� ��@lq٢74@�r�X��!?A��S]�@v_��4�ٿ�O�� ��@lq٢74@�r�X��!?A��S]�@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@��WIՄٿ�kc���@��z4@�T����!?!�����@E�C�ٿr��5���@Y�)94@�L)B��!?�z�w�U�@E�C�ٿr��5���@Y�)94@�L)B��!?�z�w�U�@d8p<�ٿ}&�)�@c��$4@�e�d�!?,���*��@d8p<�ٿ}&�)�@c��$4@�e�d�!?,���*��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@��8E��ٿ��`�5�@�dn�4@�{�V��!?�=?<��@�XC�(�ٿ���@�#54@�il!?>��Ti�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@%��D�ٿ덽����@�Z&��4@���=��!?�G�]q&�@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@̙�څٿ���=�@v+��4@�^��!?�ȏ���@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@@t�l�ٿ��KR\�@h_���4@-tߦ��!?��f��X�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@�)�*�ٿ���y�]�@��U�	4@l�RE��!?��p U�@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@`C4�݆ٿ��Z�K:�@�R�Sz4@i�`�ϐ!?j��U���@�x"�>�ٿ��L[�=�@��.�L4@Y�Y�Ր!?���Ӛ�@�x"�>�ٿ��L[�=�@��.�L4@Y�Y�Ր!?���Ӛ�@�щ�ٿ���:�@�ϱ��	4@�R���!?������@�K���ٿ�~�v���@�Ɨ<H4@�V�0ɐ!?���1Fp�@�K���ٿ�~�v���@�Ɨ<H4@�V�0ɐ!?���1Fp�@�K���ٿ�~�v���@�Ɨ<H4@�V�0ɐ!?���1Fp�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@d�$J<�ٿ��fD���@�?���4@�{�蠐!?c�]`ln�@S��f�ٿ�xM
�i�@E��(4@(}�r��!?W��D�1�@S��f�ٿ�xM
�i�@E��(4@(}�r��!?W��D�1�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@��&W�ٿ@-��89�@��J��4@�F�!?ϣ�Kܙ�@؃ï�ٿS��G��@u��O4@��nTӐ!?ϩG��@؃ï�ٿS��G��@u��O4@��nTӐ!?ϩG��@	_�@�ٿ��/�]��@o4�	4@�.����!?^�Ř�@!Ѐ���ٿ|c~���@J�҇4@�3�zq�!?ə�F�6�@!Ѐ���ٿ|c~���@J�҇4@�3�zq�!?ə�F�6�@!Ѐ���ٿ|c~���@J�҇4@�3�zq�!?ə�F�6�@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�df��ٿ6��$�"�@���4@�<��x�!?�+yG���@�ќ�ٿ�j���G�@�C#�4@8	s��!?>�6�߅�@�ќ�ٿ�j���G�@�C#�4@8	s��!?>�6�߅�@�B���ٿ�m	J�3�@q3{�t4@�So��!?����ܩ�@�B���ٿ�m	J�3�@q3{�t4@�So��!?����ܩ�@�B���ٿ�m	J�3�@q3{�t4@�So��!?����ܩ�@p�6���ٿ;#e�5(�@Q�s4@����&�!?7|�! ��@p�6���ٿ;#e�5(�@Q�s4@����&�!?7|�! ��@EC��^�ٿ�vd�cG�@���84@����\�!?�[���@EC��^�ٿ�vd�cG�@���84@����\�!?�[���@EC��^�ٿ�vd�cG�@���84@����\�!?�[���@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@+=r��ٿT�ƃ�@)�֐4@@�!�E�!?�d����@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@�^G�ٿ9Pa�#�@�Vd�4@#%��Ґ!?�������@��E?'�ٿ���3H�@��F��4@|lx*��!?U�f���@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@]}o�-�ٿ���@ύ��4@�a	���!?�7s
�
�@I����ٿ<u�9;��@�ڬa4@�}��4�!?U�
q.�@R���ٿ� ��Sb�@蚇	4@Ǡ1w
�!?�<��Y�@R���ٿ� ��Sb�@蚇	4@Ǡ1w
�!?�<��Y�@R���ٿ� ��Sb�@蚇	4@Ǡ1w
�!?�<��Y�@R���ٿ� ��Sb�@蚇	4@Ǡ1w
�!?�<��Y�@3�x̉ٿ�NTN{�@�� E�4@��r�!?�eS��@3�x̉ٿ�NTN{�@�� E�4@��r�!?�eS��@3�x̉ٿ�NTN{�@�� E�4@��r�!?�eS��@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@ħ����ٿ��U�,��@r���4@a�>I��!?ȝ2��F�@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@���C��ٿ9>�Wo>�@+�M�4@Jx����!?��-EZ��@ۡ]W��ٿ�:����@^�xC}4@6cX�͐!?��F�g�@��k��ٿл����@4�z�z4@R����!?8�O�n*�@��k��ٿл����@4�z�z4@R����!?8�O�n*�@��k��ٿл����@4�z�z4@R����!?8�O�n*�@��k��ٿл����@4�z�z4@R����!?8�O�n*�@��k��ٿл����@4�z�z4@R����!?8�O�n*�@ڍ�Oٌٿ�~;���@Yۼ�4@����!?�rĻ�7�@ڍ�Oٌٿ�~;���@Yۼ�4@����!?�rĻ�7�@ڍ�Oٌٿ�~;���@Yۼ�4@����!?�rĻ�7�@ڍ�Oٌٿ�~;���@Yۼ�4@����!?�rĻ�7�@#;̱�ٿjh����@���U4@=��^��!?b�q��@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@cq�n)�ٿ
#x��@VU-4@nӫ�ΐ!?)�s�09�@�]C�ٿ�Q��}��@��,V�4@�&R���!?�,h�G��@�&��ٿp��O���@����r4@��|�Ӑ!?�"/f��@��!3�ٿ�yw����@)�|�4@�ٖǐ!?B\�r�O�@ZL���ٿ��[}�3�@�v�͌4@B�ז�!?���ީ�@�с�ٿ@��e8�@�& GH4@2����!?�9Pɜ�@�с�ٿ@��e8�@�& GH4@2����!?�9Pɜ�@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@H�*�ٿMڌ� �@E�F�44@~���!?�{�` �@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�M�C�ٿ�^̑X��@PӦ�54@-�P�!?�ǌ�n1�@�R���ٿD���,�@5�]�4@��!N��!?�ZM���@,��ٿr4�0��@���`4@�b����!?d]h����@,��ٿr4�0��@���`4@�b����!?d]h����@,��ٿr4�0��@���`4@�b����!?d]h����@,��ٿr4�0��@���`4@�b����!?d]h����@,��ٿr4�0��@���`4@�b����!?d]h����@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@x�޴��ٿ'�	����@�Qn�4@�7����!?� ��i�@G�i���ٿѺ?�8�@c�W�4@�>���!?Ÿ��_��@�SR�x{ٿ�e>$�@��}�4@�c/[��!?�Aۨ��@�SR�x{ٿ�e>$�@��}�4@�c/[��!?�Aۨ��@I���{ٿ7�z�R�@���`4	4@�6>��!?t�Fr�@��eHٿ����*�@p���	4@�o^�!?9&�����@,��ŷ~ٿ����2�@�SE��4@3t�ӆ�!?r�Z���@,��ŷ~ٿ����2�@�SE��4@3t�ӆ�!?r�Z���@,��ŷ~ٿ����2�@�SE��4@3t�ӆ�!?r�Z���@,��ŷ~ٿ����2�@�SE��4@3t�ӆ�!?r�Z���@��X���ٿX��J`��@�55<�	4@k/q�q�!?��&l�@��X���ٿX��J`��@�55<�	4@k/q�q�!?��&l�@��X���ٿX��J`��@�55<�	4@k/q�q�!?��&l�@��X���ٿX��J`��@�55<�	4@k/q�q�!?��&l�@���ٿ������@f���4@�ŶT��!?E��ӧx�@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@���V��ٿ\�`!��@�<��4@p*4Gf�!?'����@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@7H[争ٿ�����$�@��F4@tB��s�!?�+<[���@�ܜ�ˌٿ�w��S*�@i�1$^4@�2tv�!?�X�LB��@���,�ٿ�\zi�@�s�h�4@��v�|�!?w<C�@���,�ٿ�\zi�@�s�h�4@��v�|�!?w<C�@��g�ٿ�����@�c_D4@�缑�!?{a'�@��@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@��˂�ٿ��$�5��@aT��4@r�!?�����@7�"ωٿ󦈜���@�L��,
4@/��@��!?'(:����@7�"ωٿ󦈜���@�L��,
4@/��@��!?'(:����@7�"ωٿ󦈜���@�L��,
4@/��@��!?'(:����@7�"ωٿ󦈜���@�L��,
4@/��@��!?'(:����@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@��P��ٿA��#[�@�Wт�4@!��_ݐ!?=V�ir�@g�y��ٿ;��*?T�@���*4@�Q)C�!?�����@���zٿ�^38��@a�� m4@M�s���!?v��� "�@�N���{ٿ�"�v/�@��H�4@�ps�!?2�a��@�N���{ٿ�"�v/�@��H�4@�ps�!?2�a��@�N���{ٿ�"�v/�@��H�4@�ps�!?2�a��@����q�ٿ�|�-�@�@u�4@D�i��!?]���&�@����q�ٿ�|�-�@�@u�4@D�i��!?]���&�@]��فٿ��0�$'�@��Bx0	4@�]��!?M�x�g��@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@�Q#�ٿ�y��-�@�[%4@�,3�!?�>�Q���@<#��v�ٿ@8�b��@�%U)N4@�>��!?��O�QI�@<#��v�ٿ@8�b��@�%U)N4@�>��!?��O�QI�@<#��v�ٿ@8�b��@�%U)N4@�>��!?��O�QI�@%,���ٿ��6:��@sðO	4@p81���!?ɪː��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@;�Q��ٿ��t��@�sQD4@���!�!?��Oap��@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@���,\�ٿ���uQ�@�����4@�Ʈ&��!?�Z�E�{�@z�V�Ȇٿ� ,�[F�@/>���4@���Њ�!?��}Ã�@z�V�Ȇٿ� ,�[F�@/>���4@���Њ�!?��}Ã�@z�V�Ȇٿ� ,�[F�@/>���4@���Њ�!?��}Ã�@�a�]*�ٿ�m � �@S��4	4@�����!?P��� �@�a�]*�ٿ�m � �@S��4	4@�����!?P��� �@�a�]*�ٿ�m � �@S��4	4@�����!?P��� �@�a�]*�ٿ�m � �@S��4	4@�����!?P��� �@�1�Eލٿ3��W���@�WV�4@_\���!?Aa��$��@��|�ٿ��`����@v��`;
4@_P �!?�ի:w�@��|�ٿ��`����@v��`;
4@_P �!?�ի:w�@��|�ٿ��`����@v��`;
4@_P �!?�ի:w�@��|�ٿ��`����@v��`;
4@_P �!?�ի:w�@��|�ٿ��`����@v��`;
4@_P �!?�ի:w�@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@�F5,�ٿ�}�.��@;���4@ gԚ�!?����?��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@c�d�ٿif"c��@�ƺ�4@oR�a��!?o�	Ŝ��@
�*\�ٿ�~Im�@AA0	4@���!?SpD�p�@
�*\�ٿ�~Im�@AA0	4@���!?SpD�p�@�l��ٿ1Y���5�@1ÄP�4@R&��!?%��ݽ��@�l��ٿ1Y���5�@1ÄP�4@R&��!?%��ݽ��@z���ٿnB�a��@�}�-4@�m����!?,[l��o�@z���ٿnB�a��@�}�-4@�m����!?,[l��o�@z���ٿnB�a��@�}�-4@�m����!?,[l��o�@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@�}z�ٿ��P��]�@:��4@J�+�!?�]�k8��@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@���
Ȅٿ;�6%��@���v4@��K�!?p��W�@�ڗ�ԉٿ�v����@ ��4@�2)���!?�	����@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@Hy���ٿa`��@� �4@l�߸�!?�Ө���@�<�rސٿ$J��XI�@�H��4@�;�zI�!?��dMn�@�<�rސٿ$J��XI�@�H��4@�;�zI�!?��dMn�@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@�?��ԁٿn�G�@��cn4@��Jѐ!?7+!����@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@};��уٿ��4�@�z�{4@w���!?]�Tc_$�@�q�ℂٿ����I�@�"�>�4@�-�h��!?����ړ�@ՠsA�ٿ����2�@����
4@��� Ɛ!?!�]����@ՠsA�ٿ����2�@����
4@��� Ɛ!?!�]����@ՠsA�ٿ����2�@����
4@��� Ɛ!?!�]����@ՠsA�ٿ����2�@����
4@��� Ɛ!?!�]����@2�mj�ٿE�.�VP�@@2�8�4@@�S4�!?b�Sq�u�@2�mj�ٿE�.�VP�@@2�8�4@@�S4�!?b�Sq�u�@2�mj�ٿE�.�VP�@@2�8�4@@�S4�!?b�Sq�u�@2�mj�ٿE�.�VP�@@2�8�4@@�S4�!?b�Sq�u�@$]5�ٿNX7)d�@�}�WS4@�,��!?��q�1�@$]5�ٿNX7)d�@�}�WS4@�,��!?��q�1�@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@�90<�ٿ{,��*�@��W�4@sD��!?��>���@[C)Jٿ�FN�o�@�N}Q�4@dG��!?�17��$�@�{O�وٿ�3��+�@,��	;	4@7�i��!?y�����@���k�ٿ�W��,�@���|�4@�{ݼ�!?gZ8ue��@���k�ٿ�W��,�@���|�4@�{ݼ�!?gZ8ue��@���k�ٿ�W��,�@���|�4@�{ݼ�!?gZ8ue��@���k�ٿ�W��,�@���|�4@�{ݼ�!?gZ8ue��@��'��ٿ����F�@�0I�<4@����!?Н��U��@��'��ٿ����F�@�0I�<4@����!?Н��U��@��'��ٿ����F�@�0I�<4@����!?Н��U��@��'��ٿ����F�@�0I�<4@����!?Н��U��@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@,��	
�ٿX��	�@v�ݖ4@Xy,Wϐ!?y_��*�@��.Ԇٿ�_��?�@��,4@K��!?!�����@��.Ԇٿ�_��?�@��,4@K��!?!�����@1���ٿ�����a�@�y�F4@�5�Ð!?��9X�@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@q�MeY�ٿ@y�TN!�@9����4@�t(�	�!?�*����@= �z�ٿ*�2E���@X:�4@�3u�!?��,.c�@= �z�ٿ*�2E���@X:�4@�3u�!?��,.c�@= �z�ٿ*�2E���@X:�4@�3u�!?��,.c�@z�����ٿ�P�aN��@��M�H4@��Cc�!?oޤ	�%�@��`��ٿ���A�@_n��4@��
n �!?l�����@��`��ٿ���A�@_n��4@��
n �!?l�����@��`��ٿ���A�@_n��4@��
n �!?l�����@^g�ٿn���I�@N._R4@(�t@Ր!?�/wW�@^g�ٿn���I�@N._R4@(�t@Ր!?�/wW�@^g�ٿn���I�@N._R4@(�t@Ր!?�/wW�@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@Pt;���ٿ��K��@~;�q
4@�Rn�!?>?����@_=����ٿ�B�9S�@,�$T4@�2����!?5�aĮk�@_=����ٿ�B�9S�@,�$T4@�2����!?5�aĮk�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@~@��>�ٿJvp_�@n�bj4@��uB��!?-N�<�@ܛf�&�ٿY���U��@���:	4@j�#,�!?�ǹZh�@ܛf�&�ٿY���U��@���:	4@j�#,�!?�ǹZh�@��,�Ռٿ��&����@�J0	4@�6���!?�!S�n�@��,�Ռٿ��&����@�J0	4@�6���!?�!S�n�@#qt:Çٿ��G�<�@��\�
4@,s�+.�!?wT����@�2q0�ٿ)�,�\B�@+�*4@6rs��!?ښm˪�@�2q0�ٿ)�,�\B�@+�*4@6rs��!?ښm˪�@�2q0�ٿ)�,�\B�@+�*4@6rs��!?ښm˪�@�2q0�ٿ)�,�\B�@+�*4@6rs��!?ښm˪�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@�_��n�ٿ�x�7p�@m煈4@��P �!?�6��M�@{�"��ٿn����G�@і�4@�[]x��!?"����{�@���ֱ�ٿ���1�M�@�ll�T4@����}�!?S����_�@�V���ٿO�m��O�@U�0Z�4@p�H��!?�R��I�@Zr�*!�ٿw|��@+#�*4@0joq��!?��c4���@Zr�*!�ٿw|��@+#�*4@0joq��!?��c4���@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@Fc4̈ٿi+ʬ�5�@���%4@���!?^"Q��@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@{�껋ٿ�~�^�"�@J��0�4@�^�S��!?iS����@�Lj���ٿ^��r$�@_P.C4@���U��!?L�|ZO�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@vDH1<�ٿ��)�V^�@�:�7z4@��E��!?g�@�Z�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@ٜ�ꨆٿ�po_���@".�t�4@��[y�!?�Pصn1�@9M�16�ٿZ��N�@��E�L4@DƬ��!?���x���@9M�16�ٿZ��N�@��E�L4@DƬ��!?���x���@9M�16�ٿZ��N�@��E�L4@DƬ��!?���x���@9M�16�ٿZ��N�@��E�L4@DƬ��!?���x���@9M�16�ٿZ��N�@��E�L4@DƬ��!?���x���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@�}��ٿ��]Ey��@����4@w�*:j�!?y�i���@O	��`�ٿi6 U��@m���*4@���^��!?K������@O	��`�ٿi6 U��@m���*4@���^��!?K������@O	��`�ٿi6 U��@m���*4@���^��!?K������@O	��`�ٿi6 U��@m���*4@���^��!?K������@O	��`�ٿi6 U��@m���*4@���^��!?K������@O	��`�ٿi6 U��@m���*4@���^��!?K������@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@�/w�}ٿ%#����@苑l 4@���{͐!?H�f���@2u</�ٿ�c�ÛA�@o3�&"4@lAF-�!?,#l܎o�@���a)�ٿ9\K��J�@hH�4@���ؐ!?JW��H�@+l��R�ٿ���3� �@���4@ew��!?���4��@+l��R�ٿ���3� �@���4@ew��!?���4��@+l��R�ٿ���3� �@���4@ew��!?���4��@+l��R�ٿ���3� �@���4@ew��!?���4��@��'�܈ٿ������@Y��9#
4@Rɝ��!?��h�'�@��'�܈ٿ������@Y��9#
4@Rɝ��!?��h�'�@���W��ٿ�,����@l�0��
4@h	sJ��!?��\>uQ�@���W��ٿ�,����@l�0��
4@h	sJ��!?��\>uQ�@���W��ٿ�,����@l�0��
4@h	sJ��!?��\>uQ�@���W��ٿ�,����@l�0��
4@h	sJ��!?��\>uQ�@Uax~#�ٿa�lG(;�@4O�{/
4@�+cEА!?�����Y�@�9�ٿ��P���@���Y4@F����!?~��K"~�@�9�ٿ��P���@���Y4@F����!?~��K"~�@�9�ٿ��P���@���Y4@F����!?~��K"~�@�9�ٿ��P���@���Y4@F����!?~��K"~�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��̘M�ٿ�&��%�@'�>B�4@�0��!?��pJH�@��z_��ٿ;����@q)�4@c~�!?��Z�*�@��z_��ٿ;����@q)�4@c~�!?��Z�*�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@rT J�ٿpR�n�@��;�4@d����!?XW�V�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D\���ٿ�U\���@>.Ml��3@��"ۖ�!?<�J�3!�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@D�C��ٿ����S��@t��4@���e�!?�2Y�Y�@|[�$��ٿxi�>��@`���4@�"�m�!?i f
I"�@|[�$��ٿxi�>��@`���4@�"�m�!?i f
I"�@|[�$��ٿxi�>��@`���4@�"�m�!?i f
I"�@|[�$��ٿxi�>��@`���4@�"�m�!?i f
I"�@|[�$��ٿxi�>��@`���4@�"�m�!?i f
I"�@?;<m��ٿ�{ٴV��@[X��{4@~@�:�!?��}���@?;<m��ٿ�{ٴV��@[X��{4@~@�:�!?��}���@?;<m��ٿ�{ٴV��@[X��{4@~@�:�!?��}���@?;<m��ٿ�{ٴV��@[X��{4@~@�:�!?��}���@���@��ٿ+Ok,")�@xb��4@R��_��!?W�);J��@���@��ٿ+Ok,")�@xb��4@R��_��!?W�);J��@kA��'�ٿ��Ob�@����4@,C&!ܐ!?�r�n�@kA��'�ٿ��Ob�@����4@,C&!ܐ!?�r�n�@[�ݴ!�ٿ�	�(%g�@�i�H 4@�F�hŐ!?�iZ��@[�ݴ!�ٿ�	�(%g�@�i�H 4@�F�hŐ!?�iZ��@[�ݴ!�ٿ�	�(%g�@�i�H 4@�F�hŐ!?�iZ��@{�R�E�ٿ��Kֆ`�@@�W s4@�[E��!?�mw���@�Q��ٿ�f
��@����4@�����!?���Q�f�@�Q��ٿ�f
��@����4@�����!?���Q�f�@����ٿX�����@F��4@/m�q�!?ݗ�.4�@����ٿX�����@F��4@/m�q�!?ݗ�.4�@����ٿX�����@F��4@/m�q�!?ݗ�.4�@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@~�p!�ٿ/!pZ���@�r�d��3@_tH��!?DS?���@��_F2�ٿn
y����@!'��*4@�}�ߐ!?J0B��_�@��_F2�ٿn
y����@!'��*4@�}�ߐ!?J0B��_�@��_F2�ٿn
y����@!'��*4@�}�ߐ!?J0B��_�@��_F2�ٿn
y����@!'��*4@�}�ߐ!?J0B��_�@�H_��ٿ��?1�@Y��(4@�R�cݐ!?��~��@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@�8�0y�ٿ|3p�^��@��V�,4@�Vi�;�!?K�Z���@��~��ٿʕ_���@��3�4@x��1�!?��B���@��~��ٿʕ_���@��3�4@x��1�!?��B���@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@?>dӓٿ�^y���@56�g4@� �߸�!?�I]��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@�6� '�ٿN(��@�p���4@���>��!?e]�ml��@|	�7�ٿ���@<�@DyUe��3@e�t�f�!?��z��@|	�7�ٿ���@<�@DyUe��3@e�t�f�!?��z��@|	�7�ٿ���@<�@DyUe��3@e�t�f�!?��z��@8��ӂٿ�����@�ӿ&��3@�g�φ�!?��e��/�@8��ӂٿ�����@�ӿ&��3@�g�φ�!?��e��/�@���ǆٿN!�����@����N�3@�6ׁ�!?eOm�@���ǆٿN!�����@����N�3@�6ׁ�!?eOm�@���ǆٿN!�����@����N�3@�6ׁ�!?eOm�@���ǆٿN!�����@����N�3@�6ׁ�!?eOm�@_x�Fw�ٿ˰�D~��@�j�rt 4@��dv�!?�	����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�Je�ٿ�*���@�r�A� 4@�*�5��!?����@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@�kj�F�ٿ�O��}Z�@&A\�4@5G�X�!?���LH�@Ag5�ٿ\A6���@;�1<4@[���!?���R�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@�1�3�ٿ�%�Nq=�@�+�ۏ4@��T�!?���hy�@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@ڿ�Q��ٿ�M��bG�@��4@����!?��X���@�\( ��ٿ��#A�@>��4@�O��!?�rn��@;�Ƚ��ٿrB�U��@�P�)74@�+���!?��u�@;�Ƚ��ٿrB�U��@�P�)74@�+���!?��u�@;�Ƚ��ٿrB�U��@�P�)74@�+���!?��u�@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@oX�ٿ�Q����@���Q4@�;����!?����@��jы�ٿ�����@��Tq94@u/����!?¿�s���@��jы�ٿ�����@��Tq94@u/����!?¿�s���@��jы�ٿ�����@��Tq94@u/����!?¿�s���@��jы�ٿ�����@��Tq94@u/����!?¿�s���@��jы�ٿ�����@��Tq94@u/����!?¿�s���@��jы�ٿ�����@��Tq94@u/����!?¿�s���@.�n#�ٿ�����@��\Fx�3@��W��!?�g�B��@.�n#�ٿ�����@��\Fx�3@��W��!?�g�B��@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@�� �ٿ:{j�,�@֮���4@� $Ð!?�?�)�	�@t���ٿ��i��,�@C��?�4@�L����!? D����@t���ٿ��i��,�@C��?�4@�L����!? D����@+�S��~ٿ�ԟ}�@~��&�4@���d��!?h�a/��@+�S��~ٿ�ԟ}�@~��&�4@���d��!?h�a/��@��Ue�}ٿ<{�&�@;��.4@t����!?t� �e��@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@��S�ٿ �^^�!�@)&9�n4@J)���!?�o���@�����zٿ��i%��@�L�4@f��!?��/O��@������ٿZ�J�,�@ȜY4@���!?�'��(�@������ٿZ�J�,�@ȜY4@���!?�'��(�@������ٿZ�J�,�@ȜY4@���!?�'��(�@U��O�ٿ��V�{'�@�bN��4@� Kɐ!?�IL9�6�@�<#W��ٿq\@����@HF�?Z4@DD���!?Rz/n{�@�<#W��ٿq\@����@HF�?Z4@DD���!?Rz/n{�@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@<B�|�ٿ�-�3��@僝��4@�/*J��!?R���%��@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@�F �ٿ�V�����@�AJ�k4@0o"Ð!?�n����@���܃ٿ�+����@x�u� 4@c�F~��!?H>49�@���܃ٿ�+����@x�u� 4@c�F~��!?H>49�@���܃ٿ�+����@x�u� 4@c�F~��!?H>49�@���܃ٿ�+����@x�u� 4@c�F~��!?H>49�@I���ٿG�B��@t��� 4@qm���!?�l��wb�@I���ٿG�B��@t��� 4@qm���!?�l��wb�@I���ٿG�B��@t��� 4@qm���!?�l��wb�@I���ٿG�B��@t��� 4@qm���!?�l��wb�@I���ٿG�B��@t��� 4@qm���!?�l��wb�@�����ٿSY��@�!���4@ؒ��!?I�0!��@�����ٿSY��@�!���4@ؒ��!?I�0!��@�����ٿSY��@�!���4@ؒ��!?I�0!��@�����ٿSY��@�!���4@ؒ��!?I�0!��@�����ٿSY��@�!���4@ؒ��!?I�0!��@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@L}�"��ٿ� �z���@�>ƅ4@[��W�!?�m�)�P�@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@}�ٿ�~�͖�@��Bp4@�O~���!?���Z���@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@T���ٿp�|^�/�@b��m4@�W�ե�!?��+�^��@N�U��ٿ����@�X�VT4@Q���ǐ!?���@N�U��ٿ����@�X�VT4@Q���ǐ!?���@N�U��ٿ����@�X�VT4@Q���ǐ!?���@N�U��ٿ����@�X�VT4@Q���ǐ!?���@N�U��ٿ����@�X�VT4@Q���ǐ!?���@N�U��ٿ����@�X�VT4@Q���ǐ!?���@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@��l���ٿ3��3z�@��c4@X�,�Đ!?��2-��@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@P�3�ٿȤ74���@�*e��4@b�Ύs�!?�"|S,�@?�{�y�ٿdؗȡ�@��[<�4@X]Ё��!?�����@?�{�y�ٿdؗȡ�@��[<�4@X]Ё��!?�����@?�{�y�ٿdؗȡ�@��[<�4@X]Ё��!?�����@?�{�y�ٿdؗȡ�@��[<�4@X]Ё��!?�����@�A�n�ٿH�y`P_�@A�h�4@���Ґ!?�P�7��@�A�n�ٿH�y`P_�@A�h�4@���Ґ!?�P�7��@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@,$Qtf�ٿ;/�Ф;�@q��R4@��Ү��!?pS:� H�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@$�P�ٿ�MH�7�@�OK
�4@*D��!?����C�@��8q,�ٿ0<�p���@)ȧ�P4@���ѐ!?��m��@��8q,�ٿ0<�p���@)ȧ�P4@���ѐ!?��m��@��8q,�ٿ0<�p���@)ȧ�P4@���ѐ!?��m��@��8q,�ٿ0<�p���@)ȧ�P4@���ѐ!?��m��@��� �ٿ~�8�Df�@z5��4@�<���!?b�\�~��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�*J�8�ٿ��r�c��@��'��4@�3F�x�!?j��u1��@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�|>:�ٿ`�}���@�����4@�XZDĐ!?�(�M�@�7�	�ٿ��VMM�@�ͼ�L4@t򄁻�!?RM�3�@�7�	�ٿ��VMM�@�ͼ�L4@t򄁻�!?RM�3�@�7�	�ٿ��VMM�@�ͼ�L4@t򄁻�!?RM�3�@��Dh�ٿ��G8�@7OK4@�a�{ؐ!?�ˁ���@��Dh�ٿ��G8�@7OK4@�a�{ؐ!?�ˁ���@Cs���}ٿV^4 ���@�";j�4@U�B?�!?�m�׺��@Cs���}ٿV^4 ���@�";j�4@U�B?�!?�m�׺��@*\7�Hٿ�9�wZ��@�8�4@Ҕ4ܐ!?'3p�͵�@*\7�Hٿ�9�wZ��@�8�4@Ҕ4ܐ!?'3p�͵�@��7���ٿ7���H��@(��2	4@��"��!?��A�S��@��7���ٿ7���H��@(��2	4@��"��!?��A�S��@��7���ٿ7���H��@(��2	4@��"��!?��A�S��@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@
Y�s�ٿ��SmI�@PS�� 4@��I�ϐ!?�����]�@,8/f�ٿn��f���@���i�4@���Ȑ!?k����P�@,8/f�ٿn��f���@���i�4@���Ȑ!?k����P�@,8/f�ٿn��f���@���i�4@���Ȑ!?k����P�@������ٿ��Ċg�@�xZi�4@t����!?ť6?K�@������ٿ��Ċg�@�xZi�4@t����!?ť6?K�@������ٿ��Ċg�@�xZi�4@t����!?ť6?K�@������ٿ��Ċg�@�xZi�4@t����!?ť6?K�@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@JS_тٿ�՗�x�@����64@�ŗ��!?	��+���@,��7$�ٿ��D�m�@��t��4@k% �!?�cƞ+��@,��7$�ٿ��D�m�@��t��4@k% �!?�cƞ+��@,��7$�ٿ��D�m�@��t��4@k% �!?�cƞ+��@�Ν[ȃٿ�#�����@J��nF4@��`�А!?mҼ1���@�Ν[ȃٿ�#�����@J��nF4@��`�А!?mҼ1���@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@AU-��ٿ`��ڒ�@��h�4@�q�.�!?�'��4�@7����{ٿ���e�h�@�F,�4@C�)��!?�x�(	��@w�y�}ٿ���\�@�;�O4@�p�mސ!?.�|�@w�y�}ٿ���\�@�;�O4@�p�mސ!?.�|�@w�y�}ٿ���\�@�;�O4@�p�mސ!?.�|�@w�y�}ٿ���\�@�;�O4@�p�mސ!?.�|�@w�y�}ٿ���\�@�;�O4@�p�mސ!?.�|�@؟.�(�ٿ;*z-R�@�OX
4@e���!?���}[��@؟.�(�ٿ;*z-R�@�OX
4@e���!?���}[��@؟.�(�ٿ;*z-R�@�OX
4@e���!?���}[��@g���؈ٿ�Lx���@�/=i�4@��g���!?���(�]�@��|��ٿ��'��w�@��!$4@�m3.�!?���D�[�@��|��ٿ��'��w�@��!$4@�m3.�!?���D�[�@��s^�ٿ�Ē��@��Յ4@K܉��!?��!�=�@��s^�ٿ�Ē��@��Յ4@K܉��!?��!�=�@�8魄ٿ��I� �@��sD4@�~'��!?�X�L|�@�8魄ٿ��I� �@��sD4@�~'��!?�X�L|�@��p؊ٿl1�x��@P�uB4@�ԲV|�!?W7�^�@��p؊ٿl1�x��@P�uB4@�ԲV|�!?W7�^�@J�`�a�ٿ獠4��@?�۫�4@A�yR�!?�@z�PQ�@D��Ԃٿ�˧��'�@<�v��4@�Wv6��!?�J�G�@�#a%�ٿ�_���,�@�	ˠ
4@�4hѩ�!?<!�6sX�@:l��ٿ�e&Z��@�\�4@��'��!?Ib%�@(��ٿ�-����@q���4@x�u�!?b��'���@(��ٿ�-����@q���4@x�u�!?b��'���@(��ٿ�-����@q���4@x�u�!?b��'���@(��ٿ�-����@q���4@x�u�!?b��'���@��\a+�ٿC)��:�@e�A�4@L���o�!?4g���@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@��V�ٿ5Q8��q�@��k�4@ȗY��!?�#5_��@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@�DKQ�ٿ��DXN�@�V�4@��_��!?��x�u�@��L5�ٿ�6��8�@E%e�4@�2�j�!?ф���@��1��ٿc�Q��@T5��4@6�,Ԙ�!?������@��1��ٿc�Q��@T5��4@6�,Ԙ�!?������@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@K�y�4�ٿ0������@l��u4@=�m�!?a�c��f�@��~�7�ٿ[qU\-�@|I��4@J~�!?�FL�~�@��~�7�ٿ[qU\-�@|I��4@J~�!?�FL�~�@��~�7�ٿ[qU\-�@|I��4@J~�!?�FL�~�@��~�7�ٿ[qU\-�@|I��4@J~�!?�FL�~�@��~�7�ٿ[qU\-�@|I��4@J~�!?�FL�~�@��I�8�ٿo��,�@�,��84@��}�A�!?;��ݮ@�@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@������ٿ��2ȗ�@h�'4@��JȐ!?\��"��@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@1�E:�ٿB����@�̈́o44@w��2�!?;(�G�@3�v��ٿ�F`^�b�@D��"�4@���(Ԑ!?��xg��@3�v��ٿ�F`^�b�@D��"�4@���(Ԑ!?��xg��@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@^6pXʇٿ��Usa��@4,�)�4@�}*�ǐ!?<���{�@A�}&��ٿz�iW1��@�[���4@���O��!?U&p
�@A�}&��ٿz�iW1��@�[���4@���O��!?U&p
�@A�}&��ٿz�iW1��@�[���4@���O��!?U&p
�@A�}&��ٿz�iW1��@�[���4@���O��!?U&p
�@A�}&��ٿz�iW1��@�[���4@���O��!?U&p
�@����M�ٿ#�����@�p�Y�4@�� =��!?,�t�>�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@^��لٿ�����@��[*4@=8A���!?�Ϝ�5�@]�^�y�ٿt����@6���E4@Q����!?4�\1<�@]�^�y�ٿt����@6���E4@Q����!?4�\1<�@]�^�y�ٿt����@6���E4@Q����!?4�\1<�@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@�&h�~�ٿ�����@u��5�	4@�V֐!?.�Wh���@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@F-�9�ٿp����@�\x�M4@�`B���!?���m6��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@�,T7��ٿ9Jh���@S��$�4@!��Ӑ!?��r=x��@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@v�i7�ٿ�k*b:��@�5I4@p0!�e�!?ۂ��]�@�7���ٿV�_U��@��
04@�*{Wb�!?�/�A��@�7���ٿV�_U��@��
04@�*{Wb�!?�/�A��@���j�ٿ�@w�t�@h"SN4@S.�*��!?�+��w'�@���j�ٿ�@w�t�@h"SN4@S.�*��!?�+��w'�@w�J���ٿ�ލ�^�@S b@4@+MB��!?Ԓ3�O�@w�J���ٿ�ލ�^�@S b@4@+MB��!?Ԓ3�O�@w�J���ٿ�ލ�^�@S b@4@+MB��!?Ԓ3�O�@�r0��ٿO��<���@;���4@�Ւwx�!?�V��/�@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@3���̆ٿ���7��@��K��4@3��?��!?�rfs���@���*ȅٿ�㾓�|�@i�Dw�4@�A�o{�!?,2��ߕ�@�VOZO�ٿ�C��>�@7ۙpD4@�F٤v�!?C<���@�VOZO�ٿ�C��>�@7ۙpD4@�F٤v�!?C<���@�VOZO�ٿ�C��>�@7ۙpD4@�F٤v�!?C<���@�VOZO�ٿ�C��>�@7ۙpD4@�F٤v�!?C<���@����ٿj�8��@���� 4@`��w!�!?����ʑ�@?�̯�ٿ*�mΟ��@"B�d4@�Ң�w�!?U/.�M�@H�����ٿpAf��@g,�G�4@�̽�ɐ!?��Z��Q�@0�I+�}ٿ)c�1��@0ιʹ4@�t5��!?��/;�@0�I+�}ٿ)c�1��@0ιʹ4@�t5��!?��/;�@0�I+�}ٿ)c�1��@0ιʹ4@�t5��!?��/;�@�~��(�ٿ�2$��Y�@1�a4@�L�~��!?�]�k���@�~��(�ٿ�2$��Y�@1�a4@�L�~��!?�]�k���@�~��(�ٿ�2$��Y�@1�a4@�L�~��!?�]�k���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@�M�P�ٿblҤMI�@1� �4@Ae��!?"IF���@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@k{q��ٿc� L_�@�����4@�R^܏�!?'����X�@�ov2K�ٿ��nخ�@4ʁ,�4@2���m�!?����t��@�ov2K�ٿ��nخ�@4ʁ,�4@2���m�!?����t��@�ov2K�ٿ��nخ�@4ʁ,�4@2���m�!?����t��@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@�1��
�ٿ��v5��@q;c�4@�#��!?�W��`}�@w{���ٿ��-�@�q��F4@�g@���!?��SF	�@w{���ٿ��-�@�q��F4@�g@���!?��SF	�@,�)Մٿ��=n���@�~ˉ4@z��ɐ!?�C����@,�)Մٿ��=n���@�~ˉ4@z��ɐ!?�C����@,�)Մٿ��=n���@�~ˉ4@z��ɐ!?�C����@��xf��ٿ��Q���@'��v4@@S����!?B�����@��xf��ٿ��Q���@'��v4@@S����!?B�����@��xf��ٿ��Q���@'��v4@@S����!?B�����@��xf��ٿ��Q���@'��v4@@S����!?B�����@��xf��ٿ��Q���@'��v4@@S����!?B�����@W�ʇٿh�N-#�@q8�$�4@٣�^��!?N��/���@W�ʇٿh�N-#�@q8�$�4@٣�^��!?N��/���@��L��ٿ�w�b:�@�<�^�4@'��)ِ!?&���:G�@��L��ٿ�w�b:�@�<�^�4@'��)ِ!?&���:G�@� 	F��ٿ�O��@��3� 4@�K�!��!?��N���@�ݑC�ٿ������@[~�[�4@���!?���\���@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@��i�c�ٿS��t�S�@y��C�4@��j�Ԑ!?���#w|�@�Q}��ٿ'��=>��@��Eb�4@`�X���!?�o�b�@�Q}��ٿ'��=>��@��Eb�4@`�X���!?�o�b�@�Q}��ٿ'��=>��@��Eb�4@`�X���!?�o�b�@�6^�ٿ*/.e���@8�q�4@	�_�!?�`;v@�@�6^�ٿ*/.e���@8�q�4@	�_�!?�`;v@�@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@�*l�l�ٿi�X���@��)�4@�7lÐ!?�9����@E�Z�ٿ��ؗ��@gÍ�4@�yԐ!?�C7���@E�Z�ٿ��ؗ��@gÍ�4@�yԐ!?�C7���@E�Z�ٿ��ؗ��@gÍ�4@�yԐ!?�C7���@E�Z�ٿ��ؗ��@gÍ�4@�yԐ!?�C7���@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@��C~ٿ�n����@~<��F4@�Z��ː!?Il�p��@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@�l��ٿK�� ���@�_��x4@���ΐ!?������@��[虁ٿ�l��3��@6�u4@R	�}��!?z8;u���@��[虁ٿ�l��3��@6�u4@R	�}��!?z8;u���@��[虁ٿ�l��3��@6�u4@R	�}��!?z8;u���@�i�x�ٿ�'2�h�@$?�m4@N��죐!?��'��@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@���=ńٿ�!�s.d�@aR��4@%���!?�}\rN�@��^=��ٿd�%@�@n�4�J4@�l��Ӑ!?#�#w��@��^=��ٿd�%@�@n�4�J4@�l��Ӑ!?#�#w��@��^=��ٿd�%@�@n�4�J4@�l��Ӑ!?#�#w��@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@
����ٿ���o��@L�h�k4@��Z�!?��6-���@FC}u�ٿѝC{D�@f���4@j��2��!?8���K��@ގ���ٿ�v��@NZĹ4@�4�U�!?�2K��@_gY�ٿ�����@+TZ4@a�*ϵ�!?q$��R�@C��Se�ٿ�X4(%��@���s�4@��ㄒ�!?�jG�g��@vr�Ӌٿl�R3���@�L��4@�:i%��!?.n�qc��@��}�1�ٿ��>��?�@�`��]4@d��!?	\�\�@��+�ٿ� ��VZ�@[(_4@`��Y�!?��wҵ�@��+�ٿ� ��VZ�@[(_4@`��Y�!?��wҵ�@��+�ٿ� ��VZ�@[(_4@`��Y�!?��wҵ�@�/�O�ٿ�@��7��@��:<4@�h��А!?�,}�n�@Pƫ���ٿ�gz����@��mÝ4@D�;n�!?�#�z��@���.�ٿ'���@����4@	Y� m�!?���`��@���.�ٿ'���@����4@	Y� m�!?���`��@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@��`g�ٿ՟�n׊�@�EYiw4@�\��ː!?������@u.m�}ٿ�d��=[�@m�c�4@�N��!?S#,��@u.m�}ٿ�d��=[�@m�c�4@�N��!?S#,��@u.m�}ٿ�d��=[�@m�c�4@�N��!?S#,��@�*JP�}ٿ�i�����@0 �4@ǧ結!?o�����@�*JP�}ٿ�i�����@0 �4@ǧ結!?o�����@��M�ٿ�9�I��@�5��4@o�9G��!?��*T���@��M�ٿ�9�I��@�5��4@o�9G��!?��*T���@<J�\?�ٿq�XY�T�@֋���4@B���Ő!?�ֳ��{�@<J�\?�ٿq�XY�T�@֋���4@B���Ő!?�ֳ��{�@<J�\?�ٿq�XY�T�@֋���4@B���Ő!?�ֳ��{�@<J�\?�ٿq�XY�T�@֋���4@B���Ő!?�ֳ��{�@<J�\?�ٿq�XY�T�@֋���4@B���Ő!?�ֳ��{�@R�B��ٿy���(��@b�5��4@&q���!?r�H/q�@R�B��ٿy���(��@b�5��4@&q���!?r�H/q�@"B�N2�ٿ�4����@g�k34@J��^�!?Zn���o�@"B�N2�ٿ�4����@g�k34@J��^�!?Zn���o�@"B�N2�ٿ�4����@g�k34@J��^�!?Zn���o�@N�ͣ�ٿ��%����@�[E"�4@�� ;�!?��K>�@N�ͣ�ٿ��%����@�[E"�4@�� ;�!?��K>�@N�ͣ�ٿ��%����@�[E"�4@�� ;�!?��K>�@޶hq~ٿ�����@���4@onZ�J�!?����B�@��[z�}ٿX��$5k�@��lv,4@[�v>�!?')X��O�@��[z�}ٿX��$5k�@��lv,4@[�v>�!?')X��O�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@�p��Q�ٿwF����@B
���4@�E9��!?<��城�@yӠ_�ٿ���!��@7"�d�4@|;|�!?�M{ã�@yӠ_�ٿ���!��@7"�d�4@|;|�!?�M{ã�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@d-�1�ٿ?5,3M�@��Ė�4@M1���!?0�evl�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�q�dA�ٿz@1'���@?�#�4@���c��!?�'�6�@�*���ٿ)N�}��@.��4@�ڴ۞�!?����
�@�*���ٿ)N�}��@.��4@�ڴ۞�!?����
�@�*���ٿ)N�}��@.��4@�ڴ۞�!?����
�@�*���ٿ)N�}��@.��4@�ڴ۞�!?����
�@�*���ٿ)N�}��@.��4@�ڴ۞�!?����
�@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@mn$�ٿ[���@�R��4@9�Hkː!?��"����@�����ٿG�����@p�Y�4@���ٽ�!?P�a�q�@�����ٿG�����@p�Y�4@���ٽ�!?P�a�q�@�����ٿG�����@p�Y�4@���ٽ�!?P�a�q�@�����ٿG�����@p�Y�4@���ٽ�!?P�a�q�@����ٿ�h�>t�@QYkf4@D{�IĐ!?/��.(�@����ٿ�h�>t�@QYkf4@D{�IĐ!?/��.(�@����ٿ�h�>t�@QYkf4@D{�IĐ!?/��.(�@���Xٿ���?���@�J�^�4@S[���!?��:JG��@���Xٿ���?���@�J�^�4@S[���!?��:JG��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@�)�{��ٿ�l���@K�8�X4@�γ���!?g򐺙��@Nr_���ٿ�Cv��l�@�PQ4@Z��!?b��1��@Nr_���ٿ�Cv��l�@�PQ4@Z��!?b��1��@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@"���ٿ��) 3�@.��k4@��s�q�!?hR���@ BI�[�ٿG]d��@�^ �4@1�Aא!?RD�¿�@ BI�[�ٿG]d��@�^ �4@1�Aא!?RD�¿�@/�{�G�ٿ�4��B�@���@�4@�*���!?�oWC+��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�����ٿ�A(3���@`�^�j4@�Ͽ���!?�� �a��@�=LV�ٿ��I�@D�q�4@v����!?~	B����@�ϺӮ�ٿ�Y.���@Ǩ���4@G\��Đ!?n���wT�@�ϺӮ�ٿ�Y.���@Ǩ���4@G\��Đ!?n���wT�@F��m�ٿ�܊���@k�X 4@����!?��+G�@F��m�ٿ�܊���@k�X 4@����!?��+G�@F��m�ٿ�܊���@k�X 4@����!?��+G�@F��m�ٿ�܊���@k�X 4@����!?��+G�@F��m�ٿ�܊���@k�X 4@����!?��+G�@F��m�ٿ�܊���@k�X 4@����!?��+G�@)�("�ٿ�kȕ`��@�u��4@{�����!?O�hh���@)�("�ٿ�kȕ`��@�u��4@{�����!?O�hh���@)�("�ٿ�kȕ`��@�u��4@{�����!?O�hh���@�U���ٿ(l"fv�@�|MC4@�/	��!?Ͱ�՚��@�U���ٿ(l"fv�@�|MC4@�/	��!?Ͱ�՚��@�U���ٿ(l"fv�@�|MC4@�/	��!?Ͱ�՚��@�U���ٿ(l"fv�@�|MC4@�/	��!?Ͱ�՚��@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@I�4��ٿs�g��D�@6��~�4@ ݬG�!?vjOWSb�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@~p +�ٿMj$`��@�j��4@�&��2�!?$���(�@W����ٿ��J���@���ĸ4@�R��!?��@�@�@W����ٿ��J���@���ĸ4@�R��!?��@�@�@W����ٿ��J���@���ĸ4@�R��!?��@�@�@Q$���ٿ�j�x�[�@x�T�4@������!?��as��@Q$���ٿ�j�x�[�@x�T�4@������!?��as��@Q$���ٿ�j�x�[�@x�T�4@������!?��as��@Q$���ٿ�j�x�[�@x�T�4@������!?��as��@E�~ٿ�V.K��@�:O�	4@�h���!?"Fڥ���@E�~ٿ�V.K��@�:O�	4@�h���!?"Fڥ���@E�~ٿ�V.K��@�:O�	4@�h���!?"Fڥ���@E�~ٿ�V.K��@�:O�	4@�h���!?"Fڥ���@���_�ٿ ����@T�Rce4@���䞐!??0BQl��@Oy.r|�ٿ_��3��@��:C4@}4+���!?��m�1��@Ps+Pc�ٿ7L^�3�@<�n�4@y�mk�!?b/�U�@��A�7�ٿ���i�]�@�$w�64@�ag�ǐ!?�\ګEa�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@�%5�ٿ�6��IN�@g�{=4@KP��!?kCp?�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@.�e�%�ٿ�ɸ���@J�~�y4@<�q�n�!?�Dp�,A�@���ٿ�����W�@��44@�A}��!?�c���@���ٿ�����W�@��44@�A}��!?�c���@ 2̋��ٿ�N�EX�@0��6�4@D�u��!?��k#��@ 2̋��ٿ�N�EX�@0��6�4@D�u��!?��k#��@ 2̋��ٿ�N�EX�@0��6�4@D�u��!?��k#��@s{&�b�ٿA��%��@}�l:4@��{E�!?�?���@s{&�b�ٿA��%��@}�l:4@��{E�!?�?���@s{&�b�ٿA��%��@}�l:4@��{E�!?�?���@s{&�b�ٿA��%��@}�l:4@��{E�!?�?���@s{&�b�ٿA��%��@}�l:4@��{E�!?�?���@�)Y<�ٿY�民��@=�X��4@s��C�!?�{��=�@�)Y<�ٿY�民��@=�X��4@s��C�!?�{��=�@N֍Íٿ��iv�@*�C�4@��t"�!?Û&4��@N֍Íٿ��iv�@*�C�4@��t"�!?Û&4��@N֍Íٿ��iv�@*�C�4@��t"�!?Û&4��@��ٌ�ٿ�Gc�a��@z��!&4@y�+��!?�8�P��@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@�����ٿ%x��l�@�{��	4@5V�ݠ�!?p�w'�@e����ٿ_��G�@z~�V�4@���!?۹��1�@e����ٿ_��G�@z~�V�4@���!?۹��1�@e����ٿ_��G�@z~�V�4@���!?۹��1�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@h;�Z^~ٿ	�B�@
���4@�LU/��!?�9��&�@O�IͿzٿW� �Q��@H�'³4@�� ��!?��>��@O�IͿzٿW� �Q��@H�'³4@�� ��!?��>��@O�IͿzٿW� �Q��@H�'³4@�� ��!?��>��@O�IͿzٿW� �Q��@H�'³4@�� ��!?��>��@O�IͿzٿW� �Q��@H�'³4@�� ��!?��>��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@.��=�ٿ��q5�@��;j4@�>Zս�!?\��r'��@��G���ٿe,N$�@IC�?�4@��y�א!?%xΡ��@��G���ٿe,N$�@IC�?�4@��y�א!?%xΡ��@��G���ٿe,N$�@IC�?�4@��y�א!?%xΡ��@��G���ٿe,N$�@IC�?�4@��y�א!?%xΡ��@<����ٿ��&�O2�@U(b�l4@��g��!?c�� r�@<����ٿ��&�O2�@U(b�l4@��g��!?c�� r�@<����ٿ��&�O2�@U(b�l4@��g��!?c�� r�@��� �ٿh�H P��@eƒ�h4@���0�!?7_�E6e�@��� �ٿh�H P��@eƒ�h4@���0�!?7_�E6e�@��� �ٿh�H P��@eƒ�h4@���0�!?7_�E6e�@�z}��ٿ⶝����@/W�Q� 4@�<n��!?���Y��@WM���ٿJ�]}�@���3@���1�!?�bg�7��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�Mj��ٿ�#��n�@�����4@���!?#+�N��@�6���ٿ�7�q`�@����I4@�+���!?#3�����@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@N��~ٿ.hr����@�S0�4@���!?�Ю^�E�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@��	1Zٿ��x�v�@�C�4@�|oFǐ!?��Lxל�@�,ҁٿ��pV��@�����4@4�p���!?vY����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@٣�l�ٿ�`���%�@��wcZ4@yw���!?����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@ᓏrʄٿ�[�s�@��s�4@����!?R	�����@C8���~ٿ�Z�q&w�@N�<�4@"����!?�+� l�@C8���~ٿ�Z�q&w�@N�<�4@"����!?�+� l�@C8���~ٿ�Z�q&w�@N�<�4@"����!?�+� l�@C8���~ٿ�Z�q&w�@N�<�4@"����!?�+� l�@C8���~ٿ�Z�q&w�@N�<�4@"����!?�+� l�@0k'��ٿ�����@��}��4@�� �ې!?�A����@0k'��ٿ�����@��}��4@�� �ې!?�A����@0k'��ٿ�����@��}��4@�� �ې!?�A����@0k'��ٿ�����@��}��4@�� �ې!?�A����@0k'��ٿ�����@��}��4@�� �ې!?�A����@0k'��ٿ�����@��}��4@�� �ې!?�A����@����ٿ<����@9�%��4@AwR���!?m=9F��@����ٿ<����@9�%��4@AwR���!?m=9F��@>x�교ٿY���i7�@�N�!�4@��h��!?���d��@>x�교ٿY���i7�@�N�!�4@��h��!?���d��@�oOD��ٿ.�����@�,��`4@���!?
a��@]�H���ٿ��`�oc�@��ɔ�4@�j��!?��
���@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@J�%E�ٿt]IK���@����4@��1�!?y��י��@"m�T�ٿ��t+�w�@Q$�	4@��J��!?ս�r���@"m�T�ٿ��t+�w�@Q$�	4@��J��!?ս�r���@"m�T�ٿ��t+�w�@Q$�	4@��J��!?ս�r���@�m��i�ٿ�n|�d�@#"�e�4@��,̈�!?�F����@�m��i�ٿ�n|�d�@#"�e�4@��,̈�!?�F����@���ٿ����\�@=`���3@�(-)��!?�ު��`�@���ٿ����\�@=`���3@�(-)��!?�ު��`�@���ٿ����\�@=`���3@�(-)��!?�ު��`�@�ݴn�ٿ*��Y�S�@J��3@8��ڑ�!?���,���@�ݴn�ٿ*��Y�S�@J��3@8��ڑ�!?���,���@�ݴn�ٿ*��Y�S�@J��3@8��ڑ�!?���,���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@T��K�ٿ�S#,bX�@ ����4@å0ې!?Jh���@e�1x�ٿ�J�<Ub�@QK�4@R���!?���h��@e�1x�ٿ�J�<Ub�@QK�4@R���!?���h��@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@W
v�ʂٿ��+�@��B�4@X%v��!?��a�q�@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@iL`��ٿ��qD^��@a;w4@5�$���!?�L�P��@��s&�zٿ���)��@.#�] 4@�(B���!?ٞL-z�@�yV�,yٿn������@Կa~�4@r�p{Ð!?���"�A�@�yV�,yٿn������@Կa~�4@r�p{Ð!?���"�A�@�yV�,yٿn������@Կa~�4@r�p{Ð!?���"�A�@�yV�,yٿn������@Կa~�4@r�p{Ð!?���"�A�@yp�cAvٿq�鄤��@iAS�m4@Nh;��!?�\U{�@yp�cAvٿq�鄤��@iAS�m4@Nh;��!?�\U{�@�VH=wٿ{f�����@�;9��4@��Jא!?��!×u�@�VH=wٿ{f�����@�;9��4@��Jא!?��!×u�@�VH=wٿ{f�����@�;9��4@��Jא!?��!×u�@��28~ٿ��r-߉�@S��4@����!?Y��U�@��28~ٿ��r-߉�@S��4@����!?Y��U�@��28~ٿ��r-߉�@S��4@����!?Y��U�@�xҺq�ٿ����@��"84@��Ù�!?Ĵq�9��@�xҺq�ٿ����@��"84@��Ù�!?Ĵq�9��@0�#���ٿ�R�7��@6j�o4@�l�5��!?dp��|n�@@�"��ٿ�g�b�#�@b���4@2���ǐ!?�}����@@�"��ٿ�g�b�#�@b���4@2���ǐ!?�}����@@�"��ٿ�g�b�#�@b���4@2���ǐ!?�}����@@�"��ٿ�g�b�#�@b���4@2���ǐ!?�}����@�ǎ/)�ٿ�l��M�@B��=�4@�e�w��!?%����@S��݈ٿ�2㒘��@����4@l�8r�!?�AVɦ`�@S��݈ٿ�2㒘��@����4@l�8r�!?�AVɦ`�@S��݈ٿ�2㒘��@����4@l�8r�!?�AVɦ`�@S��݈ٿ�2㒘��@����4@l�8r�!?�AVɦ`�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@�qJRٿ���Tr�@#u�S4@�7��!?� ��3�@ǐxˇٿ�u�+Tv�@�'�7"4@����]�!?��Y����@��d��zٿ�e�-<��@��aX\4@	����!?��K�U��@%V���ٿB?^�T�@���� 4@�*��{�!?�s
���@�^�Z��ٿ�qS�Z�@��c>�4@��*���!?܉��ka�@����ٿ�é\W��@_]�~� 4@bd+xؐ!?�=�L;�@����ٿ�é\W��@_]�~� 4@bd+xؐ!?�=�L;�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�n�N�ٿ�h2����@3�!�4@���I��!?���I�@�4R��ٿ#��^��@c���4@�$�!?�k�[��@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@��C�ٿI�ȼ��@�S��y4@9V�B��!?xЃ��$�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@�-��Όٿݶr����@�R=�W4@��-��!?��?W�9�@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@���Q�ٿ�Qd�p�@Ȓ�4@�)v��!?��Q#���@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@r�u��}ٿ	6M���@t�4:4@%��@��!?9�!��!�@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@�o���ٿɡ�t��@��G���3@��Ɍ�!?��z2��@"��ɀٿ��b�8��@��(�d4@������!?�#��m�@"��ɀٿ��b�8��@��(�d4@������!?�#��m�@"��ɀٿ��b�8��@��(�d4@������!?�#��m�@"��ɀٿ��b�8��@��(�d4@������!?�#��m�@8p9n�ٿ㠀���@
�o��4@��Lk��!?
��v�@+���׋ٿ�oE�`��@�r4�.4@�~�ɐ!?Y<�)���@+���׋ٿ�oE�`��@�r4�.4@�~�ɐ!?Y<�)���@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@��N�ٿĘ���r�@�n1��4@��_��!?�@�@O�=>֊ٿ�:X�Ô�@�	C��4@=����!?aW _h�@O�=>֊ٿ�:X�Ô�@�	C��4@=����!?aW _h�@O�=>֊ٿ�:X�Ô�@�	C��4@=����!?aW _h�@O�=>֊ٿ�:X�Ô�@�	C��4@=����!?aW _h�@O�=>֊ٿ�:X�Ô�@�	C��4@=����!?aW _h�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@��[x߄ٿ۱�����@�>[O�4@�l�;ؐ!?�⎶ո�@I0�
�ٿEZ�T|��@s��4@�5�oÐ!?�z4���@Ӯ� 1�ٿ_�j��@��v�4@g��!?�۸>b��@~�5��ٿ& �6���@����4@8��!?$͆ ���@~�5��ٿ& �6���@����4@8��!?$͆ ���@�3�/=�ٿ�TN���@�N��� 4@�ȴm��!?6kb9��@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@��SI�ٿ��� C&�@`C��}4@�.B9y�!?
��Fa5�@����چٿ���$��@�<�@4@����!?�E���@�؉c�ٿ�u�����@yj�44@�����!?=#9�D�@�؉c�ٿ�u�����@yj�44@�����!?=#9�D�@�o�;�ٿ��� B��@��44@�-��ې!?<�M	��@W=A��ٿ0Ӑ1[��@�X.D4@l��ߐ!?�F�_�@W=A��ٿ0Ӑ1[��@�X.D4@l��ߐ!?�F�_�@W=A��ٿ0Ӑ1[��@�X.D4@l��ߐ!?�F�_�@K��4��ٿ6���@���0t4@`K�?��!?؅(*�h�@K��4��ٿ6���@���0t4@`K�?��!?؅(*�h�@-�?��ٿ�?�j+�@:M��>4@�?��А!?�h�X�@-�?��ٿ�?�j+�@:M��>4@�?��А!?�h�X�@�����ٿ�Y����@�{��4@�j�y��!?i�{K��@�����ٿ�Y����@�{��4@�j�y��!?i�{K��@"M_j�ٿ���-�6�@�YG��4@Tt��ސ!?�S]����@"M_j�ٿ���-�6�@�YG��4@Tt��ސ!?�S]����@�m��!�ٿ�^�$'V�@�1�R�4@&ژ�͐!?��Զ?L�@�m��!�ٿ�^�$'V�@�1�R�4@&ژ�͐!?��Զ?L�@�m��!�ٿ�^�$'V�@�1�R�4@&ژ�͐!?��Զ?L�@�m��!�ٿ�^�$'V�@�1�R�4@&ژ�͐!?��Զ?L�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�9�l4�ٿ���\C�@���v4@呢ڐ!?;8��l[�@�lF��ٿ<�b��@��ۅ4@�ӻ��!?#}nT;n�@�lF��ٿ<�b��@��ۅ4@�ӻ��!?#}nT;n�@�lF��ٿ<�b��@��ۅ4@�ӻ��!?#}nT;n�@|��`�ٿ'��!���@D��4@�V�	�!?�rk�S�@|��`�ٿ'��!���@D��4@�V�	�!?�rk�S�@|��`�ٿ'��!���@D��4@�V�	�!?�rk�S�@lֱ�r�ٿ��ھn�@�ʭS�4@�l#Gِ!?dQ&�w��@lֱ�r�ٿ��ھn�@�ʭS�4@�l#Gِ!?dQ&�w��@lֱ�r�ٿ��ھn�@�ʭS�4@�l#Gِ!?dQ&�w��@lֱ�r�ٿ��ھn�@�ʭS�4@�l#Gِ!?dQ&�w��@!��\��ٿ��f����@	݄4�4@'5K��!?n���V�@!��\��ٿ��f����@	݄4�4@'5K��!?n���V�@!��\��ٿ��f����@	݄4�4@'5K��!?n���V�@!��\��ٿ��f����@	݄4�4@'5K��!?n���V�@��F��ٿJ�{T��@��lt4@U��q�!?l7�sY�@y PP�ٿ��y��@z��f4@f�܆m�!?������@y PP�ٿ��y��@z��f4@f�܆m�!?������@f�9���ٿ�=���@Q0���4@�t[ː!?^�_����@ׅ�(̑ٿ��Z��@ՠX{�4@x	�m�!?��z�
�@rV�u��ٿ������@S�yxw4@����!?��:�@rV�u��ٿ������@S�yxw4@����!?��:�@rV�u��ٿ������@S�yxw4@����!?��:�@rV�u��ٿ������@S�yxw4@����!?��:�@rV�u��ٿ������@S�yxw4@����!?��:�@����	�ٿ'�p7I'�@�[��_4@�B����!?5x`���@����ٿ�QVe�B�@�c;�/4@��wx�!?�S���4�@|YY�b�ٿa�	�p�@�ҮD�4@�%�z�!?�ݧ"�j�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@T�8X��ٿ���+Hx�@�->C}4@�ñ���!?�	-��.�@�pxQ��ٿq
�6��@�Q}ڲ4@۷j��!?�p�U:�@�pxQ��ٿq
�6��@�Q}ڲ4@۷j��!?�p�U:�@�pxQ��ٿq
�6��@�Q}ڲ4@۷j��!?�p�U:�@�pxQ��ٿq
�6��@�Q}ڲ4@۷j��!?�p�U:�@�pxQ��ٿq
�6��@�Q}ڲ4@۷j��!?�p�U:�@38N�<�ٿ}��ӷ��@�@�o4@��!?tp�i=�@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@Tf{�Đٿ.�+[��@T�4@��	�!?F�i�\��@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@���ŋٿ�>I����@�����	4@��`���!?�����/�@sH?i�ٿ#=��
��@���
4@�G��!?N��O���@���ٿ������@XՏ7F
4@�"L�Ȑ!?�zZ1��@���ٿ������@XՏ7F
4@�"L�Ȑ!?�zZ1��@���ٿ������@XՏ7F
4@�"L�Ȑ!?�zZ1��@�3n�΃ٿ%�"��@22]/�4@�+C��!?�8�C��@�3n�΃ٿ%�"��@22]/�4@�+C��!?�8�C��@�3n�΃ٿ%�"��@22]/�4@�+C��!?�8�C��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@ʈ�2��ٿ����@.X.4@��k!?։�@��@���"��ٿEp�nz�@�?���4@�e�!?�3v5%�@���"��ٿEp�nz�@�?���4@�e�!?�3v5%�@���"��ٿEp�nz�@�?���4@�e�!?�3v5%�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@T��OJ�ٿ,b�[�@G�8�#4@Ҽ;���!?�8�(�0�@�_�_�ٿ�K�!|�@���ʷ4@�mW��!?��#.���@�_�_�ٿ�K�!|�@���ʷ4@�mW��!?��#.���@�_�_�ٿ�K�!|�@���ʷ4@�mW��!?��#.���@�_�_�ٿ�K�!|�@���ʷ4@�mW��!?��#.���@�_�_�ٿ�K�!|�@���ʷ4@�mW��!?��#.���@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@Hk��Q�ٿ�aj�@r�!g_4@-P���!?y B�y�@oN��	�ٿs��[���@6���4@�;�}�!?>��L&�@oN��	�ٿs��[���@6���4@�;�}�!?>��L&�@oN��	�ٿs��[���@6���4@�;�}�!?>��L&�@oN��	�ٿs��[���@6���4@�;�}�!?>��L&�@oN��	�ٿs��[���@6���4@�;�}�!?>��L&�@�{���ٿ���|��@�_x�4@R9�3��!?�}��.�@�{���ٿ���|��@�_x�4@R9�3��!?�}��.�@~���=�ٿ5u�D_��@(D��4@tF����!?���ŷ��@~���=�ٿ5u�D_��@(D��4@tF����!?���ŷ��@~���=�ٿ5u�D_��@(D��4@tF����!?���ŷ��@@ق�4�ٿ�:I�`��@���8M�3@b~�6��!?ӈ&�@T'���yٿ`��I���@&ܰ#��3@����!?��z�E��@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@�X�yٿ*����@�p	5W 4@�w���!?6��R|�@���|ٿME�j֬�@W��4@�[�&��!?!�Ft��@���|ٿME�j֬�@W��4@�[�&��!?!�Ft��@��H��ٿ�v���@g�i`h4@�0G�ϐ!?�� Fv��@��b'�}ٿ2����.�@�(��4@����!?��mh�@C��;~�ٿ=���(�@�Q]Ui4@����!?!C5�'�@C��;~�ٿ=���(�@�Q]Ui4@����!?!C5�'�@C��;~�ٿ=���(�@�Q]Ui4@����!?!C5�'�@C��;~�ٿ=���(�@�Q]Ui4@����!?!C5�'�@C��;~�ٿ=���(�@�Q]Ui4@����!?!C5�'�@�)��ȂٿX|��@�_3�4@b&���!?�t�ov��@�)��ȂٿX|��@�_3�4@b&���!?�t�ov��@�)��ȂٿX|��@�_3�4@b&���!?�t�ov��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@-��Y��ٿ#�7���@��,j�4@��񷾐!?�GTv��@OPt���ٿ�+��@b+�W:4@E���!?���Q�G�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@U�.���ٿ�Ű�1��@��54@ۀ����!?s�f��\�@(���ٿ�6	����@�%ȉ4@��Ԑ!?��3���@(���ٿ�6	����@�%ȉ4@��Ԑ!?��3���@(���ٿ�6	����@�%ȉ4@��Ԑ!?��3���@� �n��ٿ�	۰���@��j�� 4@��˫�!?�����@� �n��ٿ�	۰���@��j�� 4@��˫�!?�����@� �n��ٿ�	۰���@��j�� 4@��˫�!?�����@� �n��ٿ�	۰���@��j�� 4@��˫�!?�����@� �n��ٿ�	۰���@��j�� 4@��˫�!?�����@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@�&u2�ٿR��>�@3��	\4@o��r��!?/�!c���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@WL�@��ٿ���a��@b��4@#Z ˘�!?��jo���@�3f��ٿ�Q�
��@��8�<4@L��!?˻����@�3f��ٿ�Q�
��@��8�<4@L��!?˻����@�3f��ٿ�Q�
��@��8�<4@L��!?˻����@�3f��ٿ�Q�
��@��8�<4@L��!?˻����@�3f��ٿ�Q�
��@��8�<4@L��!?˻����@��=��ٿ��>P���@�A?�� 4@&��Ɣ�!?B��B���@��=��ٿ��>P���@�A?�� 4@&��Ɣ�!?B��B���@��=��ٿ��>P���@�A?�� 4@&��Ɣ�!?B��B���@��=��ٿ��>P���@�A?�� 4@&��Ɣ�!?B��B���@��=��ٿ��>P���@�A?�� 4@&��Ɣ�!?B��B���@,L���ٿ��o	Bq�@��Oz84@a�r�!?����@,L���ٿ��o	Bq�@��Oz84@a�r�!?����@���&��ٿ�2�,8��@r��_&4@�j��ϐ!?��8��i�@���&��ٿ�2�,8��@r��_&4@�j��ϐ!?��8��i�@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@ �$�<�ٿ��� ��@��<4@�zݐ!?�n��0��@�� C�ٿ�+sk��@ϐMr�4@б�t��!?#y@ʼ0�@�� C�ٿ�+sk��@ϐMr�4@б�t��!?#y@ʼ0�@�� C�ٿ�+sk��@ϐMr�4@б�t��!?#y@ʼ0�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@�te�A�ٿ�-�(�@���%�4@O#ʔݐ!?�Ls�j�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@/N[=�ٿ{�b,�@F�<��4@m����!?�"[�Q%�@\�t���ٿ���:��@y��g� 4@_)l��!?�q�3�@.[��ٿ 4��ƻ�@��UU�4@��-�\�!?��䙭�@.[��ٿ 4��ƻ�@��UU�4@��-�\�!?��䙭�@.[��ٿ 4��ƻ�@��UU�4@��-�\�!?��䙭�@�?��ٿ�MkҖ�@��'l4@���IC�!?d~:O���@�?��ٿ�MkҖ�@��'l4@���IC�!?d~:O���@�?��ٿ�MkҖ�@��'l4@���IC�!?d~:O���@�O뀭�ٿ�XIvx��@'g$4�4@>��v�!?��̱���@ɋ�	��ٿ�rg���@���4 4@hO�A�!?}�OBw��@<F?Ήٿ0km|��@�G�{4@��E�!?=������@<F?Ήٿ0km|��@�G�{4@��E�!?=������@3�AV��ٿE��8���@�f�y+4@���'�!?�v�D�X�@3�AV��ٿE��8���@�f�y+4@���'�!?�v�D�X�@<�3==�ٿ��qfJ;�@�7Ɂ*	4@@X�ͤ�!?��Fz��@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@Q_�;��ٿ�ɵ����@V&-/4@\É�!?q����@}�4�p�ٿ��Vw��@��	�4@��R�ߐ!?�����@}�4�p�ٿ��Vw��@��	�4@��R�ߐ!?�����@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@,j� ��ٿ9��o�@ܣZy�4@�a
B��!?� #磾�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@�
5�ٿcC����@����4@���Q��!?y�G�@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@K�`�ٿ�%?oU�@m��(�4@\{���!?��KV��@c7��߄ٿ'��M��@�5��.4@��V6��!?��G��H�@c7��߄ٿ'��M��@�5��.4@��V6��!?��G��H�@JO6�7�ٿiF��N�@�_�:�4@Q�z^�!?�1�~Ed�@JO6�7�ٿiF��N�@�_�:�4@Q�z^�!?�1�~Ed�@JO6�7�ٿiF��N�@�_�:�4@Q�z^�!?�1�~Ed�@JO6�7�ٿiF��N�@�_�:�4@Q�z^�!?�1�~Ed�@JO6�7�ٿiF��N�@�_�:�4@Q�z^�!?�1�~Ed�@���P�ٿ�FhT��@O��Mj4@T��F�!?������@���P�ٿ�FhT��@O��Mj4@T��F�!?������@���P�ٿ�FhT��@O��Mj4@T��F�!?������@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�5��ٿΆM���@���N)4@sD�俐!?C�7�z�@�w�@C�ٿ��:�@��4@��[N�!?\�f��@�w�@C�ٿ��:�@��4@��[N�!?\�f��@�w�@C�ٿ��:�@��4@��[N�!?\�f��@RUi��ٿ^}����@S�CD4@jĿYB�!?���u'�@RUi��ٿ^}����@S�CD4@jĿYB�!?���u'�@RUi��ٿ^}����@S�CD4@jĿYB�!?���u'�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@�޹ǂٿ@C�^���@����4@�&�͐!?�����h�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@ǕH)��ٿr�nL���@<��p�4@�����!?Em;)�t�@��6�z�ٿ�S�p�Y�@��g�j4@����!?�Nn��@��6�z�ٿ�S�p�Y�@��g�j4@����!?�Nn��@��6�z�ٿ�S�p�Y�@��g�j4@����!?�Nn��@��6�z�ٿ�S�p�Y�@��g�j4@����!?�Nn��@uV(<قٿM��Q�)�@-����4@�����!?o��[$��@�jn|(}ٿr"'�KL�@1%�i�4@�hhܴ�!?�%�>�@Qu�zr�ٿ�����@�j�ş4@�~�z7�!?�,D!��@Qu�zr�ٿ�����@�j�ş4@�~�z7�!?�,D!��@Qu�zr�ٿ�����@�j�ş4@�~�z7�!?�,D!��@CM{�y�ٿh6k���@�|�I34@)��a �!?�zz5H��@CM{�y�ٿh6k���@�|�I34@)��a �!?�zz5H��@CM{�y�ٿh6k���@�|�I34@)��a �!?�zz5H��@��"L��ٿ ���ԋ�@g3z�G4@���!?�	�Fk�@��E�ٿ��2<+�@��)	4@���!?���:���@��E�ٿ��2<+�@��)	4@���!?���:���@��E�ٿ��2<+�@��)	4@���!?���:���@��E�ٿ��2<+�@��)	4@���!?���:���@��E�ٿ��2<+�@��)	4@���!?���:���@�zec�ٿ8t
3:_�@X�p6�4@e��!�!?X�z	6��@�zec�ٿ8t
3:_�@X�p6�4@e��!�!?X�z	6��@�_�J�ٿ�%���\�@4m,}O4@�"$V?�!?����A�@�_�J�ٿ�%���\�@4m,}O4@�"$V?�!?����A�@�u��`{ٿ����z�@<���"4@~����!? }�Ԟ�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@"�h�{ٿ�h�F�@���a-4@ľ: ��!?���(�K�@JL��}ٿc'`�4��@N�V4@Bs��!?�FY�]��@JL��}ٿc'`�4��@N�V4@Bs��!?�FY�]��@JL��}ٿc'`�4��@N�V4@Bs��!?�FY�]��@JL��}ٿc'`�4��@N�V4@Bs��!?�FY�]��@JL��}ٿc'`�4��@N�V4@Bs��!?�FY�]��@��s�ٿ���iL7�@	<��4@�!5mȐ!?hQ\ ��@��s�ٿ���iL7�@	<��4@�!5mȐ!?hQ\ ��@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@����D�ٿ�ՑYs�@瓈��4@G�u���!?US��%-�@*@�mh�ٿ�dC�=�@�z�4@¼&�U�!?1c�k$��@*@�mh�ٿ�dC�=�@�z�4@¼&�U�!?1c�k$��@*@�mh�ٿ�dC�=�@�z�4@¼&�U�!?1c�k$��@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@�H�E�ٿC�.����@��k�4@�w��p�!?z�Zz���@���Ƈٿ�Ag��@!�L�4@��Ϟ\�!?`>S4 �@���ٿ����@
��d4@�(+.��!? [ ���@���ٿ����@
��d4@�(+.��!? [ ���@���ٿ����@
��d4@�(+.��!? [ ���@���ٿ����@
��d4@�(+.��!? [ ���@���ٿ����@
��d4@�(+.��!? [ ���@`��Ai�ٿ����B�@�ڒaB4@�D$�|�!?��dţ�@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@	�Ϫ}ٿ-5֞�@=�X;&4@Ej�#�!?yݡ�z��@_O��yٿ�YO���@��H�4@j�/�9�!?�l���z�@0��t�{ٿp��[��@���4@��y5�!?�B�oS��@0��t�{ٿp��[��@���4@��y5�!?�B�oS��@0��t�{ٿp��[��@���4@��y5�!?�B�oS��@5��~ٿ��$���@&7��4@�ܘ�!?�'\�s
�@5��~ٿ��$���@&7��4@�ܘ�!?�'\�s
�@5��~ٿ��$���@&7��4@�ܘ�!?�'\�s
�@5��~ٿ��$���@&7��4@�ܘ�!?�'\�s
�@褰��}ٿA��%��@�j�I�4@ST\�,�!?�/�����@褰��}ٿA��%��@�j�I�4@ST\�,�!?�/�����@�W^Wp�ٿ� W&@T�@�X�	G4@�;���!?Kv�orz�@�W^Wp�ٿ� W&@T�@�X�	G4@�;���!?Kv�orz�@�W^Wp�ٿ� W&@T�@�X�	G4@�;���!?Kv�orz�@�W^Wp�ٿ� W&@T�@�X�	G4@�;���!?Kv�orz�@�W^Wp�ٿ� W&@T�@�X�	G4@�;���!?Kv�orz�@>�D%�ٿ�^[�}��@�U�#> 4@�*���!?�m���T�@>�D%�ٿ�^[�}��@�U�#> 4@�*���!?�m���T�@>�D%�ٿ�^[�}��@�U�#> 4@�*���!?�m���T�@>�D%�ٿ�^[�}��@�U�#> 4@�*���!?�m���T�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@�����ٿ���|��@o��4@����!? 7��q�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@~~�h��ٿ�I\MY�@`��n�4@����!?xT \N�@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@���O�ٿ�y~h)��@��Z4@d�X���!?M�N����@�o퇈ٿ����@��1�4@�z�H3�!?���O5h�@�o퇈ٿ����@��1�4@�z�H3�!?���O5h�@���=��ٿ$��6��@>T_1@4@-��&2�!?~�ǕiM�@���=��ٿ$��6��@>T_1@4@-��&2�!?~�ǕiM�@�;�Х�ٿe��u�@[2�s�4@t�Y��!?�w�H"��@�;�Х�ٿe��u�@[2�s�4@t�Y��!?�w�H"��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@Tg���ٿQk��@�ǒ޶4@�_�*֐!?9��
��@gp��R�ٿ�_
����@�KZ�4@Dż;��!?2���p�@gp��R�ٿ�_
����@�KZ�4@Dż;��!?2���p�@gp��R�ٿ�_
����@�KZ�4@Dż;��!?2���p�@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@;;�?�ٿv�e��@A�.4@td��!?N��e��@�jf��ٿ��5N��@)g��4@X�{��!?�vB���@��y�F�ٿ�첂��@��ec�4@����%�!?fex1�L�@��y�F�ٿ�첂��@��ec�4@����%�!?fex1�L�@��y�F�ٿ�첂��@��ec�4@����%�!?fex1�L�@��y�F�ٿ�첂��@��ec�4@����%�!?fex1�L�@��	�Ёٿ�Q}NX��@�p(��4@�ͷ��!?�~H⩖�@��	�Ёٿ�Q}NX��@�p(��4@�ͷ��!?�~H⩖�@�ɾLe�ٿ�G��e��@i7�G�4@^%����!?_i�O��@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@�mRٿ�������@��4��4@MR��!?��ª���@4�@�ٿ���)�@��S u4@�����!?�T�w��@4�@�ٿ���)�@��S u4@�����!?�T�w��@4�@�ٿ���)�@��S u4@�����!?�T�w��@4�@�ٿ���)�@��S u4@�����!?�T�w��@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@��I�ٿ�R۵?�@���{n4@��j ��!?	`��B�@Q�{�>�ٿ3��Ť�@V��4@E����!?�Ōr�t�@Q�{�>�ٿ3��Ť�@V��4@E����!?�Ōr�t�@Q�{�>�ٿ3��Ť�@V��4@E����!?�Ōr�t�@Q�{�>�ٿ3��Ť�@V��4@E����!?�Ōr�t�@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@}X'�ٿ��k١��@b�Z4@jp�'��!?����R��@���\�ٿ��j�J��@��?�w4@_TY��!?�^����@���\�ٿ��j�J��@��?�w4@_TY��!?�^����@���\�ٿ��j�J��@��?�w4@_TY��!?�^����@���\�ٿ��j�J��@��?�w4@_TY��!?�^����@<`VU��ٿ�\i/���@а��4@�rؕ��!?&�P�6��@<`VU��ٿ�\i/���@а��4@�rؕ��!?&�P�6��@�Ɲ}%�ٿ�՛3��@�⼲34@}�93��!?b��_l�@�Ɲ}%�ٿ�՛3��@�⼲34@}�93��!?b��_l�@�Ɲ}%�ٿ�՛3��@�⼲34@}�93��!?b��_l�@�Ɲ}%�ٿ�՛3��@�⼲34@}�93��!?b��_l�@�
�>Äٿt1����@C�OF�4@K����!?�IH���@�2�㾇ٿ���R��@D�m��4@�\za!?A6x�O�@�2�㾇ٿ���R��@D�m��4@�\za!?A6x�O�@�2�㾇ٿ���R��@D�m��4@�\za!?A6x�O�@�2�㾇ٿ���R��@D�m��4@�\za!?A6x�O�@�2�㾇ٿ���R��@D�m��4@�\za!?A6x�O�@���ٿ��qЉ�@�ъK4@"����!?ۋܯ���@���ٿ��qЉ�@�ъK4@"����!?ۋܯ���@���ٿ��qЉ�@�ъK4@"����!?ۋܯ���@A&;㹊ٿp2~����@o��*4@��f=Ȑ!?S��x�K�@A&;㹊ٿp2~����@o��*4@��f=Ȑ!?S��x�K�@A&;㹊ٿp2~����@o��*4@��f=Ȑ!?S��x�K�@A&;㹊ٿp2~����@o��*4@��f=Ȑ!?S��x�K�@A&;㹊ٿp2~����@o��*4@��f=Ȑ!?S��x�K�@�*Շٿ�j>=��@��Mh4@��<��!?�7Y����@��p��ٿrcL=8��@%�.��4@3$�9��!?I$��2�@a�	V!�ٿ�uQ��@� `,&4@�Q��p�!?��:��&�@a�	V!�ٿ�uQ��@� `,&4@�Q��p�!?��:��&�@�7~(�ٿ9���@��gB4@EkSQE�!?\��x��@�7~(�ٿ9���@��gB4@EkSQE�!?\��x��@�7~(�ٿ9���@��gB4@EkSQE�!?\��x��@�7~(�ٿ9���@��gB4@EkSQE�!?\��x��@!����{ٿ���j��@I]�I|4@#��A�!?�r���@!����{ٿ���j��@I]�I|4@#��A�!?�r���@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@z�c�ٿ�����@)g��A4@�|��ݐ!?�l�$�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@0�ݙ��ٿX*1L��@�RjS�4@	D�!?m��:�=�@�2��ٿq;�dp��@�ݿV4@�M���!?��z^�@�|�5�ٿ&}'��)�@U�Jx4@���!?B�pLz�@�|�5�ٿ&}'��)�@U�Jx4@���!?B�pLz�@[i�ٿR�ѪW��@F�G=�4@R�y��!?K9k�!��@[i�ٿR�ѪW��@F�G=�4@R�y��!?K9k�!��@[i�ٿR�ѪW��@F�G=�4@R�y��!?K9k�!��@[i�ٿR�ѪW��@F�G=�4@R�y��!?K9k�!��@����@�ٿ�����,�@)��64@��1��!?����/�@����@�ٿ�����,�@)��64@��1��!?����/�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@�h�*Մٿj�6�b��@�~	��4@�lO �!?Њ^0C�@��� !�ٿ�������@��/]4@d�殐!?&
�����@��� !�ٿ�������@��/]4@d�殐!?&
�����@4� �ٿw��]`��@�E�f4@�!v��!?H��I u�@4� �ٿw��]`��@�E�f4@�!v��!?H��I u�@4� �ٿw��]`��@�E�f4@�!v��!?H��I u�@a!��l�ٿ̯a�/�@P!_�4@����А!?���lk�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@'�O���ٿ��Si�l�@�P1�4@���ߺ�!?�N\a�@�����zٿU�bj���@ =)}4@Y8�*��!?���D�!�@�����zٿU�bj���@ =)}4@Y8�*��!?���D�!�@�����zٿU�bj���@ =)}4@Y8�*��!?���D�!�@��մ��ٿ�/�ʉ�@��ʫ4@��{9X�!?��\�#��@��մ��ٿ�/�ʉ�@��ʫ4@��{9X�!?��\�#��@��մ��ٿ�/�ʉ�@��ʫ4@��{9X�!?��\�#��@û�k��ٿ��c���@j�3�/4@{���!?��T?�@û�k��ٿ��c���@j�3�/4@{���!?��T?�@��5�ٿ��'���@��U�i4@�ɟ�!?�W?R3�@��5�ٿ��'���@��U�i4@�ɟ�!?�W?R3�@��5�ٿ��'���@��U�i4@�ɟ�!?�W?R3�@�F���ٿ�y�NE��@�v��@4@��3ѐ!?P/��8��@�F���ٿ�y�NE��@�v��@4@��3ѐ!?P/��8��@�F���ٿ�y�NE��@�v��@4@��3ѐ!?P/��8��@�pz�ٿ<P�����@ [4@l�`�S�!?�)`O���@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@OU�|ٿ��Y�>�@��0��3@@�˭��!?Ϭ����@q5�~*�ٿ$*xq���@�&�4@/�l�!?�^�*P�@q5�~*�ٿ$*xq���@�&�4@/�l�!?�^�*P�@q5�~*�ٿ$*xq���@�&�4@/�l�!?�^�*P�@q5�~*�ٿ$*xq���@�&�4@/�l�!?�^�*P�@־�W�ٿkv�;���@G7��4@�7��!?�z�;+�@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@ɩ���ٿ����q"�@����4@��eۅ�!?(�3M��@y���Ƀٿ)����@�i{�4@=���w�!?{��n��@y���Ƀٿ)����@�i{�4@=���w�!?{��n��@y���Ƀٿ)����@�i{�4@=���w�!?{��n��@k�kc�}ٿ�*Z��@��74@R�����!?^`���@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@؄I3=�ٿ[�k\�@ï�wy4@ַ����!?����D�@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@~r� U�ٿ��J�f�@ys�4@��ɉ�!?L��T��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@�>
�ٿ��<!B��@����t4@�=����!?kc�9k��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@ &Ü�ٿ=I�x_��@�AC�4@)�[���!?]0�N��@�5��N�ٿ2�L�1�@�!�V4@"�a�!?u�~F�6�@�5��N�ٿ2�L�1�@�!�V4@"�a�!?u�~F�6�@�5��N�ٿ2�L�1�@�!�V4@"�a�!?u�~F�6�@�5��N�ٿ2�L�1�@�!�V4@"�a�!?u�~F�6�@�5��N�ٿ2�L�1�@�!�V4@"�a�!?u�~F�6�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@(M2 �ٿ8���M��@@�6�4@��N@��!?B~��x�@�ўf�ٿ�V
���@j����4@Pq�{��!?���ӆ�@�ўf�ٿ�V
���@j����4@Pq�{��!?���ӆ�@�ўf�ٿ�V
���@j����4@Pq�{��!?���ӆ�@$lv=|�ٿ(�f�"K�@��-�4@e7?��!?|&cz�@$lv=|�ٿ(�f�"K�@��-�4@e7?��!?|&cz�@�@�s��ٿ� py�@F()f
4@�]N$5�!?����{�@B+MBc�ٿ����@��!)�	4@��"��!?(��x��@B+MBc�ٿ����@��!)�	4@��"��!?(��x��@B+MBc�ٿ����@��!)�	4@��"��!?(��x��@mu�tM�ٿ!��f�1�@NH�M4@M�?�!?�Y�K�@mu�tM�ٿ!��f�1�@NH�M4@M�?�!?�Y�K�@��:�6�ٿ�Y"w�d�@��hU�4@*���!?��dC�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�����ٿ9��2��@ ���n4@&�q��!?ٟ�-�@�|F(�ٿ�!BS'��@�s_�_4@���U|�!?=.�7���@x����ٿk(]�Ѷ�@�JR�4@%&ECB�!?��`U n�@)]�+�ٿP-���5�@@���
4@�����!?; �L�@)]�+�ٿP-���5�@@���
4@�����!?; �L�@?�]�ٿ%��+:��@a�(4@�|��V�!?`���"�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@��'iɅٿ8`,��@k���24@I��=x�!?Y)@�I�@NW.܃ٿ��	��+�@�5w4@�*��!?�
�)��@NW.܃ٿ��	��+�@�5w4@�*��!?�
�)��@NW.܃ٿ��	��+�@�5w4@�*��!?�
�)��@NW.܃ٿ��	��+�@�5w4@�*��!?�
�)��@+�m~ٿ,-�3���@"j�a4@�q��D�!?h�1�@+�m~ٿ,-�3���@"j�a4@�q��D�!?h�1�@+�m~ٿ,-�3���@"j�a4@�q��D�!?h�1�@+�m~ٿ,-�3���@"j�a4@�q��D�!?h�1�@+�m~ٿ,-�3���@"j�a4@�q��D�!?h�1�@z�h=�ٿO�p���@��~4@��:�,�!?w�$k��@z�h=�ٿO�p���@��~4@��:�,�!?w�$k��@z�h=�ٿO�p���@��~4@��:�,�!?w�$k��@z�h=�ٿO�p���@��~4@��:�,�!?w�$k��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@����}ٿ2kd��@:xO�
4@�t�K�!?Ʌ��+��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@�IO��}ٿ�ؤ�p�@����4@F�q�<�!?����`��@����1�ٿ��@e"��@�c�L�4@�J�#H�!?j#/��Y�@���v��ٿrc8�*��@�q���4@ K�!?D��v���@��GJf�ٿ�ܛXZ��@pH.��4@�Z'b�!?��,���@+?���ٿ9�ƱNW�@ �G�4@ق���!?'�I���@�ǣ�ٿ���!o�@u
E�4@�Qz�א!?��~1���@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@���럇ٿno�(��@��h�0	4@(���!?k���!��@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@�,�*/�ٿ�˱��@w�09Z4@��/У�!?gI�㵶�@��D��ٿ������@rz��4@C�W-��!?������@��D��ٿ������@rz��4@C�W-��!?������@��D��ٿ������@rz��4@C�W-��!?������@��D��ٿ������@rz��4@C�W-��!?������@��D��ٿ������@rz��4@C�W-��!?������@��D��ٿ������@rz��4@C�W-��!?������@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@�'Bi4�ٿyM�̲��@b����4@�����!?C����@a���ٿ=�4&���@~���4@�}5n�!?t�X���@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@��^�ڀٿ�)'c�@Q��� 4@o��ә�!?��)m��@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@=Oo�(�ٿ���բ�@��W9�4@b�����!?{�*���@�TY���ٿaޞO{�@5�Y,4@������!?����F�@�TY���ٿaޞO{�@5�Y,4@������!?����F�@�TY���ٿaޞO{�@5�Y,4@������!?����F�@�TY���ٿaޞO{�@5�Y,4@������!?����F�@�Y��F�ٿ����@��b��4@�F |��!?������@�Y��F�ٿ����@��b��4@�F |��!?������@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@z{O��ٿ7�O�ҭ�@3���c4@���^��!?[����q�@�1�㋂ٿ�~�"�T�@��.��4@WM;��!?��Q���@�1�㋂ٿ�~�"�T�@��.��4@WM;��!?��Q���@�1�㋂ٿ�~�"�T�@��.��4@WM;��!?��Q���@E���ٿ3��F?-�@nk(�y4@f�4��!?;����+�@E���ٿ3��F?-�@nk(�y4@f�4��!?;����+�@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@)7K��ٿ33�4I�@]�\�4@��4���!?�H�[��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@w�v1�ٿ�˴>�W�@Qi�+�4@:.w8��!?��Fe��@ӎ�ٿxrs�a�@�VT�S4@jH���!?,Q���@ӎ�ٿxrs�a�@�VT�S4@jH���!?,Q���@ӎ�ٿxrs�a�@�VT�S4@jH���!?,Q���@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@g����ٿ$[5҂�@`��G�4@⑸&_�!?�ҭ�w��@K�<�4�ٿK	�W��@qx��d4@z�c1I�!?�*��k�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@~�&���ٿ�W� ��@����	4@4xfޙ�!?��*S�@wnaz�ٿL��Є�@�Y7_�4@�Hm��!?����@wnaz�ٿL��Є�@�Y7_�4@�Hm��!?����@wnaz�ٿL��Є�@�Y7_�4@�Hm��!?����@wnaz�ٿL��Є�@�Y7_�4@�Hm��!?����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@�r����ٿ�_\�q�@��Ziw4@�^M���!?:L����@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@��R��ٿ�D�]u�@�u��4@=b�ɐ!?�az[�`�@OK+���ٿ �e	2��@�V�A4@O	���!?&���ު�@OK+���ٿ �e	2��@�V�A4@O	���!?&���ު�@�C]�ٿ<�r"���@�>"E4@c^+��!?Ka-QX�@�C]�ٿ<�r"���@�>"E4@c^+��!?Ka-QX�@�C]�ٿ<�r"���@�>"E4@c^+��!?Ka-QX�@�C]�ٿ<�r"���@�>"E4@c^+��!?Ka-QX�@���3�ٿȺD6��@g
�4@��N<��!?-��L��@���3�ٿȺD6��@g
�4@��N<��!?-��L��@���3�ٿȺD6��@g
�4@��N<��!?-��L��@���3�ٿȺD6��@g
�4@��N<��!?-��L��@���3�ٿȺD6��@g
�4@��N<��!?-��L��@I4��҇ٿS�)N+��@5���d�3@~\��ΐ!?�ȸ9���@I4��҇ٿS�)N+��@5���d�3@~\��ΐ!?�ȸ9���@(����ٿ:o�`9�@�����4@e�8�Ӑ!?cAԒP@�@(����ٿ:o�`9�@�����4@e�8�Ӑ!?cAԒP@�@(����ٿ:o�`9�@�����4@e�8�Ӑ!?cAԒP@�@(����ٿ:o�`9�@�����4@e�8�Ӑ!?cAԒP@�@(����ٿ:o�`9�@�����4@e�8�Ӑ!?cAԒP@�@z��ٿxߘ���@��/�� 4@n�N,"�!?�C���@z��ٿxߘ���@��/�� 4@n�N,"�!?�C���@x=
�b�ٿ��N��@#�R}��3@�+���!?�r�����@x=
�b�ٿ��N��@#�R}��3@�+���!?�r�����@��ۅٿ�O�%��@W:e^�4@�xvb�!?�r��=��@T�_�~ٿ{*��M�@�J�=�4@:�'^J�!?����@T�_�~ٿ{*��M�@�J�=�4@:�'^J�!?����@T�_�~ٿ{*��M�@�J�=�4@:�'^J�!?����@T�_�~ٿ{*��M�@�J�=�4@:�'^J�!?����@T�_�~ٿ{*��M�@�J�=�4@:�'^J�!?����@�>�1�ٿ��f���@��}�4@��t͐!?���W��@�>�1�ٿ��f���@��}�4@��t͐!?���W��@jm��|ٿ�"%���@��/3�4@�i���!?�������@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@P�Ɂ�ٿ#9����@�[У4@�+pL�!?����@��Y��ٿ n���2�@Ͱ:y�4@H�H0�!?ȡ҈j�@��Y��ٿ n���2�@Ͱ:y�4@H�H0�!?ȡ҈j�@ދ�z��ٿ�TX.f�@4Ӛ�4@Q��Đ!?<�=� �@ދ�z��ٿ�TX.f�@4Ӛ�4@Q��Đ!?<�=� �@��z��ٿ��O���@�L�4@A���!?*x���@��z��ٿ��O���@�L�4@A���!?*x���@��z��ٿ��O���@�L�4@A���!?*x���@��z��ٿ��O���@�L�4@A���!?*x���@�/���ٿKLM��T�@L��(04@�0�#��!?�z���@�/���ٿKLM��T�@L��(04@�0�#��!?�z���@�/���ٿKLM��T�@L��(04@�0�#��!?�z���@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@c9�y �ٿ��[��@���ܯ4@�0�]�!?WNZ�p�@ɡ��c�ٿo5w���@����4@�͇��!?����j�@ɡ��c�ٿo5w���@����4@�͇��!?����j�@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@�O\�ٿ�h� �k�@;����4@;���!?5������@5��ٿ�����v�@�¦�d4@7)Ő!?� ��*�@5��ٿ�����v�@�¦�d4@7)Ő!?� ��*�@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@�ݤ�Ɋٿ�8D6���@�W֧N4@WK{�w�!?��~)��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@��1�e�ٿw�ءq(�@�c_ 	4@A�a k�!?&��O��@B@K�ٿ�
�g���@S,(�4@�+�q�!?&���i��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@.)���ٿ���#U�@x93� 4@K��I��!?�SV$��@�.��^�ٿ�[���@M��{4@�e_�Ð!?��8��@���d��ٿ��<��@{���4@K����!?�f�*8F�@�����~ٿ%�Wj2��@����4@d8����!?����#k�@�����~ٿ%�Wj2��@����4@d8����!?����#k�@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@� l���ٿ'���R�@��D�4@p����!?&09���@��Yw�ٿq�Om�>�@;EtШ4@᳅���!?��9/�@�ݠ瞃ٿ��$��@?'��a	4@��H'ѐ!?b�y��D�@�p���ٿW�+�ڦ�@�YC��	4@����ڐ!?���\.�@�p���ٿW�+�ڦ�@�YC��	4@����ڐ!?���\.�@�����ٿ'�.�b�@3~��4@4����!?�NM<7�@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@��!�ٿ�g�U��@z��4@�cz�!?�EQ�W��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@�h�|ٿɒ�F�A�@�/��4@��S-��!?�dvWe��@~&rY�vٿD=�7��@����|4@"���2�!?�-d	��@~&rY�vٿD=�7��@����|4@"���2�!?�-d	��@	�]|ٿ�ߍ��_�@�;g�_4@4!��S�!?���>�@	�]|ٿ�ߍ��_�@�;g�_4@4!��S�!?���>�@\n�MY�ٿ8����@�ٰ�4@�G�۵�!?����:�@¾KDZ�ٿ��ܕ���@�kv��4@ķ��Ȑ!?+���,�@¾KDZ�ٿ��ܕ���@�kv��4@ķ��Ȑ!?+���,�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@��`���ٿ>O���@�ϴ[! 4@��ٯ^�!?��@�:W�@A�pĀٿ9Υ�g�@��o�4@sŢ�!?��<|�@A�pĀٿ9Υ�g�@��o�4@sŢ�!?��<|�@A�pĀٿ9Υ�g�@��o�4@sŢ�!?��<|�@�����ٿ���1,v�@'��$�4@aJ*�v�!?�=:��@�_��~ٿK+S����@�sC� 4@�]���!?�c�&��@�_��~ٿK+S����@�sC� 4@�]���!?�c�&��@�_��~ٿK+S����@�sC� 4@�]���!?�c�&��@�_��~ٿK+S����@�sC� 4@�]���!?�c�&��@14�i�ٿ���]���@,�&�4@��zF�!?�剛A�@~�(�ٌٿ��@���@����4@G6�ӗ�!?A_��)��@~�(�ٌٿ��@���@����4@G6�ӗ�!?A_��)��@~�(�ٌٿ��@���@����4@G6�ӗ�!?A_��)��@~�(�ٌٿ��@���@����4@G6�ӗ�!?A_��)��@:�Lفٿ;bPTSy�@Xg��4@m�:��!?��P?I��@�� �ȁٿ��6���@���@4@}>+�!?Χ*e��@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�i�Dh�ٿ�2h,��@)e��4@֠�h�!?31`Lq�@�����ٿ�nx�n�@��Oa}4@챹�r�!?P�υY�@�����ٿ�nx�n�@��Oa}4@챹�r�!?P�υY�@�����ٿ�nx�n�@��Oa}4@챹�r�!?P�υY�@�����ٿ�nx�n�@��Oa}4@챹�r�!?P�υY�@�S����ٿ\bݿi?�@j��}�4@Q�׎��!?���f���@�S����ٿ\bݿi?�@j��}�4@Q�׎��!?���f���@�S����ٿ\bݿi?�@j��}�4@Q�׎��!?���f���@�S����ٿ\bݿi?�@j��}�4@Q�׎��!?���f���@�
S�i�ٿ�Jq���@+v�� 4@X�E���!?�K��G�@�
S�i�ٿ�Jq���@+v�� 4@X�E���!?�K��G�@M���ٿ=�ҺiR�@�g��/�3@ŪN�!?�b-=͔�@M���ٿ=�ҺiR�@�g��/�3@ŪN�!?�b-=͔�@M���ٿ=�ҺiR�@�g��/�3@ŪN�!?�b-=͔�@M���ٿ=�ҺiR�@�g��/�3@ŪN�!?�b-=͔�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@}ASa�ٿ�޽���@�חG��3@i6��ݐ!?i~���U�@,۪��ٿ"���qf�@�6
�M4@���\��!?H!�I-�@,۪��ٿ"���qf�@�6
�M4@���\��!?H!�I-�@,۪��ٿ"���qf�@�6
�M4@���\��!?H!�I-�@,۪��ٿ"���qf�@�6
�M4@���\��!?H!�I-�@,۪��ٿ"���qf�@�6
�M4@���\��!?H!�I-�@�L�M�ٿw9q�sC�@��-u�4@xD����!?�UDB��@�L�M�ٿw9q�sC�@��-u�4@xD����!?�UDB��@�G�U�ٿÔ1>��@�1���4@Ƴ����!?�[�"�@�G�U�ٿÔ1>��@�1���4@Ƴ����!?�[�"�@�G�U�ٿÔ1>��@�1���4@Ƴ����!?�[�"�@��f��ٿ��"q)�@�9?E4@P~��d�!?� ��@���c�ٿћe<2�@F�]4@B_Bك�!?��v�c��@v�@��ٿɫ�dr�@���4@�p����!?s�,�<�@T�����ٿ,風C�@��{:4@0�Z]�!?n���@T�����ٿ,風C�@��{:4@0�Z]�!?n���@T�����ٿ,風C�@��{:4@0�Z]�!?n���@T�����ٿ,風C�@��{:4@0�Z]�!?n���@T�����ٿ,風C�@��{:4@0�Z]�!?n���@T�����ٿ,風C�@��{:4@0�Z]�!?n���@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@S���ٿ���W�i�@Oi{�4@P:�ݐ!?
�U�Ơ�@��E��ٿC�җ�@ ���Q4@y��q�!?㕲���@��E��ٿC�җ�@ ���Q4@y��q�!?㕲���@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@x�"�1�ٿ�F�p�@b���q4@U�u�!?)RQ%�@�WR?�ٿ����@+g�:h4@�W��!?�"���@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@4�����ٿ%[c+r�@���̚4@9ن��!?o�a-�^�@X����ٿ��[�5��@$��u�4@HTAQ��!?h�1Ǩ�@X����ٿ��[�5��@$��u�4@HTAQ��!?h�1Ǩ�@%�<;��ٿ��Ge��@Q�c�-4@f�$�n�!?n���3��@%�<;��ٿ��Ge��@Q�c�-4@f�$�n�!?n���3��@%�<;��ٿ��Ge��@Q�c�-4@f�$�n�!?n���3��@������ٿ�(;.0�@�∮�4@-��AȐ!?TP�k�&�@�c-��ٿ�:.*E�@�W���4@Z�<ː!?��8 �P�@��o�y�ٿ�!T89�@^�ԏ�4@Q�����!?�0����@��o�y�ٿ�!T89�@^�ԏ�4@Q�����!?�0����@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@�Om��{ٿU}���@Y�a��4@x�A��!?��`��@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@���Ӂٿ��u
�@W䍼4@�*<3��!?����ŷ�@������ٿ�J�X��@� ��4@1˟���!?�c`���@������ٿ�J�X��@� ��4@1˟���!?�c`���@������ٿ�J�X��@� ��4@1˟���!?�c`���@������ٿ�J�X��@� ��4@1˟���!?�c`���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@/srԑٿ�(D-4��@U��4@49��!?Fi���@��V�Ȋٿ}�A���@�G�~]4@-�4�!?��F8��@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�c�ՇٿU���EL�@4\�G4@��*:�!?�#���@�a��,�ٿ�uܭ͢�@j�/8�4@OJ�Ő�!?Ɗ,���@����y�ٿ���ӫ��@A��(�4@mB2��!?]��F��@����y�ٿ���ӫ��@A��(�4@mB2��!?]��F��@��/��ٿ�x��Ǿ�@j[�ϥ4@z�a�!?D�Dז4�@��/��ٿ�x��Ǿ�@j[�ϥ4@z�a�!?D�Dז4�@��/��ٿ�x��Ǿ�@j[�ϥ4@z�a�!?D�Dז4�@��/��ٿ�x��Ǿ�@j[�ϥ4@z�a�!?D�Dז4�@�C=偊ٿQ��Il��@�6��34@�Şc3�!?��X��@u��}�ٿyk]Y�!�@�'�K4@L�=��!?ۿ�z�8�@u��}�ٿyk]Y�!�@�'�K4@L�=��!?ۿ�z�8�@� ���ٿ�m�y8��@G�&�4@�x���!?[�p�@��R�ٿ��,� ��@Ɇ<�V4@���(��!?��
���@\*���ٿ6�E��@�P=	4@�$��!?�����	�@\*���ٿ6�E��@�P=	4@�$��!?�����	�@\*���ٿ6�E��@�P=	4@�$��!?�����	�@\*���ٿ6�E��@�P=	4@�$��!?�����	�@\*���ٿ6�E��@�P=	4@�$��!?�����	�@\*���ٿ6�E��@�P=	4@�$��!?�����	�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@��K�ٿ
�Į���@��C4@�r��a�!?�,Uv̬�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@J�'�>�ٿ/�i�:��@K����4@�$���!?���^�J�@�2@|�ٿ�g�@R6�`�4@����q�!?Q|�g��@�2@|�ٿ�g�@R6�`�4@����q�!?Q|�g��@�2@|�ٿ�g�@R6�`�4@����q�!?Q|�g��@�2@|�ٿ�g�@R6�`�4@����q�!?Q|�g��@1� ��|ٿi:��@���4@��"P�!?2�S�k��@1� ��|ٿi:��@���4@��"P�!?2�S�k��@1� ��|ٿi:��@���4@��"P�!?2�S�k��@1� ��|ٿi:��@���4@��"P�!?2�S�k��@1� ��|ٿi:��@���4@��"P�!?2�S�k��@��q��vٿ�Sh>�@�r�9(4@���V��!?��0�d�@�����zٿ��$�{��@�Vtl}4@�l!��!?E�]���@�����zٿ��$�{��@�Vtl}4@�l!��!?E�]���@�����zٿ��$�{��@�Vtl}4@�l!��!?E�]���@w�6�ٿߌ��=!�@�:K�T4@>*��ސ!?:c���@w�6�ٿߌ��=!�@�:K�T4@>*��ސ!?:c���@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@{̧m+�ٿ4��,k9�@��"��4@B9����!?���M�Y�@a�=l�ٿUl�!?�@=����4@��%O��!?��	��@a�=l�ٿUl�!?�@=����4@��%O��!?��	��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��;D_�ٿ�*���@�@X�4@h�����!?a��I��@��C�R�ٿ���1|�@_hkw� 4@�:����!?�"� j�@@�Bn�ٿ�m�����@gé�� 4@�IC#'�!?�LY����@@�Bn�ٿ�m�����@gé�� 4@�IC#'�!?�LY����@@�Bn�ٿ�m�����@gé�� 4@�IC#'�!?�LY����@@�Bn�ٿ�m�����@gé�� 4@�IC#'�!?�LY����@@�Bn�ٿ�m�����@gé�� 4@�IC#'�!?�LY����@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@��_̈ٿ5�n��@�/-5�3@�j1��!?�j�*�@���Y�ٿ��mj
�@y��!�3@f	J���!?�u:4��@���Y�ٿ��mj
�@y��!�3@f	J���!?�u:4��@���Y�ٿ��mj
�@y��!�3@f	J���!?�u:4��@���Y�ٿ��mj
�@y��!�3@f	J���!?�u:4��@/���ٿ�',�T��@f���q�3@�s�o�!?�Z�Ӯ�@/���ٿ�',�T��@f���q�3@�s�o�!?�Z�Ӯ�@/���ٿ�',�T��@f���q�3@�s�o�!?�Z�Ӯ�@ "9�V�ٿ[u%R��@n���j4@�pk7��!?1�m��@ "9�V�ٿ[u%R��@n���j4@�pk7��!?1�m��@ "9�V�ٿ[u%R��@n���j4@�pk7��!?1�m��@ "9�V�ٿ[u%R��@n���j4@�pk7��!?1�m��@ "9�V�ٿ[u%R��@n���j4@�pk7��!?1�m��@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@/�uH0�ٿ}���C�@;׃;4@+F|͐!?u���t�@����z�ٿ��.�/�@��f&�4@��sՐ!?D��U���@����z�ٿ��.�/�@��f&�4@��sՐ!?D��U���@(it�4�ٿ	�ۖ���@zn�/4@���.�!?z����@(it�4�ٿ	�ۖ���@zn�/4@���.�!?z����@(it�4�ٿ	�ۖ���@zn�/4@���.�!?z����@��ó��ٿw�Η��@���a4@�����!?�]�q��@��ó��ٿw�Η��@���a4@�����!?�]�q��@��ó��ٿw�Η��@���a4@�����!?�]�q��@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@^��3Ҋٿ���8��@�"�<�4@����ؐ!?-��B�@8d8�X�ٿ�I���@�H	-
4@e^�!?n�#n���@8d8�X�ٿ�I���@�H	-
4@e^�!?n�#n���@2���ٿ�0�'{��@o���|4@����!?��I�:�@2���ٿ�0�'{��@o���|4@����!?��I�:�@2���ٿ�0�'{��@o���|4@����!?��I�:�@e��\�ٿ��N뛷�@F�j�	4@<�V��!?x���xz�@e��\�ٿ��N뛷�@F�j�	4@<�V��!?x���xz�@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@���ٿK.��"�@$�l[`4@S��Lِ!?CN$���@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@]/�\^�ٿQ)����@v�\4@�\�鱐!?j��}�	�@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@\�fo%�ٿ i�L0�@���4@C����!?;���@Q8� ��ٿ�1dW�d�@�E� 4@C���ܐ!?͉Y^��@sq��ٿkE�Lm�@���1|4@���ِ!?���M%��@sq��ٿkE�Lm�@���1|4@���ِ!?���M%��@sq��ٿkE�Lm�@���1|4@���ِ!?���M%��@sq��ٿkE�Lm�@���1|4@���ِ!?���M%��@sq��ٿkE�Lm�@���1|4@���ِ!?���M%��@Y>R]�ٿ3�Tk���@�Ǳ�4@9J��Ԑ!?�r�S�N�@Y>R]�ٿ3�Tk���@�Ǳ�4@9J��Ԑ!?�r�S�N�@Y>R]�ٿ3�Tk���@�Ǳ�4@9J��Ԑ!?�r�S�N�@Y>R]�ٿ3�Tk���@�Ǳ�4@9J��Ԑ!?�r�S�N�@�ӎ�1�ٿܫ��z"�@�]8�4@�w����!?̡����@��3�V�ٿ�C�\��@
􁻆4@k"�I��!?(ޥA%�@��3�V�ٿ�C�\��@
􁻆4@k"�I��!?(ޥA%�@��3�V�ٿ�C�\��@
􁻆4@k"�I��!?(ޥA%�@��3�V�ٿ�C�\��@
􁻆4@k"�I��!?(ޥA%�@��3�V�ٿ�C�\��@
􁻆4@k"�I��!?(ޥA%�@��0��ٿr���X��@�����4@��(���!?��#�P��@��0��ٿr���X��@�����4@��(���!?��#�P��@��0��ٿr���X��@�����4@��(���!?��#�P��@PP՝h�ٿ�ҧ9��@�ʚ8�4@e��!?�Y`�=��@PP՝h�ٿ�ҧ9��@�ʚ8�4@e��!?�Y`�=��@PP՝h�ٿ�ҧ9��@�ʚ8�4@e��!?�Y`�=��@PP՝h�ٿ�ҧ9��@�ʚ8�4@e��!?�Y`�=��@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@��jM�ٿ�-&,��@I�8#4@w�x��!?�]Dp�K�@"�E���ٿ��Ft�.�@���U�4@�b���!?G��d��@"�E���ٿ��Ft�.�@���U�4@�b���!?G��d��@"�E���ٿ��Ft�.�@���U�4@�b���!?G��d��@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@>r�}W�ٿ[_�ɀ��@�A�F�4@�>����!?GU�����@W�ĆٿsK�����@���< 4@}��<��!?�Nޠ_�@|��)D�ٿ.�(����@1����4@��v� �!?�'��o�@|��)D�ٿ.�(����@1����4@��v� �!?�'��o�@|��)D�ٿ.�(����@1����4@��v� �!?�'��o�@|��)D�ٿ.�(����@1����4@��v� �!?�'��o�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�R#}8�ٿ_�����@	� 4@#�@���!?�Ԑ��T�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@�s����ٿf�(�@��.8�4@TH{E��!?�����9�@Kj��ٿ���#n*�@�K#�U4@��D+��!?����d�@Kj��ٿ���#n*�@�K#�U4@��D+��!?����d�@Kj��ٿ���#n*�@�K#�U4@��D+��!?����d�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@�CQ�ٿ���d�@m�q4@�v{�ː!?���,�@E^���ٿ[k�c�@�~�TR4@�J��!?�W���@E^���ٿ[k�c�@�~�TR4@�J��!?�W���@g���)�ٿ�w�n;�@Y�S�4@��k{2�!?�^Y)��@ha�t�~ٿ��Fed�@z��k4@��;�!?���d��@ha�t�~ٿ��Fed�@z��k4@��;�!?���d��@ha�t�~ٿ��Fed�@z��k4@��;�!?���d��@ha�t�~ٿ��Fed�@z��k4@��;�!?���d��@ha�t�~ٿ��Fed�@z��k4@��;�!?���d��@~��F�ٿ~���H�@�2'P�4@<�=-�!?���PsB�@~��F�ٿ~���H�@�2'P�4@<�=-�!?���PsB�@~��F�ٿ~���H�@�2'P�4@<�=-�!?���PsB�@~��F�ٿ~���H�@�2'P�4@<�=-�!?���PsB�@��_ۉٿ�ꝝ.��@j4$� 4@TU���!?�$�$��@��_ۉٿ�ꝝ.��@j4$� 4@TU���!?�$�$��@��_ۉٿ�ꝝ.��@j4$� 4@TU���!?�$�$��@��_ۉٿ�ꝝ.��@j4$� 4@TU���!?�$�$��@���ԊٿI�>w��@�Q�;�4@i��f �!?�c2=2R�@���ԊٿI�>w��@�Q�;�4@i��f �!?�c2=2R�@���ԊٿI�>w��@�Q�;�4@i��f �!?�c2=2R�@���ԊٿI�>w��@�Q�;�4@i��f �!?�c2=2R�@Jh�r��ٿ01���@P���4@݆dk��!?Wk~���@Jh�r��ٿ01���@P���4@݆dk��!?Wk~���@Jh�r��ٿ01���@P���4@݆dk��!?Wk~���@Jh�r��ٿ01���@P���4@݆dk��!?Wk~���@\0���|ٿ�ůpU�@	m�4@��B�̐!?%z����@\0���|ٿ�ůpU�@	m�4@��B�̐!?%z����@�`D���ٿa��p�@�nή 4@<t��!?�i����@�`D���ٿa��p�@�nή 4@<t��!?�i����@�`D���ٿa��p�@�nή 4@<t��!?�i����@�`D���ٿa��p�@�nή 4@<t��!?�i����@b���ٿ*&����@�4S�4@�MF�!?�-�c+��@	P���ٿ��؞��@~��q.4@���%�!?��@&�@	P���ٿ��؞��@~��q.4@���%�!?��@&�@	P���ٿ��؞��@~��q.4@���%�!?��@&�@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@g �U �ٿCt��@����4@��?�ΐ!?]�6����@�(�G��ٿ<�Pl���@�-�M�4@�z�!?�4� �@�(�G��ٿ<�Pl���@�-�M�4@�z�!?�4� �@�(�G��ٿ<�Pl���@�-�M�4@�z�!?�4� �@�Р���ٿ%!k#��@�iZ��4@e�e
�!?EHB����@�Р���ٿ%!k#��@�iZ��4@e�e
�!?EHB����@�Р���ٿ%!k#��@�iZ��4@e�e
�!?EHB����@�Р���ٿ%!k#��@�iZ��4@e�e
�!?EHB����@-�1M�ٿ.̔���@�Z5(4@��=z��!?�����@-�1M�ٿ.̔���@�Z5(4@��=z��!?�����@-�1M�ٿ.̔���@�Z5(4@��=z��!?�����@-�1M�ٿ.̔���@�Z5(4@��=z��!?�����@-�1M�ٿ.̔���@�Z5(4@��=z��!?�����@&e)�ٿ��#���@��lb4@�
��!?�O�(��@�j#|iٿS)y��f�@頾/4@�i��Ґ!?�ױ6^�@�j#|iٿS)y��f�@頾/4@�i��Ґ!?�ױ6^�@�j#|iٿS)y��f�@頾/4@�i��Ґ!?�ױ6^�@���(�ٿ�\W����@5�`(p4@Y��N�!?P�n"r��@���(�ٿ�\W����@5�`(p4@Y��N�!?P�n"r��@���(�ٿ�\W����@5�`(p4@Y��N�!?P�n"r��@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@n_u(�ٿu�\���@���4@R�P��!?�'k��>�@����2�ٿ3ɜ,.��@I����4@`�qm�!?
����@����2�ٿ3ɜ,.��@I����4@`�qm�!?
����@����2�ٿ3ɜ,.��@I����4@`�qm�!?
����@����2�ٿ3ɜ,.��@I����4@`�qm�!?
����@ݘ���ٿ��5�p��@o��4@j�b���!?p#���R�@ݘ���ٿ��5�p��@o��4@j�b���!?p#���R�@ݘ���ٿ��5�p��@o��4@j�b���!?p#���R�@ݘ���ٿ��5�p��@o��4@j�b���!?p#���R�@ݘ���ٿ��5�p��@o��4@j�b���!?p#���R�@�5����ٿ�bR�@(���4@V�<w��!? <|'�`�@�5����ٿ�bR�@(���4@V�<w��!? <|'�`�@�5����ٿ�bR�@(���4@V�<w��!? <|'�`�@�5����ٿ�bR�@(���4@V�<w��!? <|'�`�@�5����ٿ�bR�@(���4@V�<w��!? <|'�`�@t��ٿ������@��,b4@x�R�!?E���[�@t��ٿ������@��,b4@x�R�!?E���[�@]L�q�ٿD�9���@Y
D{4@�?ް��!?��(���@W��p[�ٿBJi����@�]�"�4@�egJ̐!?)����'�@W��p[�ٿBJi����@�]�"�4@�egJ̐!?)����'�@��)n�ٿ	�rv��@l,��4@�T�$��!?^x��!�@��)n�ٿ	�rv��@l,��4@�T�$��!?^x��!�@��)n�ٿ	�rv��@l,��4@�T�$��!?^x��!�@E��Ćٿ�j$:�h�@�@_n4@kh�Ґ!?<�=EO��@E��Ćٿ�j$:�h�@�@_n4@kh�Ґ!?<�=EO��@aZ|p��ٿW��9|�@�n�*4@�{+��!?Ev<}��@|x�Z�ٿiqU��j�@�z��4@�9+Đ!?�����@|x�Z�ٿiqU��j�@�z��4@�9+Đ!?�����@|x�Z�ٿiqU��j�@�z��4@�9+Đ!?�����@|x�Z�ٿiqU��j�@�z��4@�9+Đ!?�����@|x�Z�ٿiqU��j�@�z��4@�9+Đ!?�����@�2�ٿd��]G�@8�8l24@��|uƐ!?�V����@�2�ٿd��]G�@8�8l24@��|uƐ!?�V����@�2�ٿd��]G�@8�8l24@��|uƐ!?�V����@�b�,j�ٿ�S�w���@Ht~��4@�q���!?�_E)Z�@�b�,j�ٿ�S�w���@Ht~��4@�q���!?�_E)Z�@�b�,j�ٿ�S�w���@Ht~��4@�q���!?�_E)Z�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@��o�ٿ!�yb�@>RQQ 4@��v���!?^,UPi�@>����ٿf�B���@D��Y� 4@=�@���!?���dh��@>����ٿf�B���@D��Y� 4@=�@���!?���dh��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@���F��ٿ�b2a�_�@�<x�4@ȦX�!?���u��@�nD3r�ٿ��y��o�@�X�%4@w9^z�!?l��H�w�@�nD3r�ٿ��y��o�@�X�%4@w9^z�!?l��H�w�@�nD3r�ٿ��y��o�@�X�%4@w9^z�!?l��H�w�@�nD3r�ٿ��y��o�@�X�%4@w9^z�!?l��H�w�@�nD3r�ٿ��y��o�@�X�%4@w9^z�!?l��H�w�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@Zu�Ar�ٿS�]��@bMz�4@`�wI��!?<m`L׻�@���ٿ�TG��@[���4@�� �!?�M�T���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@7�#�ٿx+���@��)4@t}S�א!?�,�G���@���$-�ٿʖO���@̡2�4@Sц���!?�� ���@���$-�ٿʖO���@̡2�4@Sц���!?�� ���@���$-�ٿʖO���@̡2�4@Sц���!?�� ���@����ٿn������@�Pb�4@dԙ1̐!?�c�a���@����ٿn������@�Pb�4@dԙ1̐!?�c�a���@���O�ٿnDF2�*�@X���!4@���<�!?���a���@���O�ٿnDF2�*�@X���!4@���<�!?���a���@���O�ٿnDF2�*�@X���!4@���<�!?���a���@����ٿ��L�i�@?�r��4@\	�Đ!?l�D;E�@����ٿ��L�i�@?�r��4@\	�Đ!?l�D;E�@3EǏ��ٿ�I��!�@��h�]4@B�c�!?���?��@X�L�ٿ�d����@�/�.	4@Q Q��!?􏥃(��@X�L�ٿ�d����@�/�.	4@Q Q��!?􏥃(��@X�L�ٿ�d����@�/�.	4@Q Q��!?􏥃(��@*����ٿ�ϐK2�@�k?��4@s����!?%��܇�@*����ٿ�ϐK2�@�k?��4@s����!?%��܇�@*����ٿ�ϐK2�@�k?��4@s����!?%��܇�@j$n�2�ٿV��W�i�@���b�4@G%e��!?6�z�
�@x���!�ٿ��|��]�@[�آ	4@�7#���!?KC����@x���!�ٿ��|��]�@[�آ	4@�7#���!?KC����@�I�;!�ٿ�wp�V��@����4@O�t���!?dԻ�%�@�I�;!�ٿ�wp�V��@����4@O�t���!?dԻ�%�@"O駴�ٿ|��n��@Xs.�
4@pf��ΐ!?j�0�@"O駴�ٿ|��n��@Xs.�
4@pf��ΐ!?j�0�@"O駴�ٿ|��n��@Xs.�
4@pf��ΐ!?j�0�@��t�ڈٿP���@ �؏�	4@�e�Ő!?,����:�@��t�ڈٿP���@ �؏�	4@�e�Ő!?,����:�@��t�ڈٿP���@ �؏�	4@�e�Ő!?,����:�@T/5ѻ�ٿQl� l�@�;��4@
�R��!?�#�}��@�-���ٿ�s1��@`ZZgb4@�a@;��!?��L[���@�-���ٿ�s1��@`ZZgb4@�a@;��!?��L[���@�-���ٿ�s1��@`ZZgb4@�a@;��!?��L[���@�-���ٿ�s1��@`ZZgb4@�a@;��!?��L[���@���rN�ٿ6��%�@0�=O4@^��ߐ!?<�<���@���rN�ٿ6��%�@0�=O4@^��ߐ!?<�<���@���rN�ٿ6��%�@0�=O4@^��ߐ!?<�<���@���rN�ٿ6��%�@0�=O4@^��ߐ!?<�<���@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@�1�O�ٿ׎H<L��@����4@�S�&�!?�.eE'�@R:�q�ٿg������@�*�ţ4@bc�cߐ!?�<�<��@������ٿ����@�UZ 4@D�͙�!?�J3����@������ٿ����@�UZ 4@D�͙�!?�J3����@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@D�?�N{ٿ]B:Kq��@�A���4@~k��Đ!?$l�Z�@�����ٿw��|��@M���`4@s�g��!?]�d��	�@X�1�e�ٿ>:���c�@A�!�4@��zʸ�!?ei����@�;��~�ٿ��`��@�(��w4@,��A��!?���%��@�q�*�ٿ�fF{� �@�?`tH4@^��M��!?y�BMH��@�q�*�ٿ�fF{� �@�?`tH4@^��M��!?y�BMH��@�q�*�ٿ�fF{� �@�?`tH4@^��M��!?y�BMH��@�q�*�ٿ�fF{� �@�?`tH4@^��M��!?y�BMH��@�q�*�ٿ�fF{� �@�?`tH4@^��M��!?y�BMH��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@&_{��ٿ�T���@�.��4@t�F�!?��;, ��@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�NÇٿ(�E��-�@�d4@�Z���!?�5�I�0�@�\�Յٿ�NzQ�E�@��4@�s�9!?����9��@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@��ɿ�ٿ���c5�@�f�Ճ	4@+ޡ��!?Ē�Nǵ�@%��ϱ�ٿ3��n6�@�f�`�	4@~&6\֐!?�շ5��@%��ϱ�ٿ3��n6�@�f�`�	4@~&6\֐!?�շ5��@%��ϱ�ٿ3��n6�@�f�`�	4@~&6\֐!?�շ5��@��tT��ٿ,d��%�@w�76�4@!�x��!?�o�-�)�@��tT��ٿ,d��%�@w�76�4@!�x��!?�o�-�)�@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�5۠�ٿ-�D��"�@3ξ4�	4@�� �!?�:F��@�	L�/�ٿ�b�}!�@�_,�|4@�i޺�!? p�����@�	L�/�ٿ�b�}!�@�_,�|4@�i޺�!? p�����@���uˏٿr�Q�W\�@��xF<4@��d��!?���3��@���uˏٿr�Q�W\�@��xF<4@��d��!?���3��@s�'�Dٿ	]����@&�(�J4@�8W�!?wMJ����@A�0�ٿJ`����@ȴ���3@2u˕�!?���c��@��lN��ٿ��N>S��@��H� 4@Ej�!?:�'��e�@8�'�A�ٿ�Pp����@��j��4@G6����!?3�DE#��@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�'v"��ٿ�Dl���@#Ú�* 4@s?��!?Ys0���@�B1�ٿ)0x�)�@3�I��3@J�و�!?�=�Sx�@�\^��ٿ(���2�@DK�}4@�-���!?�#��@�\^��ٿ(���2�@DK�}4@�-���!?�#��@	�K���ٿ���J�@�fiC	4@D���ϐ!?�4j�1�@�+4��}ٿ� ��&�@(W��	4@��Xj�!?�?��:>�@�+4��}ٿ� ��&�@(W��	4@��Xj�!?�?��:>�@L����ٿ�,��h�@�~$ 	4@�O���!?_�gTv0�@y2&R�ٿA���i�@Փ�P'4@uB�%��!?<���lX�@y2&R�ٿA���i�@Փ�P'4@uB�%��!?<���lX�@y2&R�ٿA���i�@Փ�P'4@uB�%��!?<���lX�@y2&R�ٿA���i�@Փ�P'4@uB�%��!?<���lX�@�#����ٿkzWh/C�@9���4@�'�8�!?�0�"���@�#����ٿkzWh/C�@9���4@�'�8�!?�0�"���@�#����ٿkzWh/C�@9���4@�'�8�!?�0�"���@�#����ٿkzWh/C�@9���4@�'�8�!?�0�"���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@��k�,�ٿ�vYz&�@�_�B4@�mŐ!?Դ�t���@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@�qD��ٿ������@���Ѫ4@���ݐ!?R��&(N�@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@n�2��ٿe�ka(�@�݋�4@1T"oِ!?��k}���@�Tht��ٿ��Q�{�@�ﭢ�4@���ǐ!?qo����@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@lx�;B�ٿ�߅�9�@�F��~4@9t���!?���4Fs�@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�r�<��ٿ��M�*�@⁧��4@�CJ���!?U����@�G���ٿV��^��@[@�4@��� Ґ!?{����@�G���ٿV��^��@[@�4@��� Ґ!?{����@�G���ٿV��^��@[@�4@��� Ґ!?{����@�G���ٿV��^��@[@�4@��� Ґ!?{����@�G���ٿV��^��@[@�4@��� Ґ!?{����@�KaQ��ٿ���DN.�@��a�O 4@G�R�!?WIg?���@�KaQ��ٿ���DN.�@��a�O 4@G�R�!?WIg?���@�KaQ��ٿ���DN.�@��a�O 4@G�R�!?WIg?���@�KaQ��ٿ���DN.�@��a�O 4@G�R�!?WIg?���@P��N!�ٿ�]4�/�@��#��4@~���!?V�C��@P��N!�ٿ�]4�/�@��#��4@~���!?V�C��@P��N!�ٿ�]4�/�@��#��4@~���!?V�C��@5�^o�ٿ��A����@4ꄷ 4@n���!?��Xh�|�@C��l��ٿ�-U<8q�@��d��4@�Q��!?/�Z����@C��l��ٿ�-U<8q�@��d��4@�Q��!?/�Z����@C��l��ٿ�-U<8q�@��d��4@�Q��!?/�Z����@u��7�ٿ�o* �`�@�Ai5J 4@@��׮�!?B��1�.�@U?qA�ٿ*,o�:�@��7	�4@C�ٳ�!?�H.��z�@U?qA�ٿ*,o�:�@��7	�4@C�ٳ�!?�H.��z�@U?qA�ٿ*,o�:�@��7	�4@C�ٳ�!?�H.��z�@��~N)�ٿ�)n?��@�?�I�	4@��x��!?�k�C��@��~N)�ٿ�)n?��@�?�I�	4@��x��!?�k�C��@%	 ��ٿ�zP��4�@�e.if4@+�J�}�!?C��y/L�@%	 ��ٿ�zP��4�@�e.if4@+�J�}�!?C��y/L�@%	 ��ٿ�zP��4�@�e.if4@+�J�}�!?C��y/L�@�u�$]�ٿ�nѵ4�@U�D�4@Ks7䕐!?;l�;B3�@�u�$]�ٿ�nѵ4�@U�D�4@Ks7䕐!?;l�;B3�@�u�$]�ٿ�nѵ4�@U�D�4@Ks7䕐!?;l�;B3�@�u�$]�ٿ�nѵ4�@U�D�4@Ks7䕐!?;l�;B3�@��`7�ٿv^�F#D�@K���.
4@8�7D��!?���ɟk�@��`7�ٿv^�F#D�@K���.
4@8�7D��!?���ɟk�@��`7�ٿv^�F#D�@K���.
4@8�7D��!?���ɟk�@��`7�ٿv^�F#D�@K���.
4@8�7D��!?���ɟk�@��`7�ٿv^�F#D�@K���.
4@8�7D��!?���ɟk�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@%��ٿ7��mc��@���J4@�g�C��!?VptY�a�@!5��m�ٿwۯl��@����4@5)�r��!?;Hy�l�@!5��m�ٿwۯl��@����4@5)�r��!?;Hy�l�@!5��m�ٿwۯl��@����4@5)�r��!?;Hy�l�@Nj�qٿ�e�QY��@"�PD<4@��*�ѐ!?(V"gA�@�`�ٿ��Q0�@��Wm4@��4�!?އR�@�`�ٿ��Q0�@��Wm4@��4�!?އR�@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@���#�ٿ�fV�"��@��m4@���1ݐ!?w��9��@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@G��/�ٿT��^��@?h	�n4@���!?��L7���@�ч�W�ٿ�0�q*��@�斀4@
X�E��!?-k7�u�@�ч�W�ٿ�0�q*��@�斀4@
X�E��!?-k7�u�@m�mq��ٿ�Y�M{�@N�`ž4@���ǐ!?T��H��@z$�ۅ�ٿӁ�	Q�@����4@�z)Aݐ!?D��N.��@XC��ވٿ۳�����@�Vt�4@�/��!?���/��@�&��ٿ¦�O�U�@5�o�4@u˦k�!?͢���V�@�&��ٿ¦�O�U�@5�o�4@u˦k�!?͢���V�@�&��ٿ¦�O�U�@5�o�4@u˦k�!?͢���V�@�&��ٿ¦�O�U�@5�o�4@u˦k�!?͢���V�@�&��ٿ¦�O�U�@5�o�4@u˦k�!?͢���V�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@��j6ۉٿm��9��@�a�4@��z��!?q�`Cԧ�@f�J�Ɍٿ_��<�B�@2�>�4@�G"��!?�|�@f�J�Ɍٿ_��<�B�@2�>�4@�G"��!?�|�@��W�ٿf��\U�@@+Ȇ�4@�!R��!?s� ��@��W�ٿf��\U�@@+Ȇ�4@�!R��!?s� ��@F�ސЋٿ�*���4�@�ӽ�4@������!?�$����@F�ސЋٿ�*���4�@�ӽ�4@������!?�$����@�V�EE�ٿ���C}�@_�8�4@�mÐ!?���J��@ʞ�ٿ�9Ԓ���@�����4@���"�!?t3ɶ�@z\m�]�ٿw�Ƞ�@r�D��4@'��(�!?RWc�s�@z\m�]�ٿw�Ƞ�@r�D��4@'��(�!?RWc�s�@z\m�]�ٿw�Ƞ�@r�D��4@'��(�!?RWc�s�@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@/޵ (�ٿUi^��@���m�4@��}.�!?�bD"���@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@�Q�&�ٿ-��B��@� O�O4@s)��А!?�����@��VQa�ٿ�FT<���@r6W,[4@�����!?z9ݗ���@��JO��ٿ�C�ص��@o:Q��4@�6���!?��t���@��JO��ٿ�C�ص��@o:Q��4@�6���!?��t���@��JO��ٿ�C�ص��@o:Q��4@�6���!?��t���@��JO��ٿ�C�ص��@o:Q��4@�6���!?��t���@��JO��ٿ�C�ص��@o:Q��4@�6���!?��t���@ʏ��6}ٿ�̍���@El]�4@��B���!?���� �@ʏ��6}ٿ�̍���@El]�4@��B���!?���� �@��E|ٿb��<��@3�6�4@�$2�ڐ!?���X�@j�'�ٿ_� g�v�@�KZ��4@��	��!?��|�`�@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@�%�$��ٿ$��s��@�J�"%4@��c���!?\�S� ��@9Դ�a�ٿoEd8'��@X�ƀ4@�:���!?�4�s��@9Դ�a�ٿoEd8'��@X�ƀ4@�:���!?�4�s��@9Դ�a�ٿoEd8'��@X�ƀ4@�:���!?�4�s��@9Դ�a�ٿoEd8'��@X�ƀ4@�:���!?�4�s��@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�S�yڈٿ���!~�@��O�L4@������!?(�^�̳�@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@�n��Q�ٿ��'�[�@���T4@L�(���!?X�����@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@G n��ٿ���݃��@e��7X4@r���͐!?�:��Sx�@K����ٿ2+ՃW~�@�x��� 4@��Ꮠ!?�.ܝ%�@K����ٿ2+ՃW~�@�x��� 4@��Ꮠ!?�.ܝ%�@6�K�ٿ��U����@h�*ms4@^�	��!?4捇��@6�K�ٿ��U����@h�*ms4@^�	��!?4捇��@6�K�ٿ��U����@h�*ms4@^�	��!?4捇��@J���ٿUWb��^�@���74@r�`�s�!?]�ڽ>��@,�qg�ٿ $����@���4@wcM{�!?�m7����@,�qg�ٿ $����@���4@wcM{�!?�m7����@,�qg�ٿ $����@���4@wcM{�!?�m7����@
�MF�ٿ���o�@ ���4@�I��ؐ!?���q��@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@�$L�+�ٿ�N:F�@;�U`g4@Ly؞�!? 8�(�2�@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@oG�#�ٿ
��U��@��^�4@<���ې!?7Q!	N��@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@F�œ��ٿ�\G��@^3��4@�vH預!?��M�)�@�L7�	�ٿ��X�Z�@s����4@^Wֆ��!?m�tc��@�)<� �ٿ^ X0_��@���24@z����!?���v���@�)<� �ٿ^ X0_��@���24@z����!?���v���@�)<� �ٿ^ X0_��@���24@z����!?���v���@�)<� �ٿ^ X0_��@���24@z����!?���v���@�)<� �ٿ^ X0_��@���24@z����!?���v���@�)<� �ٿ^ X0_��@���24@z����!?���v���@"9�Ήٿϖt���@��z44@�+c0;�!?��E>���@"9�Ήٿϖt���@��z44@�+c0;�!?��E>���@"9�Ήٿϖt���@��z44@�+c0;�!?��E>���@"9�Ήٿϖt���@��z44@�+c0;�!?��E>���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@
���ٿ^u�A,��@�U��4@4�y�ې!?�{���@��ݠ��ٿ��U�X�@�˫�4@��>"�!?�IN8(��@��ݠ��ٿ��U�X�@�˫�4@��>"�!?�IN8(��@�G$VG�ٿC�{��"�@=QѝQ4@4B����!?����<z�@�G$VG�ٿC�{��"�@=QѝQ4@4B����!?����<z�@�G$VG�ٿC�{��"�@=QѝQ4@4B����!?����<z�@�G$VG�ٿC�{��"�@=QѝQ4@4B����!?����<z�@�3�/�ٿסIGP�@~�fG�4@��v$��!?4w�V7��@�3�/�ٿסIGP�@~�fG�4@��v$��!?4w�V7��@�3�/�ٿסIGP�@~�fG�4@��v$��!?4w�V7��@�3�/�ٿסIGP�@~�fG�4@��v$��!?4w�V7��@�3�/�ٿסIGP�@~�fG�4@��v$��!?4w�V7��@ƗWD@�ٿ�k�:��@+�T4@���Z��!?&l�7m3�@ƗWD@�ٿ�k�:��@+�T4@���Z��!?&l�7m3�@ƗWD@�ٿ�k�:��@+�T4@���Z��!?&l�7m3�@#ID���ٿ>���l��@��f�v4@��PR �!?�؏����@#ID���ٿ>���l��@��f�v4@��PR �!?�؏����@#ID���ٿ>���l��@��f�v4@��PR �!?�؏����@#ID���ٿ>���l��@��f�v4@��PR �!?�؏����@#ID���ٿ>���l��@��f�v4@��PR �!?�؏����@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@E6	��ٿ�]	i��@���[w4@���B�!?j
3m���@�ol~�ٿ [��8�@wN;�]4@/����!?�OPtj8�@�ol~�ٿ [��8�@wN;�]4@/����!?�OPtj8�@�ol~�ٿ [��8�@wN;�]4@/����!?�OPtj8�@�ə�a�ٿ��ۅ��@99�&*4@�Iܐ!?���L�"�@cDe�@�ٿ3]qٲ�@q=�Iy4@'#��!?��1�@�@l��ćٿ=����@ ^k4@��g���!?�t*�<��@m���5�ٿ�շ����@<��4@2D3���!?�b%%�@m���5�ٿ�շ����@<��4@2D3���!?�b%%�@m���5�ٿ�շ����@<��4@2D3���!?�b%%�@8��fp�ٿ�@'��*�@����Z4@�e����!?Gr��;�@8��fp�ٿ�@'��*�@����Z4@�e����!?Gr��;�@8��fp�ٿ�@'��*�@����Z4@�e����!?Gr��;�@8��fp�ٿ�@'��*�@����Z4@�e����!?Gr��;�@~��4�ٿ����ݺ�@��L^�4@�NTq�!?i&q���@~��4�ٿ����ݺ�@��L^�4@�NTq�!?i&q���@~��4�ٿ����ݺ�@��L^�4@�NTq�!?i&q���@�Xf~�|ٿݧQ�@���A4@�˲�!?$��`FK�@�%ʇٿȚB(^�@�E��4@�����!?�__�#�@�%ʇٿȚB(^�@�E��4@�����!?�__�#�@�%ʇٿȚB(^�@�E��4@�����!?�__�#�@�%ʇٿȚB(^�@�E��4@�����!?�__�#�@b7��͂ٿ�pi2k/�@?���?4@V�gŐ!?�
���-�@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�����ٿ���}=�@ݮ*�4@e�Nnِ!?]�\R��@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@�g��׊ٿ�ځ�m�@f�[/+4@tT��!?z� �V�@oU��Mٿn���B�@���4@�����!?��b���@oU��Mٿn���B�@���4@�����!?��b���@����.�ٿ,�N$�,�@8*+�{4@��0��!?e��˶��@����.�ٿ,�N$�,�@8*+�{4@��0��!?e��˶��@����.�ٿ,�N$�,�@8*+�{4@��0��!?e��˶��@����.�ٿ,�N$�,�@8*+�{4@��0��!?e��˶��@�s/��ٿ���(�@t>]y+4@w|=�ѐ!?�S>u��@�s/��ٿ���(�@t>]y+4@w|=�ѐ!?�S>u��@�s/��ٿ���(�@t>]y+4@w|=�ѐ!?�S>u��@�s/��ٿ���(�@t>]y+4@w|=�ѐ!?�S>u��@�l���ٿ���c��@���4@�
W�'�!?Γ����@�l���ٿ���c��@���4@�
W�'�!?Γ����@�|��(ٿX���e�@1����4@�J��!?��겼)�@�|��(ٿX���e�@1����4@�J��!?��겼)�@�|��(ٿX���e�@1����4@�J��!?��겼)�@�|��(ٿX���e�@1����4@�J��!?��겼)�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@_A�mV{ٿ���O�8�@�T�Wq4@i�un��!?驶�6{�@�ȍ��{ٿě9��@�<h�S4@}�-�!??��{��@7	�{��ٿ��wZ��@y,�!�4@�"���!?�6'fE�@7	�{��ٿ��wZ��@y,�!�4@�"���!?�6'fE�@7	�{��ٿ��wZ��@y,�!�4@�"���!?�6'fE�@7	�{��ٿ��wZ��@y,�!�4@�"���!?�6'fE�@7	�{��ٿ��wZ��@y,�!�4@�"���!?�6'fE�@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@H��#��ٿ/n0̵��@���:4@i��!? S��E��@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@ͮ�!S�ٿG
=*��@cE{�/4@\i͓ �!?w��5�f�@-��i�ٿ�7��m�@�+��q4@�g%@�!?] L4�T�@-��i�ٿ�7��m�@�+��q4@�g%@�!?] L4�T�@Tlrt��ٿI��,��@PX(��4@�ۉ�ڐ!?��</�X�@Tlrt��ٿI��,��@PX(��4@�ۉ�ڐ!?��</�X�@Tlrt��ٿI��,��@PX(��4@�ۉ�ڐ!?��</�X�@Tlrt��ٿI��,��@PX(��4@�ۉ�ڐ!?��</�X�@Tlrt��ٿI��,��@PX(��4@�ۉ�ڐ!?��</�X�@vHtO�ٿ�zdz^�@�b��N4@��I�!?W`��	��@vHtO�ٿ�zdz^�@�b��N4@��I�!?W`��	��@vHtO�ٿ�zdz^�@�b��N4@��I�!?W`��	��@'?��P�ٿH�V�$��@{8��<�3@�W6�!?�a����@'?��P�ٿH�V�$��@{8��<�3@�W6�!?�a����@'?��P�ٿH�V�$��@{8��<�3@�W6�!?�a����@�'�w~ٿ�"eo���@����.4@L;u��!?���i��@�'�w~ٿ�"eo���@����.4@L;u��!?���i��@@=��j�ٿ��n`%F�@+d��x4@*>��o�!?��&F���@@=��j�ٿ��n`%F�@+d��x4@*>��o�!?��&F���@�Ze(�ٿˉB)G��@���>4@�*pi�!?���\��@�Ze(�ٿˉB)G��@���>4@�*pi�!?���\��@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@���'d�ٿ;rs��@�����4@H�zVʐ!?>f��w�@��ν�{ٿ�2��&��@OP�4@�.���!?ָ�����@��ν�{ٿ�2��&��@OP�4@�.���!?ָ�����@�̤ٿ���	5��@��"�	4@�� ��!?X�ϰ+�@�̤ٿ���	5��@��"�	4@�� ��!?X�ϰ+�@�K,�ρٿ�p��m��@T+G�	4@t��O�!?v��#�=�@�K,�ρٿ�p��m��@T+G�	4@t��O�!?v��#�=�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@��(-V�ٿO����@Wr�4@�9=�{�!? X�Y�@�"�m��ٿ�����^�@;X�TI4@7�CG��!?�����P�@�"�m��ٿ�����^�@;X�TI4@7�CG��!?�����P�@�"�m��ٿ�����^�@;X�TI4@7�CG��!?�����P�@޽�1S�ٿ�We���@�� �4@hn(��!?�E�����@޽�1S�ٿ�We���@�� �4@hn(��!?�E�����@޽�1S�ٿ�We���@�� �4@hn(��!?�E�����@޽�1S�ٿ�We���@�� �4@hn(��!?�E�����@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@qAɅ�ٿ�Y�V��@'�"��4@����!?[�߬1k�@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@��c��ٿ�gB�T��@�``V�4@�R���!?]�ܧ��@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@7�.�Јٿ,xe(s��@Hm��4@�$�1�!?�3N�@��Gޅٿe��vC��@����%4@|�P�1�!?�`7%f��@�9S�ٿ���Cn�@�8�i�4@�g</�!?v|��)��@�9S�ٿ���Cn�@�8�i�4@�g</�!?v|��)��@�9S�ٿ���Cn�@�8�i�4@�g</�!?v|��)��@���-G�ٿ���\�@#*�U�4@��A�!?K�k®��@���-G�ٿ���\�@#*�U�4@��A�!?K�k®��@M��b}ٿ%	UK)�@(H�$�	4@�7���!?�h7��@M��b}ٿ%	UK)�@(H�$�	4@�7���!?�h7��@M��b}ٿ%	UK)�@(H�$�	4@�7���!?�h7��@M��b}ٿ%	UK)�@(H�$�	4@�7���!?�h7��@�y�b��ٿWT�''��@ A�cK
4@X>���!?�M����@�y�b��ٿWT�''��@ A�cK
4@X>���!?�M����@9RÀ�ٿM
Ba��@@_�`�	4@=,=���!?=m�)z�@9RÀ�ٿM
Ba��@@_�`�	4@=,=���!?=m�)z�@�3��ٿ�>�>�	�@�%>�|4@P�lߐ!?�p�-u{�@i4����ٿ�{���@��K@�	4@�Ǥ�!?���)gl�@i4����ٿ�{���@��K@�	4@�Ǥ�!?���)gl�@i4����ٿ�{���@��K@�	4@�Ǥ�!?���)gl�@i4����ٿ�{���@��K@�	4@�Ǥ�!?���)gl�@K��E�ٿ�y%"��@=���@4@�Nؐ!?�|��
��@K��E�ٿ�y%"��@=���@4@�Nؐ!?�|��
��@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@^C�K|ٿE;�m��@�{n4@��H��!?�n~�A<�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@��xh��ٿ�4�%��@E���4@@�+���!?5�#0�R�@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@�n}��ٿ�W�e��@_�-{4@���OԐ!?Z�H��@Ϛ��z�ٿ�}yU���@x���0 4@}tg���!?*��g�(�@Ϛ��z�ٿ�}yU���@x���0 4@}tg���!?*��g�(�@���̂ٿ	d(N�5�@K���� 4@r/��Ȑ!?��'�k�@���̂ٿ	d(N�5�@K���� 4@r/��Ȑ!?��'�k�@aU1��ٿwC�d���@j�&F4@��mC��!?�ܛؑ�@aU1��ٿwC�d���@j�&F4@��mC��!?�ܛؑ�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@i�ca{�ٿd�����@�1=e�4@Ec��!?���z]�@�]�%�~ٿ5q���@������3@��W�!?^9���@�]�%�~ٿ5q���@������3@��W�!?^9���@�]�%�~ٿ5q���@������3@��W�!?^9���@�]�%�~ٿ5q���@������3@��W�!?^9���@Z�\c�}ٿ����X��@H���z4@皂�Ɛ!?��)	G��@Z�\c�}ٿ����X��@H���z4@皂�Ɛ!?��)	G��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@/�Ɉٿ��A+Q�@����4@���tʐ!?m�"�"��@��t��ٿ���d���@p��c4@#�6G��!?�h�l��@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@�E��ٿ����f��@�'
4@��5���!?3Z����@���ga�ٿ"	}��@�]��4@C��ޤ�!?��%���@���ga�ٿ"	}��@�]��4@C��ޤ�!?��%���@���ga�ٿ"	}��@�]��4@C��ޤ�!?��%���@���ga�ٿ"	}��@�]��4@C��ޤ�!?��%���@���/��ٿ�ԵR��@H6�@M4@�M���!?��$���@j��'_�ٿ���O��@K��Hb4@5����!?����.u�@j��'_�ٿ���O��@K��Hb4@5����!?����.u�@j��'_�ٿ���O��@K��Hb4@5����!?����.u�@j��'_�ٿ���O��@K��Hb4@5����!?����.u�@j��'_�ٿ���O��@K��Hb4@5����!?����.u�@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@�����ٿ�Z����@Q(��4@yڀ��!?:6[�L��@&j3�;�ٿ�@�����@��Q�4@����ː!?�l���@&j3�;�ٿ�@�����@��Q�4@����ː!?�l���@&j3�;�ٿ�@�����@��Q�4@����ː!?�l���@3�;�L�ٿ�g����@U{e�4@�Q���!?/��Wq��@3�;�L�ٿ�g����@U{e�4@�Q���!?/��Wq��@3�;�L�ٿ�g����@U{e�4@�Q���!?/��Wq��@3�;�L�ٿ�g����@U{e�4@�Q���!?/��Wq��@"ظGۉٿ)4i h�@ǚS4@�5�ָ�!?�d���@"ظGۉٿ)4i h�@ǚS4@�5�ָ�!?�d���@"ظGۉٿ)4i h�@ǚS4@�5�ָ�!?�d���@"ظGۉٿ)4i h�@ǚS4@�5�ָ�!?�d���@�ɏg�ٿ���&�@�Sx��4@�ۻ
̐!?2���:��@C?��
�ٿfX�4��@A�����3@	]�͐!?�Z�c���@C?��
�ٿfX�4��@A�����3@	]�͐!?�Z�c���@�h���zٿd�����@ @N64@/��Ȑ!?;f����@p��ѿ�ٿ��� ��@��i� 4@V�]-֐!?QP�ƫ��@]"�+�ٿឿ���@	���4@3����!?����{�@]"�+�ٿឿ���@	���4@3����!?����{�@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@����O�ٿ���CtN�@�B�L� 4@8U��!?p�o���@J���(�ٿ��f�p�@H��L4@��a/ܐ!?���BZ"�@J���(�ٿ��f�p�@H��L4@��a/ܐ!?���BZ"�@/���|ٿ�S�o��@쯻Zn4@�4��!??����@/���|ٿ�S�o��@쯻Zn4@�4��!??����@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@ޟ9�p�ٿ�ҟgr��@z��ţ4@O�ʼ�!?L�U��@�U��!�ٿ�VҬF�@���4@;&�z�!?q�E���@W6�)�ٿ��
ZT��@8�i�4@B܃�!?&B#)	m�@W6�)�ٿ��
ZT��@8�i�4@B܃�!?&B#)	m�@W6�)�ٿ��
ZT��@8�i�4@B܃�!?&B#)	m�@W6�)�ٿ��
ZT��@8�i�4@B܃�!?&B#)	m�@['��ٿ鉺\��@�]L�4@��$���!?̹��\�@['��ٿ鉺\��@�]L�4@��$���!?̹��\�@['��ٿ鉺\��@�]L�4@��$���!?̹��\�@['��ٿ鉺\��@�]L�4@��$���!?̹��\�@['��ٿ鉺\��@�]L�4@��$���!?̹��\�@�s�~ٿ�G5L/��@|]&U�4@ϊH��!?c������@�s�~ٿ�G5L/��@|]&U�4@ϊH��!?c������@�s�~ٿ�G5L/��@|]&U�4@ϊH��!?c������@�s�~ٿ�G5L/��@|]&U�4@ϊH��!?c������@��I�ٿLO,t�@����4@V�c��!?ʹ�����@��I�ٿLO,t�@����4@V�c��!?ʹ�����@��I�ٿLO,t�@����4@V�c��!?ʹ�����@��I�ٿLO,t�@����4@V�c��!?ʹ�����@���R�ٿ%ޤ��@�L3P�4@�[�޽�!?���֩2�@���R�ٿ%ޤ��@�L3P�4@�[�޽�!?���֩2�@����@�ٿ��c�%q�@{EQk4@Wҡ���!?-��:K�@����@�ٿ��c�%q�@{EQk4@Wҡ���!?-��:K�@����@�ٿ��c�%q�@{EQk4@Wҡ���!?-��:K�@����@�ٿ��c�%q�@{EQk4@Wҡ���!?-��:K�@�2/��ٿ!Ý�\��@�"QKy4@�,����!?!R+�\:�@�2/��ٿ!Ý�\��@�"QKy4@�,����!?!R+�\:�@�2/��ٿ!Ý�\��@�"QKy4@�,����!?!R+�\:�@�2/��ٿ!Ý�\��@�"QKy4@�,����!?!R+�\:�@�$G���ٿ��3a�I�@S��4@1ۜwݐ!?T��V���@�[F��ٿ	l���@�����4@w����!?� [\��@%�ٿp�D8��@>.�04@y͇�!?jT�N�@%�ٿp�D8��@>.�04@y͇�!?jT�N�@�|����ٿ�W�N��@N�Ge4@%R���!?pD$ڋ��@�|����ٿ�W�N��@N�Ge4@%R���!?pD$ڋ��@�|����ٿ�W�N��@N�Ge4@%R���!?pD$ڋ��@�|����ٿ�W�N��@N�Ge4@%R���!?pD$ڋ��@�|����ٿ�W�N��@N�Ge4@%R���!?pD$ڋ��@����ٿ�n�4��@�2*��4@dI�<��!?n�_yY��@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@�DS7�ٿ��K/N�@���K�4@9̬0}�!?P�����@T�NKЌٿ�V{`���@��/)�4@����:�!?�WDle��@T�NKЌٿ�V{`���@��/)�4@����:�!?�WDle��@T�NKЌٿ�V{`���@��/)�4@����:�!?�WDle��@T�NKЌٿ�V{`���@��/)�4@����:�!?�WDle��@T�NKЌٿ�V{`���@��/)�4@����:�!?�WDle��@�����ٿ��;fq�@��!��4@>�}m:�!?�yd�q�@��-`�ٿ���.��@���4@�;���!?.+�_[�@��-`�ٿ���.��@���4@�;���!?.+�_[�@��-`�ٿ���.��@���4@�;���!?.+�_[�@��-`�ٿ���.��@���4@�;���!?.+�_[�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@�rݵ�ٿ]e�h#�@H�l04@�����!?�e��qy�@iATn��ٿ��">�@����3@��Lt��!?����I�@iATn��ٿ��">�@����3@��Lt��!?����I�@iATn��ٿ��">�@����3@��Lt��!?����I�@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@�=�q �ٿ�{�(�@�]Ku4@N<$,d�!?�rf����@��a#3�ٿ�wt����@���]c4@���Z�!?��r� ��@<�+�
�ٿg�CB��@����m4@��yې!?��I%�@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@����ٿ���K�@Q�^�4@�(�b!?�L�!��@Z�0B�ٿ�Dn�@9���h4@C�z��!?v��Q��@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@Y|�H�ٿ!C����@��R�4@���ͣ�!??����@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@
��bb�ٿ��X���@5��}�4@G���l�!?�Õp���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@���Ǉٿ09z�57�@'\M�"4@��S��!?��s���@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@��pU�ٿ��9���@SNS�/4@q�����!?7��� �@�ۇ��ٿ2�_q�.�@z��|��3@+�U��!?v�u �j�@�ۇ��ٿ2�_q�.�@z��|��3@+�U��!?v�u �j�@�ۇ��ٿ2�_q�.�@z��|��3@+�U��!?v�u �j�@�ۇ��ٿ2�_q�.�@z��|��3@+�U��!?v�u �j�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@��Dt,�ٿ�f,E��@HN	&4@D��
��!?��~�<J�@���q�ٿD�5n1��@�S�� 4@1�����!?��;�a��@�&�\8�ٿ���&��@��s4@w�{"z�!?���2��@�&�\8�ٿ���&��@��s4@w�{"z�!?���2��@�&�\8�ٿ���&��@��s4@w�{"z�!?���2��@�>Wb!�ٿ �����@誾�{4@������!?	� ����@�-řٿ��ȃ�E�@''�Z54@���T��!?P"���@�-řٿ��ȃ�E�@''�Z54@���T��!?P"���@�-řٿ��ȃ�E�@''�Z54@���T��!?P"���@�-řٿ��ȃ�E�@''�Z54@���T��!?P"���@���L�ٿ�J䬝��@sqo}�4@(��e��!?�%�$��@�;�G��ٿ��~���@D`ߋ&4@Obhܐ!?��o����@�;�G��ٿ��~���@D`ߋ&4@Obhܐ!?��o����@�;�G��ٿ��~���@D`ߋ&4@Obhܐ!?��o����@�;�G��ٿ��~���@D`ߋ&4@Obhܐ!?��o����@�;�G��ٿ��~���@D`ߋ&4@Obhܐ!?��o����@Οlc�ٿ���q���@KMIu&4@�Ӧ+א!?_L�]��@Οlc�ٿ���q���@KMIu&4@�Ӧ+א!?_L�]��@Οlc�ٿ���q���@KMIu&4@�Ӧ+א!?_L�]��@IS5FZ�ٿ]L&js�@"ʙJ4@��?���!?]?�:���@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��"r��ٿ�F�� ��@��`T�4@ɬ6��!?�ڋ}�@��n��ٿO�w���@�\�"g4@���T��!?}��P��@D:V��ٿ�¼�-�@4�w�4@��k�!?h�����@D:V��ٿ�¼�-�@4�w�4@��k�!?h�����@D:V��ٿ�¼�-�@4�w�4@��k�!?h�����@D:V��ٿ�¼�-�@4�w�4@��k�!?h�����@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@[���ٿ���)Q�@��~�[4@{^���!?�C胀G�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�/Âٿ�vFF���@��N4@0����!?]���8�@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@�ؒ߁ٿ�����@����4@4�A:�!?�),c9��@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@1-���ٿ��]�e��@����c4@�G�Ŀ�!?͂e���@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@w&�9#�ٿZU�a��@�{�{4@��ǐ!?0�u^��@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@]W-.h�ٿ���$���@o�=�x4@� Ӫ��!?#*���&�@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@�!Vr�ٿos&lH��@D�5�4@�+�S��!?|WGN��@��܄J}ٿd�c� ��@���T�4@a�^�֐!?��Ol9�@��܄J}ٿd�c� ��@���T�4@a�^�֐!?��Ol9�@��܄J}ٿd�c� ��@���T�4@a�^�֐!?��Ol9�@*�bs?�ٿ_�W�@B_}�34@�P�!?��FH/
�@*�bs?�ٿ_�W�@B_}�34@�P�!?��FH/
�@*�bs?�ٿ_�W�@B_}�34@�P�!?��FH/
�@*�bs?�ٿ_�W�@B_}�34@�P�!?��FH/
�@*�bs?�ٿ_�W�@B_}�34@�P�!?��FH/
�@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@Su��[}ٿ�����@��{J4@w�vPʐ!?0&�4��@:����~ٿ����@���4@�^R���!?J?����@:����~ٿ����@���4@�^R���!?J?����@��B��ٿ��Y���@gpx$+4@��dL�!?�a���@��B��ٿ��Y���@gpx$+4@��dL�!?�a���@��B��ٿ��Y���@gpx$+4@��dL�!?�a���@��B��ٿ��Y���@gpx$+4@��dL�!?�a���@l���t�ٿ������@A+Yr�	4@���ސ!?��+,D9�@l���t�ٿ������@A+Yr�	4@���ސ!?��+,D9�@��7uA�ٿWU�U&��@H��/4@	 	�!?����@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@�D��ٿu�y����@��^�<4@�*d��!?`}�Ɉ��@����ٿY�S[��@��; �4@�Zb\z�!?�r�`��@����ٿY�S[��@��; �4@�Zb\z�!?�r�`��@@����ٿ�~f-�q�@i�<&4@�mf��!?�5����@@����ٿ�~f-�q�@i�<&4@�mf��!?�5����@V1���ٿ+^�\�	�@�<_�4@�i8A��!?R>F���@1�� �ٿ:k�2�#�@+lް4@r��<�!?1]��!�@1�� �ٿ:k�2�#�@+lް4@r��<�!?1]��!�@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@A�y���ٿ�rK]-��@�
LS4@^<U�Ð!?7�92���@X�7��ٿjr[�*�@�>�
4@ �\��!?	��8��@?@��ٿ�� p/�@ ���-4@�c\~�!?YБ�Mu�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@���x	�ٿk��^Z��@�����4@�Q�c��!?��F�C%�@����ٿ�|�m��@�w:�4@݁��!?����@����ٿ�|�m��@�w:�4@݁��!?����@����ٿ�|�m��@�w:�4@݁��!?����@(�6�ٿ� ύ�]�@����q4@���
�!?�sD�m`�@(�6�ٿ� ύ�]�@����q4@���
�!?�sD�m`�@(�6�ٿ� ύ�]�@����q4@���
�!?�sD�m`�@(�6�ٿ� ύ�]�@����q4@���
�!?�sD�m`�@(�6�ٿ� ύ�]�@����q4@���
�!?�sD�m`�@���<�ٿH�D��@�u�4@i<1sw�!?��,���@���yٿ��/�I��@k�R84@���s�!?r�+���@��~��~ٿ�}$��@8�#�C4@���T9�!?8����@�wB/��ٿ�Ċn�@zvaLz4@��J�!?7�\����@ER.$�ٿ�#���@�/U١4@���a�!?+�� e�@ER.$�ٿ�#���@�/U١4@���a�!?+�� e�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@�A��
�ٿg�0��@��bݓ4@�GkG��!?���:A�@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@*��!z�ٿ(�S����@���L4@ǫiĐ!?��~��@�� ��ٿþ�˼�@��x��4@���D�!?ud��@�� ��ٿþ�˼�@��x��4@���D�!?ud��@�l���ٿ��fj-�@��?��4@��@��!?�L`��@�l���ٿ��fj-�@��?��4@��@��!?�L`��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�����ٿ&!Cu�P�@4v��.4@	�p��!?�ߧ�3��@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@�1�A�ٿ* �:C�@��t�<4@8/�q��!?�l.qAO�@��p�ٿ�8i�@�BFq�4@ث����!?���d?��@n-ҤN�ٿm�(�@B�2�4@�����!?�"���@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@�%|(��ٿ1�� �@h�x6F4@(g�ǐ�!?eVנ �@!�ٿrc�e���@���Q�4@!�𻪐!?6�^hcu�@!�ٿrc�e���@���Q�4@!�𻪐!?6�^hcu�@!�ٿrc�e���@���Q�4@!�𻪐!?6�^hcu�@/>5��ٿ'Dx�MO�@ݐ�4@'�m���!?±���@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@6<4H�ٿ��Æ�_�@�ߤ��4@*K�ݐ!?�5F߯��@ ���,�ٿ�����9�@��aW4@M�W��!?���O�G�@ ���,�ٿ�����9�@��aW4@M�W��!?���O�G�@���y�ٿ�����O�@�MmT�4@kuBi(�!?��r�@} ˪�ٿ~�Ci��@�����4@����7�!?�bR`0q�@>'��ٿ;9��*��@��4@22��!?�%A��@�^���{ٿ0�l���@���X 4@)H�cƐ!?*���H�@�^���{ٿ0�l���@���X 4@)H�cƐ!?*���H�@�����ٿ��8��@b��ې�3@��֩�!?#[v��@p|��ٿ�Õ]���@��ǌ4@9�$��!?5��wz�@T�����ٿ�^d���@�S�g4@j��X��!?����C�@T�����ٿ�^d���@�S�g4@j��X��!?����C�@T�����ٿ�^d���@�S�g4@j��X��!?����C�@T�����ٿ�^d���@�S�g4@j��X��!?����C�@���,ˆٿ4��g�@UH,@>4@U���!?
dK�w��@���,ˆٿ4��g�@UH,@>4@U���!?
dK�w��@���,ˆٿ4��g�@UH,@>4@U���!?
dK�w��@��>FɄٿ�D�UW�@ �{T�3@�'��!?�F�@��W�T�ٿV�+��@�*�PR4@�s���!?��W~p�@A�����ٿ�p����@���sS4@�$��!?W�"YH�@���m�~ٿ������@�#��S4@e��2�!?7ĵ�і�@���m�~ٿ������@�#��S4@e��2�!?7ĵ�і�@bnx�w|ٿ�֌ҩ�@�4Km 4@���V�!?.�C���@bnx�w|ٿ�֌ҩ�@�4Km 4@���V�!?.�C���@bnx�w|ٿ�֌ҩ�@�4Km 4@���V�!?.�C���@z+�ޫ�ٿ���5��@7j�0�4@�;��5�!?�m�j��@z+�ޫ�ٿ���5��@7j�0�4@�;��5�!?�m�j��@z+�ޫ�ٿ���5��@7j�0�4@�;��5�!?�m�j��@P����ٿv|C�9�@w.�x}4@�]Z���!?[V +���@���"�~ٿ���Y���@1��y5 4@W�<�Ґ!?�K!���@���"�~ٿ���Y���@1��y5 4@W�<�Ґ!?�K!���@���L~ٿ-�S�	�@ӀТ 4@Dv�X��!?ljf	���@�VT܎{ٿg�����@z#+���3@��9j�!?Q�+*V7�@*��Q�ٿr������@^�_Z4@+U�)�!?���~G��@*��Q�ٿr������@^�_Z4@+U�)�!?���~G��@*��Q�ٿr������@^�_Z4@+U�)�!?���~G��@*��Q�ٿr������@^�_Z4@+U�)�!?���~G��@*��Q�ٿr������@^�_Z4@+U�)�!?���~G��@hڸ@��ٿ��4=��@2�V94@�F�(9�!?�D-o�@hڸ@��ٿ��4=��@2�V94@�F�(9�!?�D-o�@hڸ@��ٿ��4=��@2�V94@�F�(9�!?�D-o�@hڸ@��ٿ��4=��@2�V94@�F�(9�!?�D-o�@hڸ@��ٿ��4=��@2�V94@�F�(9�!?�D-o�@	 Ki"�ٿQǆ$�'�@��v4@H��=�!?y�%���@	 Ki"�ٿQǆ$�'�@��v4@H��=�!?y�%���@	 Ki"�ٿQǆ$�'�@��v4@H��=�!?y�%���@	 Ki"�ٿQǆ$�'�@��v4@H��=�!?y�%���@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@�,Z�̊ٿT ��%��@���X�4@�:����!?���fR�@|�	�ٿ�(Z���@=�o�4@��@�!?O�@"|��@|�	�ٿ�(Z���@=�o�4@��@�!?O�@"|��@|�	�ٿ�(Z���@=�o�4@��@�!?O�@"|��@|�	�ٿ�(Z���@=�o�4@��@�!?O�@"|��@�uQ��ٿ;�zH�@<n-��4@�.a_Ր!?%A��t�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@�Id7<�ٿEb����@̌V��4@ �uv��!??���{0�@��~�ٿ��1�@����4@n.&��!?&��"�~�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@Ѕ+���ٿQ�����@LV 	�4@f{�䤐!?k�D�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@м
�ٿ��v��*�@�W��U4@G����!?�4���z�@R.ǐ��ٿ�m�R���@�d��� 4@.?���!?�IE�i��@��Z�ٿ�*-�8�@��=4@k�E��!?SvFs��@��Z�ٿ�*-�8�@��=4@k�E��!?SvFs��@��Z�ٿ�*-�8�@��=4@k�E��!?SvFs��@��Z�ٿ�*-�8�@��=4@k�E��!?SvFs��@��Z�ٿ�*-�8�@��=4@k�E��!?SvFs��@��[^F~ٿN��_�@P�w4@*����!?N]�#��@��[^F~ٿN��_�@P�w4@*����!?N]�#��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@&�ӁٿL��?��@�7�d4@.dt���!?��ς��@�,��|ٿ1���C��@�-.�	4@E�ݯ�!?[��ft��@�,��|ٿ1���C��@�-.�	4@E�ݯ�!?[��ft��@V�_ӷ�ٿ��>��v�@Wbt9 4@&b-��!?�Y����@V�_ӷ�ٿ��>��v�@Wbt9 4@&b-��!?�Y����@)Ex�ٿ��e�#��@�Zq}� 4@͚"�!�!?>����@��Uz	�ٿ"����@%�Ip� 4@�!z��!?��g��G�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@ Q0܉ٿ�ut�@��r9� 4@!VU�C�!?-��%U�@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@�Gb���ٿd��/G�@�dK��4@1Z��ϐ!?�_#��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@o�g��ٿ�٭r��@?�]v�4@����!?�"JC��@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@��,�ٿ�&���@����4@�%<Ԑ!?��{��7�@�k�(�ٿE��{�@���:4@h��㷐!?|�[�b�@�k�(�ٿE��{�@���:4@h��㷐!?|�[�b�@�k�(�ٿE��{�@���:4@h��㷐!?|�[�b�@�k�(�ٿE��{�@���:4@h��㷐!?|�[�b�@is��wٿ\�u�~�@b�>�4@������!?�;�/�@is��wٿ\�u�~�@b�>�4@������!?�;�/�@is��wٿ\�u�~�@b�>�4@������!?�;�/�@is��wٿ\�u�~�@b�>�4@������!?�;�/�@t���ٿP��~���@q�o�;4@(�%�0�!?�X��p�@z`�^�ٿ�^ a?D�@{;C�;4@^��h�!?��N��@z`�^�ٿ�^ a?D�@{;C�;4@^��h�!?��N��@"1�"j�ٿ�W�{q��@�o�94@�$Â��!?��k�(��@"1�"j�ٿ�W�{q��@�o�94@�$Â��!?��k�(��@"1�"j�ٿ�W�{q��@�o�94@�$Â��!?��k�(��@"1�"j�ٿ�W�{q��@�o�94@�$Â��!?��k�(��@�u_�Z�ٿ�HU���@o��\4@p�_���!?Ee�͜�@�u_�Z�ٿ�HU���@o��\4@p�_���!?Ee�͜�@�u_�Z�ٿ�HU���@o��\4@p�_���!?Ee�͜�@�u_�Z�ٿ�HU���@o��\4@p�_���!?Ee�͜�@�u_�Z�ٿ�HU���@o��\4@p�_���!?Ee�͜�@,�R]�ٿ�Z����@'�fQ4@L���ސ!?�%�Ξ�@�2�[E�ٿ�3�r���@�[Q� 4@�L6&@�!?�縑���@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@���˸ٿ<��7��@�WVׅ4@���Ő!?JQ"諃�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@��ˀ��ٿR������@��Z4@��E��!?�>.�++�@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@�?uv�ٿJ��`k��@�5?4@y�J��!?C�x��@J5&�҃ٿO���2��@D�=-�4@R����!?��a���@��q��ٿ�u�h�@��Ҋ�4@u�SY��!?�TG��@��q��ٿ�u�h�@��Ҋ�4@u�SY��!?�TG��@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@�cc]�ٿ�g���@�Q ��4@��Y��!?�~G���@{�7!��ٿ���4��@��O��4@���̐!?1Za���@{�7!��ٿ���4��@��O��4@���̐!?1Za���@��ԍٿ8k���@h�I�Q4@��6���!?�X"����@/~�&�ٿn����@���=<4@�����!?ˠ%�h��@��@$�ٿ�E��Qa�@W��}�4@��z�א!?ގ�5��@��@$�ٿ�E��Qa�@W��}�4@��z�א!?ގ�5��@��@$�ٿ�E��Qa�@W��}�4@��z�א!?ގ�5��@7�<v�ٿ��{'��@��ʫo4@$<>��!?���py��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@tc�,˂ٿt�n��`�@qǡ�X4@Gg���!?�A_c��@P�;�&�ٿu������@)�%4@)�5���!?�'����@P�;�&�ٿu������@)�%4@)�5���!?�'����@�Vv�m�ٿ�N�R�@��4@+��ɐ!?+j���@�Vv�m�ٿ�N�R�@��4@+��ɐ!?+j���@�Vv�m�ٿ�N�R�@��4@+��ɐ!?+j���@�Vv�m�ٿ�N�R�@��4@+��ɐ!?+j���@/�o2�ٿlp#����@�`���4@Õ_��!?7Z2�F��@/�o2�ٿlp#����@�`���4@Õ_��!?7Z2�F��@/�o2�ٿlp#����@�`���4@Õ_��!?7Z2�F��@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@,:y��ٿ
�D���@V���4@WT���!?�X����@h��pهٿ�3b��@E�b64@X�':�!?x7����@h��pهٿ�3b��@E�b64@X�':�!?x7����@h��pهٿ�3b��@E�b64@X�':�!?x7����@�"u�G�ٿ��˗&�@�ة4@C�g��!?I�r�O�@�"u�G�ٿ��˗&�@�ة4@C�g��!?I�r�O�@�"u�G�ٿ��˗&�@�ة4@C�g��!?I�r�O�@�I��8�ٿ�\�c>�@g���4@W���!?Ho�*v��@�I��8�ٿ�\�c>�@g���4@W���!?Ho�*v��@�I��8�ٿ�\�c>�@g���4@W���!?Ho�*v��@�I��8�ٿ�\�c>�@g���4@W���!?Ho�*v��@��`�a�ٿe���(�@"ۡbJ4@�,����!?�[�u���@��`�a�ٿe���(�@"ۡbJ4@�,����!?�[�u���@��`�a�ٿe���(�@"ۡbJ4@�,����!?�[�u���@��`�a�ٿe���(�@"ۡbJ4@�,����!?�[�u���@��`�a�ٿe���(�@"ۡbJ4@�,����!?�[�u���@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�2*,Q�ٿz`1?�@���Y�4@�3t��!?�]��8S�@�08N�ٿ�.�g�@��hJ�4@ 	hTŐ!?��8��@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@x��,�ٿ��%�4�@lA��4@��`o�!?`�C\�@�}7���ٿ��/:ͧ�@�kw�N4@K��9ߐ!?��@��@,���ٿ�%�����@���%4@�n���!?8d�

{�@,���ٿ�%�����@���%4@�n���!?8d�

{�@|S����ٿ4�g����@�rk�4@ȴg|��!?nv�V�@|S����ٿ4�g����@�rk�4@ȴg|��!?nv�V�@&��P��ٿ��!�6x�@nl��k4@���3��!?�,1���@&��P��ٿ��!�6x�@nl��k4@���3��!?�,1���@&��P��ٿ��!�6x�@nl��k4@���3��!?�,1���@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@�#X��ٿC��$H�@e ���4@%�JH!?�S�6��@_`;�˂ٿg>�Ȯ��@(&��4@XR_��!?l�6@O�@_`;�˂ٿg>�Ȯ��@(&��4@XR_��!?l�6@O�@_`;�˂ٿg>�Ȯ��@(&��4@XR_��!?l�6@O�@_`;�˂ٿg>�Ȯ��@(&��4@XR_��!?l�6@O�@_`;�˂ٿg>�Ȯ��@(&��4@XR_��!?l�6@O�@c�]Hm�ٿ��@��#�@�4�G4@H"�l̐!?��񇠈�@c�]Hm�ٿ��@��#�@�4�G4@H"�l̐!?��񇠈�@c�]Hm�ٿ��@��#�@�4�G4@H"�l̐!?��񇠈�@�g�Fވٿ��i��@�����4@(#��ؐ!?ʧI����@�g�Fވٿ��i��@�����4@(#��ؐ!?ʧI����@�g�Fވٿ��i��@�����4@(#��ؐ!?ʧI����@�KA���ٿ���>�@^A77\4@�t �ɐ!?�C�g��@�='[ƈٿ,��Mn9�@�ҥ�4@�;jÐ!?��چ�@�ӥ1�ٿ���'��@^u)~�4@ka�ǐ!?%o���@�ӥ1�ٿ���'��@^u)~�4@ka�ǐ!?%o���@�}��ٿ3�$I�@�\y8�4@=�|?��!?G���լ�@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@f�]���ٿȅ�>0�@��r34@���;x�!?����u��@+p��#�ٿQ!���@��̱}4@��գ�!?��SP��@�J��݉ٿL>g"ǥ�@��I}�4@��p՗�!?<[�L���@�J��݉ٿL>g"ǥ�@��I}�4@��p՗�!?<[�L���@�CD�ٿ��W`��@�W���4@������!?�F����@��1�9�ٿ������@h&��4@)�JQŐ!?���Jk��@��1�9�ٿ������@h&��4@)�JQŐ!?���Jk��@%"-�ٿ#S�x�N�@�y��4@6�[�!?'0�\S��@�^�
��ٿ�T)����@����4@v]%/+�!?�X��E�@�^�
��ٿ�T)����@����4@v]%/+�!?�X��E�@�^�
��ٿ�T)����@����4@v]%/+�!?�X��E�@�^�
��ٿ�T)����@����4@v]%/+�!?�X��E�@��&Azٿbt~7�@�w�b�4@1���ڐ!?<%V)� �@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@}��}ٿLeU���@Gh�~4@���ΐ!?�����@�D�,�}ٿ�=%7���@?VOa.4@p`^b�!?��O:���@;8�:�ٿW�0s֋�@�)~��4@ ի!Ґ!?!M�<� �@;8�:�ٿW�0s֋�@�)~��4@ ի!Ґ!?!M�<� �@;8�:�ٿW�0s֋�@�)~��4@ ի!Ґ!?!M�<� �@q4�0�ٿ��u�U�@�̧Z�4@k��uݐ!?�K.g�@q4�0�ٿ��u�U�@�̧Z�4@k��uݐ!?�K.g�@q4�0�ٿ��u�U�@�̧Z�4@k��uݐ!?�K.g�@�8t$L�ٿ�l�UU�@��h�4@�b��!?r����@�8t$L�ٿ�l�UU�@��h�4@�b��!?r����@�8t$L�ٿ�l�UU�@��h�4@�b��!?r����@�8t$L�ٿ�l�UU�@��h�4@�b��!?r����@����ٿ?o�\b+�@U�]�4@}�8Gؐ!?�H}>��@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@=��[��ٿ��f�B��@�0�Y4@�1t=�!?����#�@��tٿP��\���@�wF��4@a�;�!?��֒��@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@4��9��ٿ���9t�@Lrďw4@7�)��!?һ��L�@�P:՟�ٿ�K� ;�@43��Z4@O=ٞ��!?���e��@�P:՟�ٿ�K� ;�@43��Z4@O=ٞ��!?���e��@�P:՟�ٿ�K� ;�@43��Z4@O=ٞ��!?���e��@�P:՟�ٿ�K� ;�@43��Z4@O=ٞ��!?���e��@�P:՟�ٿ�K� ;�@43��Z4@O=ٞ��!?���e��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@C�G��ٿ�d,>r��@' ��4@���I��!?m�u��@xS����ٿ+,pC� �@�t�;4@���g��!?(3oe��@xS����ٿ+,pC� �@�t�;4@���g��!?(3oe��@xS����ٿ+,pC� �@�t�;4@���g��!?(3oe��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@�>�
݆ٿ��ӫȇ�@e�Ӡ�4@A�Ў�!?K�<��@f�jN�ٿ�O�A�F�@�n���4@�-���!?|�~�L�@f�jN�ٿ�O�A�F�@�n���4@�-���!?|�~�L�@f�jN�ٿ�O�A�F�@�n���4@�-���!?|�~�L�@f�jN�ٿ�O�A�F�@�n���4@�-���!?|�~�L�@f�jN�ٿ�O�A�F�@�n���4@�-���!?|�~�L�@-Tx!�ٿ�~+�2�@�*��4@�Ǉ���!?/r,]g�@-Tx!�ٿ�~+�2�@�*��4@�Ǉ���!?/r,]g�@-Tx!�ٿ�~+�2�@�*��4@�Ǉ���!?/r,]g�@�=�i�ٿ�n�D2O�@p�P�4@��}Ȑ!?��(B��@�=�i�ٿ�n�D2O�@p�P�4@��}Ȑ!?��(B��@������ٿ3�g�"��@�+<w4@Y��k�!?��{���@������ٿ3�g�"��@�+<w4@Y��k�!?��{���@������ٿ3�g�"��@�+<w4@Y��k�!?��{���@������ٿ3�g�"��@�+<w4@Y��k�!?��{���@������ٿ3�g�"��@�+<w4@Y��k�!?��{���@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@��ʄٿ��jm���@;�@��4@"�O��!?�j%�6^�@v��R�ٿ�\���@s���54@����!?L��n�@v��R�ٿ�\���@s���54@����!?L��n�@v��R�ٿ�\���@s���54@����!?L��n�@v��R�ٿ�\���@s���54@����!?L��n�@v��R�ٿ�\���@s���54@����!?L��n�@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@d�(�Êٿ%s:5��@˝�;_4@U�G��!?�@)��@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@�Ȉ�!�ٿ�e���@�/v�4@$�ǘ��!?T��� �@G�L���ٿ)�^�T��@�&)�4@����Ґ!?�r��@6�@G�L���ٿ)�^�T��@�&)�4@����Ґ!?�r��@6�@G�L���ٿ)�^�T��@�&)�4@����Ґ!?�r��@6�@G�L���ٿ)�^�T��@�&)�4@����Ґ!?�r��@6�@����҆ٿ�u'��@�z�x4@9�1��!?��S�t��@����҆ٿ�u'��@�z�x4@9�1��!?��S�t��@����҆ٿ�u'��@�z�x4@9�1��!?��S�t��@�M�l�ٿ�[����@�X��A4@4PG���!?�Y���@II�͋ٿ���HrY�@��/�[4@rU�Q��!?�a�؝��@�h*�ٿ�	�,�@�Db��4@H ��g�!?�VR[��@���ٿ$^��,L�@���:4@����!?R�z�K��@���ٿ$^��,L�@���:4@����!?R�z�K��@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@t�����ٿ��Nԧq�@'ɽ`�4@rG5jѐ!?��8��X�@VJ^N��ٿϾ��g�@�7>4@]�si�!?r�.��@kA�-�ٿ
�,E��@�=R�4@8�㚒�!?pE�`w�@kA�-�ٿ
�,E��@�=R�4@8�㚒�!?pE�`w�@kA�-�ٿ
�,E��@�=R�4@8�㚒�!?pE�`w�@��h��ٿ��K��@�N�^4@�K_k��!?�����@鵩��ٿ�l.�i�@���"4@ �"?��!?�pP/�k�@鵩��ٿ�l.�i�@���"4@ �"?��!?�pP/�k�@�_=c��ٿ]�y�R�@D��>�4@S�Ѧ�!?h.�7F��@�_=c��ٿ]�y�R�@D��>�4@S�Ѧ�!?h.�7F��@��Ջ��ٿp�o��7�@O�*�e4@�_P���!?�5p��@��Ջ��ٿp�o��7�@O�*�e4@�_P���!?�5p��@��H���ٿ:�%�A�@�ba
4@�����!?ҡN��@��H���ٿ:�%�A�@�ba
4@�����!?ҡN��@W`z�}�ٿ��.A��@��0��4@�Z��ɐ!?��s��^�@W`z�}�ٿ��.A��@��0��4@�Z��ɐ!?��s��^�@W`z�}�ٿ��.A��@��0��4@�Z��ɐ!?��s��^�@��]<�ٿT�I�F5�@�ߥ�4@��͐!?�c���@��]<�ٿT�I�F5�@�ߥ�4@��͐!?�c���@zҸ�T�ٿ���~�@�8�� 4@ �\��!?��n�l�@�c��ٿ�p��@�;fF4@����r�!?�W�&��@�c��ٿ�p��@�;fF4@����r�!?�W�&��@�c��ٿ�p��@�;fF4@����r�!?�W�&��@߭�ՄٿwM%WB�@�D�� 4@���#E�!?����B�@߭�ՄٿwM%WB�@�D�� 4@���#E�!?����B�@��!�:�ٿ	���l�@���64@��*4�!?PL��� �@��B�ٿ���s�@2��:\4@q�6\�!?trd%@�@��B�ٿ���s�@2��:\4@q�6\�!?trd%@�@��B�ٿ���s�@2��:\4@q�6\�!?trd%@�@��B�ٿ���s�@2��:\4@q�6\�!?trd%@�@��B�ٿ���s�@2��:\4@q�6\�!?trd%@�@�dt��ٿ�S��_`�@r29b4@y2
R��!?U��>���@�dt��ٿ�S��_`�@r29b4@y2
R��!?U��>���@�dt��ٿ�S��_`�@r29b4@y2
R��!?U��>���@>1�P��ٿ�l��T�@���"4@[�`�!?�UU;���@a�y�y�ٿ�V��f��@0�-�4@���ʐ!?T�v�e��@��$7*�ٿ9��]���@���y4@�k���!?h~�
��@3����ٿ�B�K��@���$�4@�߇ѐ!?�6��|�@3����ٿ�B�K��@���$�4@�߇ѐ!?�6��|�@z�iʊٿ��\:��@!B-�4@�~���!?O�%�5y�@z�iʊٿ��\:��@!B-�4@�~���!?O�%�5y�@?�yF:�ٿ8����/�@(sA�4@MWf��!?!TG��@?�yF:�ٿ8����/�@(sA�4@MWf��!?!TG��@��S�؋ٿtV����@;��+4@*:�ǐ!?K{��)��@��S�؋ٿtV����@;��+4@*:�ǐ!?K{��)��@$[��ٿ���{��@�P�.4@����!?G<�3�y�@$[��ٿ���{��@�P�.4@����!?G<�3�y�@$[��ٿ���{��@�P�.4@����!?G<�3�y�@$[��ٿ���{��@�P�.4@����!?G<�3�y�@���N��ٿQ�z��y�@f��.4@;��8��!?�f��+�@���N��ٿQ�z��y�@f��.4@;��8��!?�f��+�@���N��ٿQ�z��y�@f��.4@;��8��!?�f��+�@���N��ٿQ�z��y�@f��.4@;��8��!?�f��+�@���N��ٿQ�z��y�@f��.4@;��8��!?�f��+�@y�̜h�ٿw��ŧ�@:W��,	4@�:��Ð!?
��Z��@<�,���ٿ���W�@�β�!4@�]�ʐ!?���@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@�ub���ٿ=�y����@�r,�4@gY��ܐ!?\�c�	��@P0��ٿ#%k H�@(�n�D4@~��!?�
n�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@���q��ٿ�����@��4@�����!?@j�g]�@}]��r�ٿ��T�3\�@�q4@讏�
�!?�W<��F�@}]��r�ٿ��T�3\�@�q4@讏�
�!?�W<��F�@}]��r�ٿ��T�3\�@�q4@讏�
�!?�W<��F�@}]��r�ٿ��T�3\�@�q4@讏�
�!?�W<��F�@�~'�.�ٿxbUT��@N`c%4@X���!?gqZ�@�~'�.�ٿxbUT��@N`c%4@X���!?gqZ�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@��L��ٿ2v�p�[�@��=�#4@�}��א!?ha�0x�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@'}mۦ�ٿ9���.E�@��!ލ4@�d	蕐!?�-��В�@ˌ�Dӈٿ��M����@�t�4@��!?G���#�@+��C�ٿ��T���@�����4@hn� �!?%�aO��@+��C�ٿ��T���@�����4@hn� �!?%�aO��@
@���ٿ�~K�6��@	�ͯ�4@|�j���!?��V71�@
@���ٿ�~K�6��@	�ͯ�4@|�j���!?��V71�@
@���ٿ�~K�6��@	�ͯ�4@|�j���!?��V71�@
@���ٿ�~K�6��@	�ͯ�4@|�j���!?��V71�@��^�ւٿNg��@�[ ƴ4@V��k�!?�����m�@��^�ւٿNg��@�[ ƴ4@V��k�!?�����m�@��^�ւٿNg��@�[ ƴ4@V��k�!?�����m�@��H	`�ٿ	��j��@�ȹm4@��徐!?��5���@��H	`�ٿ	��j��@�ȹm4@��徐!?��5���@��H	`�ٿ	��j��@�ȹm4@��徐!?��5���@��H	`�ٿ	��j��@�ȹm4@��徐!?��5���@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@��QŅٿ|�k��@�ʵ�4@ļ|�!?K(�/QL�@dpM�҈ٿ�v��5��@u6Y�4@n�*2�!?�W���@dpM�҈ٿ�v��5��@u6Y�4@n�*2�!?�W���@���ѽ�ٿ�	,t;�@U��e54@��;���!?�)`k~��@7�nh�ٿ�C v�;�@&+�4@7|�Ȑ!?��뗸x�@7�nh�ٿ�C v�;�@&+�4@7|�Ȑ!?��뗸x�@^��C��ٿ��|���@j�u�4@�c��ې!?׵"��@^��C��ٿ��|���@j�u�4@�c��ې!?׵"��@��Pׇٿ�7�WkM�@�Kl4@ߛD�!?�^���@��Pׇٿ�7�WkM�@�Kl4@ߛD�!?�^���@��Pׇٿ�7�WkM�@�Kl4@ߛD�!?�^���@u�k1�ٿ�+����@l��M�4@��;̻�!?�C^Wr�@u�k1�ٿ�+����@l��M�4@��;̻�!?�C^Wr�@u�k1�ٿ�+����@l��M�4@��;̻�!?�C^Wr�@u�k1�ٿ�+����@l��M�4@��;̻�!?�C^Wr�@u�k1�ٿ�+����@l��M�4@��;̻�!?�C^Wr�@`�[>p�ٿaG��t�@Y�M4@�;Z͐!?$�$�%��@�[�!��ٿ	�U ��@<�q4@��7��!?�Y�c<��@����ٿ����\��@`8t4@���G��!?,��{<	�@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@uX�B��ٿ}��-3��@�E��j4@RE���!?����?��@*�+ٿ�4�&��@j�.4@ؠF:��!?��q�b��@*�+ٿ�4�&��@j�.4@ؠF:��!?��q�b��@*�+ٿ�4�&��@j�.4@ؠF:��!?��q�b��@*�+ٿ�4�&��@j�.4@ؠF:��!?��q�b��@*�+ٿ�4�&��@j�.4@ؠF:��!?��q�b��@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@3�K!:�ٿ���c�@T�ul�4@K�ѹ�!?�u��(�@V�*Y�ٿ�O����@K��8�4@.UV��!?��ン��@V�*Y�ٿ�O����@K��8�4@.UV��!?��ン��@V�*Y�ٿ�O����@K��8�4@.UV��!?��ン��@V�*Y�ٿ�O����@K��8�4@.UV��!?��ン��@V�*Y�ٿ�O����@K��8�4@.UV��!?��ン��@�����ٿ4�+�D�@�'�4@�dn��!?i�Ӏ0��@�����ٿ4�+�D�@�'�4@�dn��!?i�Ӏ0��@�����ٿ4�+�D�@�'�4@�dn��!?i�Ӏ0��@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@�AE!��ٿ��h2z��@�|��4@0���!?Q�Z��i�@1ax���ٿ�nGz�@��h�4@%�Z�!?]�vF��@1ax���ٿ�nGz�@��h�4@%�Z�!?]�vF��@F�ZJ׊ٿ�8`j���@o��g 4@���ւ�!?ڸ����@F�ZJ׊ٿ�8`j���@o��g 4@���ւ�!?ڸ����@DJg��ٿ��~����@���4@k�9�Ԑ!?�S�����@DJg��ٿ��~����@���4@k�9�Ԑ!?�S�����@DJg��ٿ��~����@���4@k�9�Ԑ!?�S�����@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@>򁛥�ٿ�K��K�@�u���4@�#G&��!?YMö�@Ub�K�ٿ�����@�#}�~4@nv�!?�W��g�@"�ߪ�ٿ)�g D�@ 	��4@v@�`�!?��c��s�@"�ߪ�ٿ)�g D�@ 	��4@v@�`�!?��c��s�@Z�1BՌٿP��o�@�y�k4@K;�x��!?�ν	?}�@Z�1BՌٿP��o�@�y�k4@K;�x��!?�ν	?}�@Z�1BՌٿP��o�@�y�k4@K;�x��!?�ν	?}�@Z�1BՌٿP��o�@�y�k4@K;�x��!?�ν	?}�@B�Gǧ�ٿ���9'�@���4@��up�!?2@v|��@��R	�ٿ�<U)���@G$۵�4@�i���!?�O����@�qT�Նٿ;��#��@�^��4@�,j<�!?�8t�n��@�qT�Նٿ;��#��@�^��4@�,j<�!?�8t�n��@w�v3�ٿh*ʓf��@�鲴V4@��w���!?�7k?��@w�v3�ٿh*ʓf��@�鲴V4@��w���!?�7k?��@w�v3�ٿh*ʓf��@�鲴V4@��w���!?�7k?��@w�v3�ٿh*ʓf��@�鲴V4@��w���!?�7k?��@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�6U6��ٿ$H�7�@�@��ÒF4@ �Đ!?�K��;�@�+��ٿљ�Hk�@��=64@l�T��!?$����<�@�+��ٿљ�Hk�@��=64@l�T��!?$����<�@�+��ٿљ�Hk�@��=64@l�T��!?$����<�@���ٿ��Jl�@��4@�~h_��!?����K��@���ٿ��Jl�@��4@�~h_��!?����K��@���ٿ��Jl�@��4@�~h_��!?����K��@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@~�7i0�ٿe-��.��@+�p�<4@A��w��!?K��!h8�@,R1���ٿ�r��V9�@�.ޑ4@�*W���!?P%�>���@&�~�ٿ��)�@k u�I4@�Zj-��!?�گ/���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@0���,~ٿ��=��@<	`\� 4@m %@��!?+`%3���@.e-�)�ٿ�˽�uk�@���d� 4@!�L���!?K�zߖ�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@��vo�ٿ!�= �)�@
��W 4@G�jѐ!?�5B�@�A�^�ٿ!f���@�VT��3@�A���!?�N�����@�A�^�ٿ!f���@�VT��3@�A���!?�N�����@�A�^�ٿ!f���@�VT��3@�A���!?�N�����@e8��L�ٿ���k�C�@L���� 4@X���!?�@� �@u^��ٿ�bA�|��@e���$4@��~��!?z��� ��@u^��ٿ�bA�|��@e���$4@��~��!?z��� ��@u^��ٿ�bA�|��@e���$4@��~��!?z��� ��@��@r�ٿ�|�s�M�@����4@�����!?X�^���@��@r�ٿ�|�s�M�@����4@�����!?X�^���@��@r�ٿ�|�s�M�@����4@�����!?X�^���@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@V�wЏٿ�6����@���34@�.p�!?#kIa�@p���ٿ����@D�1��4@S��q�!?�e�κ��@p���ٿ����@D�1��4@S��q�!?�e�κ��@p���ٿ����@D�1��4@S��q�!?�e�κ��@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@h;���ٿ�[s���@�K��	4@� �ʐ!?6V�bD@�@�YMr�ٿ��d�@d�zh�4@w6-[�!?��V��D�@�YMr�ٿ��d�@d�zh�4@w6-[�!?��V��D�@�YMr�ٿ��d�@d�zh�4@w6-[�!?��V��D�@ ���h�ٿ��|~V�@�-�4@w2�죐!?oB�"/��@ZPtLO�ٿr�-lt�@��*�_4@�f	!?�SQ��@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�q~멆ٿ�F=5�c�@�c�4@�6j��!?�&��ђ�@�z�AG�ٿ��q��B�@�aFV4@�����!?�&c��@�z�AG�ٿ��q��B�@�aFV4@�����!?�&c��@�z�AG�ٿ��q��B�@�aFV4@�����!?�&c��@�3cd�ٿ��v)���@������3@	�����!?��g�w�@�3cd�ٿ��v)���@������3@	�����!?��g�w�@�3cd�ٿ��v)���@������3@	�����!?��g�w�@�3cd�ٿ��v)���@������3@	�����!?��g�w�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@�4��ٿ��R�y�@�^4@�?�֐!?���BJ�@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��LiщٿU$&#���@���uG4@=[NĐ!?(�7�w��@��Mkc�ٿ�A�� �@�U���4@��/`��!?�
>��@��Mkc�ٿ�A�� �@�U���4@��/`��!?�
>��@��Mkc�ٿ�A�� �@�U���4@��/`��!?�
>��@�+$�уٿ��\F���@X����4@�F��Y�!?�a����@�+$�уٿ��\F���@X����4@�F��Y�!?�a����@�h�7�ٿ� r}��@5�64@�d��t�!?
�>��@�h�7�ٿ� r}��@5�64@�d��t�!?
�>��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�e��4�ٿ��L��@�z)��4@�3�_2�!?��K!8��@�1Lq;�ٿ�s�C�@�y�R4@U��k�!?���`�O�@�1Lq;�ٿ�s�C�@�y�R4@U��k�!?���`�O�@�1Lq;�ٿ�s�C�@�y�R4@U��k�!?���`�O�@-3Z�1�ٿa,'�#�@�\=nw4@�%ߚW�!?�;K��<�@�B[@�ٿtι(��@uH�h4@*3�?}�!?l0����@�B[@�ٿtι(��@uH�h4@*3�?}�!?l0����@�B[@�ٿtι(��@uH�h4@*3�?}�!?l0����@�B[@�ٿtι(��@uH�h4@*3�?}�!?l0����@�}����ٿ��P%��@��O�4@T��1��!?�g�YԵ�@�}����ٿ��P%��@��O�4@T��1��!?�g�YԵ�@�}����ٿ��P%��@��O�4@T��1��!?�g�YԵ�@�}����ٿ��P%��@��O�4@T��1��!?�g�YԵ�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@;WC8��ٿtEn���@=Ɨ�Z4@�۱�!?����kT�@_r�u�ٿ�3��@�i��4@���ѐ!?:�e)hN�@_r�u�ٿ�3��@�i��4@���ѐ!?:�e)hN�@_r�u�ٿ�3��@�i��4@���ѐ!?:�e)hN�@_r�u�ٿ�3��@�i��4@���ѐ!?:�e)hN�@7���u�ٿY�w?�{�@�Qs�4@��`��!?�{���@�W���ٿ�ҺK���@���U4@���毐!?�au*ˇ�@�W���ٿ�ҺK���@���U4@���毐!?�au*ˇ�@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@�ʒ���ٿ��A_��@�#�+�4@�C�x��!?�������@��#2�ٿv�DU@��@n����4@������!?��Q'���@��#2�ٿv�DU@��@n����4@������!?��Q'���@V�7X��ٿ�����
�@~On4@���@�!?gm�/=`�@V�7X��ٿ�����
�@~On4@���@�!?gm�/=`�@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@8�qtd�ٿ�
\�2��@��+�4@����E�!?❙���@�����ٿL�n�_�@V!�]4@-"ם!�!?t����@	�{���ٿ�Q���o�@͕�:�4@�c� �!?̨";���@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�Ը3	�ٿr��j�@NaX4@����'�!?�z�ܐ��@�~U��~ٿ�c�%u�@(Ѥ��4@c��0�!?R8N� �@�~U��~ٿ�c�%u�@(Ѥ��4@c��0�!?R8N� �@�~U��~ٿ�c�%u�@(Ѥ��4@c��0�!?R8N� �@�~U��~ٿ�c�%u�@(Ѥ��4@c��0�!?R8N� �@�~U��~ٿ�c�%u�@(Ѥ��4@c��0�!?R8N� �@���Q��ٿ�H�S-�@��Rl�4@��:Y�!?{c��@���Q��ٿ�H�S-�@��Rl�4@��:Y�!?{c��@���Q��ٿ�H�S-�@��Rl�4@��:Y�!?{c��@���Q��ٿ�H�S-�@��Rl�4@��:Y�!?{c��@o����}ٿ�M��ޡ�@>l�K4@ş��!?&�jmXU�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@[�?T�|ٿ��qj�@3���4@D��w��!?�"�%�@����D~ٿF6���@8;�n4@����!?}kB�[�@����D~ٿF6���@8;�n4@����!?}kB�[�@����D~ٿF6���@8;�n4@����!?}kB�[�@����D~ٿF6���@8;�n4@����!?}kB�[�@̣aߕ|ٿ�vT���@��{4@��t�ʐ!?�����o�@�ꐵ�}ٿG�����@��G4@��'��!?��Ɵ[��@�ꐵ�}ٿG�����@��G4@��'��!?��Ɵ[��@�ꐵ�}ٿG�����@��G4@��'��!?��Ɵ[��@�ꐵ�}ٿG�����@��G4@��'��!?��Ɵ[��@�ꐵ�}ٿG�����@��G4@��'��!?��Ɵ[��@K��(�tٿ0x><��@�&-4�4@姭|��!?�c�1�@K��(�tٿ0x><��@�&-4�4@姭|��!?�c�1�@K��(�tٿ0x><��@�&-4�4@姭|��!?�c�1�@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@�,�}ٿQ����^�@��_n4@H�P���!?X{�?���@gm/(5ٿ�#��b�@�M@"4@�x굗�!??�c�@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@��${ٿNg�s�@a�R�4@��ɐ!?�
;?���@�ɇ.r�ٿ
t��Z�@��a��4@Un���!?�ϮE��@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@C��ٿ�r�=��@�M��A4@�~��Ȑ!?\de2ѓ�@�d���ٿZ�9�\�@�9�k4@Թ�4��!?�DU)�@�d���ٿZ�9�\�@�9�k4@Թ�4��!?�DU)�@�d���ٿZ�9�\�@�9�k4@Թ�4��!?�DU)�@�d���ٿZ�9�\�@�9�k4@Թ�4��!?�DU)�@S��[�ٿ�Q���@��G4@B��O�!?��43x��@S��[�ٿ�Q���@��G4@B��O�!?��43x��@S��[�ٿ�Q���@��G4@B��O�!?��43x��@u3ڟzٿN�����@���G�4@Zv����!?��=��l�@u3ڟzٿN�����@���G�4@Zv����!?��=��l�@u3ڟzٿN�����@���G�4@Zv����!?��=��l�@u3ڟzٿN�����@���G�4@Zv����!?��=��l�@�s����ٿ�";��@Y��� 4@��a��!?~,Q�U�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���!�ٿ]�+� �@���Q�4@�Ey ��!?&� 1�@���ٿ��@��@��QT4@%�B��!?N#v��p�@���ٿ��@��@��QT4@%�B��!?N#v��p�@���2,}ٿ�#�VA�@�q�Eg4@����Ӑ!?j
]͍�@��N}ٿ�&��!��@���<4@�����!?8��֫�@��dN�{ٿTµ����@���E4@���i��!?I@�q�z�@��dN�{ٿTµ����@���E4@���i��!?I@�q�z�@<����ٿ�l�R�;�@d��Kq4@�@u!�!?S���@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@,��t�ٿ�wے��@�5z�W4@�pKX	�!?x�
�m�@��3�ٿ2Ξ�H�@i� ��4@�c}�ѐ!?�!0*��@��3�ٿ2Ξ�H�@i� ��4@�c}�ѐ!?�!0*��@��3�ٿ2Ξ�H�@i� ��4@�c}�ѐ!?�!0*��@��tIj}ٿw�J��@'cY:�4@��8���!?���ׂ�@��tIj}ٿw�J��@'cY:�4@��8���!?���ׂ�@@�kN��ٿ��?��N�@���E�4@�	���!?l��O���@@�kN��ٿ��?��N�@���E�4@�	���!?l��O���@@�kN��ٿ��?��N�@���E�4@�	���!?l��O���@@�kN��ٿ��?��N�@���E�4@�	���!?l��O���@@�kN��ٿ��?��N�@���E�4@�	���!?l��O���@�e�ٿ�4J��(�@_<(4@����!?�V�6���@xGp��ٿ�s�Kz�@���<4@�-�ې!?���Y���@xGp��ٿ�s�Kz�@���<4@�-�ې!?���Y���@xGp��ٿ�s�Kz�@���<4@�-�ې!?���Y���@xGp��ٿ�s�Kz�@���<4@�-�ې!?���Y���@�6yP�ٿ����,�@�6(u�4@Ύ"q�!?c0���v�@\\��~ٿw0�`��@�}�l4@q����!?�AĖ��@\\��~ٿw0�`��@�}�l4@q����!?�AĖ��@\\��~ٿw0�`��@�}�l4@q����!?�AĖ��@�3���ٿ�#�z3��@f����4@S�{̐!?���M�@�3���ٿ�#�z3��@f����4@S�{̐!?���M�@�3���ٿ�#�z3��@f����4@S�{̐!?���M�@�3���ٿ�#�z3��@f����4@S�{̐!?���M�@�3���ٿ�#�z3��@f����4@S�{̐!?���M�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@����ٿ�a���@��v+24@��8��!?3M/.�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@������ٿ��"U{�@X��}4@���}ސ!?���e�@�w`���ٿК�����@+h}��4@�\"��!?@�n)�@�w`���ٿК�����@+h}��4@�\"��!?@�n)�@@��׈ٿ��ۡ3�@]�8N)
4@�|�X��!?1Ut�DO�@Q�MX��ٿ;���@�̧4@�U6&ǐ!?)� �Ps�@Q�MX��ٿ;���@�̧4@�U6&ǐ!?)� �Ps�@Q�MX��ٿ;���@�̧4@�U6&ǐ!?)� �Ps�@Q�MX��ٿ;���@�̧4@�U6&ǐ!?)� �Ps�@�F�^�ٿВF���@���1�4@/XA�!?��<����@�F�^�ٿВF���@���1�4@/XA�!?��<����@��+��ٿ����@PB���4@~����!?�z�ER��@��+��ٿ����@PB���4@~����!?�z�ER��@�#VT}ٿE�*D��@Gp�4@@-؉�!?R��ͨ��@�#VT}ٿE�*D��@Gp�4@@-؉�!?R��ͨ��@�#VT}ٿE�*D��@Gp�4@@-؉�!?R��ͨ��@Z��1�ٿ�{����@���k	4@C+��!?�
��@Z��1�ٿ�{����@���k	4@C+��!?�
��@Z��1�ٿ�{����@���k	4@C+��!?�
��@Z��1�ٿ�{����@���k	4@C+��!?�
��@~"J���ٿ���(uF�@���g|4@LB��!?�I��@l��p��ٿ�1|���@Q��4@�'H^�!?���퐛�@l��p��ٿ�1|���@Q��4@�'H^�!?���퐛�@���[��ٿ�,�p��@�i4@)�����!?�m�Nڧ�@���[��ٿ�,�p��@�i4@)�����!?�m�Nڧ�@���[��ٿ�,�p��@�i4@)�����!?�m�Nڧ�@�#6���ٿ/���Ī�@����4@n��>�!??\Vh���@�#6���ٿ/���Ī�@����4@n��>�!??\Vh���@�#6���ٿ/���Ī�@����4@n��>�!??\Vh���@�#6���ٿ/���Ī�@����4@n��>�!??\Vh���@����*�ٿ�W��{�@n�ɩj4@V~���!?@�g�@����*�ٿ�W��{�@n�ɩj4@V~���!?@�g�@����*�ٿ�W��{�@n�ɩj4@V~���!?@�g�@����*�ٿ�W��{�@n�ɩj4@V~���!?@�g�@����*�ٿ�W��{�@n�ɩj4@V~���!?@�g�@�/�*��ٿݚ��@�S�A,4@8[&[�!?�d�$�z�@�ֺ�ٿRO�Ǽ�@���4@د���!?��e^��@�ֺ�ٿRO�Ǽ�@���4@د���!?��e^��@�ֺ�ٿRO�Ǽ�@���4@د���!?��e^��@�ֺ�ٿRO�Ǽ�@���4@د���!?��e^��@�ֺ�ٿRO�Ǽ�@���4@د���!?��e^��@ֹ�+�ٿM.�ȴ*�@�AD	~4@g@{y�!?@�!��@ֹ�+�ٿM.�ȴ*�@�AD	~4@g@{y�!?@�!��@ֹ�+�ٿM.�ȴ*�@�AD	~4@g@{y�!?@�!��@ֹ�+�ٿM.�ȴ*�@�AD	~4@g@{y�!?@�!��@ֹ�+�ٿM.�ȴ*�@�AD	~4@g@{y�!?@�!��@�R�X�ٿ�;O����@�6��� 4@f?\.�!?NnWl���@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@k1��i�ٿ���/��@�5Z@�4@5�� �!?s����Q�@ߣ�n�ٿ�`���A�@�%�4@�O����!?H�;���@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@tC`��ٿ��7����@��)�4@��\Y�!?OF��@�6aa�ٿ��=M
��@��z��4@YWw�!?l����@�N��>�ٿg�Q�H�@�d"�4@����D�!?r�m@T}�@�N��>�ٿg�Q�H�@�d"�4@����D�!?r�m@T}�@�N��>�ٿg�Q�H�@�d"�4@����D�!?r�m@T}�@�N��>�ٿg�Q�H�@�d"�4@����D�!?r�m@T}�@����ٿ$k�W�@֦�4@�.1#�!?�B]����@����ٿ$k�W�@֦�4@�.1#�!?�B]����@����ٿ$k�W�@֦�4@�.1#�!?�B]����@����ٿ$k�W�@֦�4@�.1#�!?�B]����@����ٿ$k�W�@֦�4@�.1#�!?�B]����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@�\p��ٿ|�푼��@�*j*j4@DɎ�6�!?�����@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@uE���|ٿ��ͤ��@�/u��4@qSXސ!?�E���@A%��ٿ��}���@b�X&4@�l��ߐ!?�.�Rb�@A%��ٿ��}���@b�X&4@�l��ߐ!?�.�Rb�@���Ix�ٿ�Jǜ_��@Ymx4@%�@\"�!?ư�V��@���Ix�ٿ�Jǜ_��@Ymx4@%�@\"�!?ư�V��@���Ix�ٿ�Jǜ_��@Ymx4@%�@\"�!?ư�V��@���Ix�ٿ�Jǜ_��@Ymx4@%�@\"�!?ư�V��@���yʃٿ@0S��#�@W�﮵4@lɬ2А!?"0��j��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@>��҈ٿ��ic��@֚c��4@�6�8{�!? �d-1��@u�~٦�ٿ������@�B3�4@Ħ*E��!?��Y���@l~_�l�ٿ��qs��@��h4@�U�)�!?����)��@���s�ٿ~�&���@W��\�4@d<���!?j{�a{`�@���s�ٿ~�&���@W��\�4@d<���!?j{�a{`�@���s�ٿ~�&���@W��\�4@d<���!?j{�a{`�@���s�ٿ~�&���@W��\�4@d<���!?j{�a{`�@T�z��ٿ~G�� �@�Y��4@��:Đ!?��ݍX��@T�z��ٿ~G�� �@�Y��4@��:Đ!?��ݍX��@T�z��ٿ~G�� �@�Y��4@��:Đ!?��ݍX��@T�z��ٿ~G�� �@�Y��4@��:Đ!?��ݍX��@T�z��ٿ~G�� �@�Y��4@��:Đ!?��ݍX��@��j�ٿ��6��@d��F�4@b�!?J9�#��@�?��m�ٿ���p�@g�CHI4@�઼�!?�)�D��@�?��m�ٿ���p�@g�CHI4@�઼�!?�)�D��@�?��m�ٿ���p�@g�CHI4@�઼�!?�)�D��@�?��m�ٿ���p�@g�CHI4@�઼�!?�)�D��@�?��m�ٿ���p�@g�CHI4@�઼�!?�)�D��@�Elg�ٿ_�ܠ���@�����4@�<���!?�����@�Elg�ٿ_�ܠ���@�����4@�<���!?�����@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@��g��ٿu*�b��@pQF�4@x�v���!?�P���A�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@3&dƃ�ٿ�/5շ�@�)��4@�ߵ��!?��S\�@��هٿX����$�@�X��T4@ǿ;���!?��O3�@��هٿX����$�@�X��T4@ǿ;���!?��O3�@��هٿX����$�@�X��T4@ǿ;���!?��O3�@��هٿX����$�@�X��T4@ǿ;���!?��O3�@��هٿX����$�@�X��T4@ǿ;���!?��O3�@�V���ٿ׻� ���@FJ6�c4@��a�!?��l�q�@Su���}ٿ�Ɔ#5��@ �SA4@�~~"�!?6M�{'��@Su���}ٿ�Ɔ#5��@ �SA4@�~~"�!?6M�{'��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@��N�σٿ� k�98�@�*��4@Yts���!?z.� o��@�ݎaD�ٿ"W�����@Ӽh4@�Е*�!?���AAN�@�ݎaD�ٿ"W�����@Ӽh4@�Е*�!?���AAN�@�ݎaD�ٿ"W�����@Ӽh4@�Е*�!?���AAN�@)��$��ٿ� �U�@���E# 4@��%�!?J�bB�@)��$��ٿ� �U�@���E# 4@��%�!?J�bB�@��u!ÏٿL2m5Q_�@�4��4@�}0|�!?�淯�|�@Pjɭ-�ٿ�P�j���@ZN|I~4@�b��E�!?W샛x�@��_��ٿς����@���:14@
Rw[�!?�MN�ӱ�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@�l~�4�ٿGn�wn�@9�x�4@ez���!?�E�Zm2�@$-���ٿw�l^x�@����4@@��r��!?����}�@$-���ٿw�l^x�@����4@@��r��!?����}�@$-���ٿw�l^x�@����4@@��r��!?����}�@���ٿ�j�+��@�D�4@&�r�0�!?_�`���@!p7�ٿڀ�Ť�@�|���4@Ć��ݐ!?d!�ؤ,�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@p���A�ٿ��FD���@��>�4@{��J��!?qm^q�?�@��̊ٿ���Ԧ�@�R
4@������!?�U�����@��G�͈ٿSa$�5j�@�֢��4@���ժ�!?��j�h��@��G�͈ٿSa$�5j�@�֢��4@���ժ�!?��j�h��@��G�͈ٿSa$�5j�@�֢��4@���ժ�!?��j�h��@CWf'�ٿ�%��u��@����4@��V¸�!?�G^mw�@CWf'�ٿ�%��u��@����4@��V¸�!?�G^mw�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@�J��g�ٿ!�G�D�@����4@��R���!?��C��o�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@��3~,�ٿ���j���@|kc,4@��J�;�!?QL�0�@�@^��("~ٿ��;��@�>%r�4@
E��!?@JK4j6�@^��("~ٿ��;��@�>%r�4@
E��!?@JK4j6�@^��("~ٿ��;��@�>%r�4@
E��!?@JK4j6�@^��("~ٿ��;��@�>%r�4@
E��!?@JK4j6�@�sEF~ٿ��J��e�@䲏��4@j��8ސ!?8��0s�@�sEF~ٿ��J��e�@䲏��4@j��8ސ!?8��0s�@�����ٿI\��mY�@�|�4@�k��!?a�+z!�@�����ٿI\��mY�@�|�4@�k��!?a�+z!�@�����ٿI\��mY�@�|�4@�k��!?a�+z!�@*s-G	�ٿ�X~����@_B�Y�4@�r�C�!?������@��?�~ٿ"��B#U�@�Ǜ�4@t���!?�f,�N��@�"nb�ٿ)���@���4@�D����!?2��yTY�@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@��Q���ٿv��Ο�@H����4@�i?���!?�O:���@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@�:^�ٿy� �_�@� �&�4@��*r��!?�>�\	�@)��b�ٿ3�o���@��j*~4@���୐!?N������@)��b�ٿ3�o���@��j*~4@���୐!?N������@)��b�ٿ3�o���@��j*~4@���୐!?N������@)��b�ٿ3�o���@��j*~4@���୐!?N������@�.WMM�ٿ�os��	�@�%q�C4@�'��!?��ƴ0�@�.WMM�ٿ�os��	�@�%q�C4@�'��!?��ƴ0�@���ŅٿU����@�A�y4@`�S��!?:U�:J�@���ŅٿU����@�A�y4@`�S��!?:U�:J�@���ŅٿU����@�A�y4@`�S��!?:U�:J�@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�!��6�ٿx��T���@�+=4@%u,��!?b��@�"l���ٿ:��V��@�^LI�4@�EG�!?��|u�*�@�6Π)�ٿ͉�l��@q�;x�4@�Nѐ!?�Zs�٤�@
�Ԋٿ)z����@V[��4@LPג��!?��;\po�@
�Ԋٿ)z����@V[��4@LPג��!?��;\po�@
�Ԋٿ)z����@V[��4@LPג��!?��;\po�@
�Ԋٿ)z����@V[��4@LPג��!?��;\po�@
�Ԋٿ)z����@V[��4@LPג��!?��;\po�@�����ٿ�	���<�@���Q�	4@����{�!?��tFf�@�����ٿ�	���<�@���Q�	4@����{�!?��tFf�@�����ٿ�	���<�@���Q�	4@����{�!?��tFf�@�����ٿ�	���<�@���Q�	4@����{�!?��tFf�@0H�чٿ���;N��@w]�B-4@��9��!?��z&��@0H�чٿ���;N��@w]�B-4@��9��!?��z&��@0H�чٿ���;N��@w]�B-4@��9��!?��z&��@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@� x���ٿ��ʝ��@�q>�4@� 2U��!?��/���@�~���ٿ	�g.���@_�(�4@
��c�!?�`l�	�@�~���ٿ	�g.���@_�(�4@
��c�!?�`l�	�@�iu�ٿ\K�6��@l?Q04@)�Kp^�!?:�R�r�@�iu�ٿ\K�6��@l?Q04@)�Kp^�!?:�R�r�@��`Ij�ٿ�2-9���@Ӄ�4@�	ʐ!?A�σ�)�@]YI�ٿK����!�@j}4@�qQ[?�!?�䟢��@]YI�ٿK����!�@j}4@�qQ[?�!?�䟢��@]YI�ٿK����!�@j}4@�qQ[?�!?�䟢��@�UfE~~ٿ��m%��@S_4@��r�Ґ!?�£�`��@�UfE~~ٿ��m%��@S_4@��r�Ґ!?�£�`��@�UfE~~ٿ��m%��@S_4@��r�Ґ!?�£�`��@�UfE~~ٿ��m%��@S_4@��r�Ґ!?�£�`��@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@?��捀ٿ�I���z�@��`ҵ4@*��̐!?c;5�~�@�:��0~ٿG�L����@�\C�4@�ׇ���!?�H�(Y��@�:��0~ٿG�L����@�\C�4@�ׇ���!?�H�(Y��@�LJ��ٿ�8B�ӊ�@f,�e-4@���А!?�hn���@�LJ��ٿ�8B�ӊ�@f,�e-4@���А!?�hn���@�LJ��ٿ�8B�ӊ�@f,�e-4@���А!?�hn���@�LJ��ٿ�8B�ӊ�@f,�e-4@���А!?�hn���@�LJ��ٿ�8B�ӊ�@f,�e-4@���А!?�hn���@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@��q��ٿUBU��@QK�O4@d��e��!?�A ��@����҅ٿ��=�|�@{�Fz�4@Fr-���!?G�a����@����҅ٿ��=�|�@{�Fz�4@Fr-���!?G�a����@����҅ٿ��=�|�@{�Fz�4@Fr-���!?G�a����@��9�ٿ���cp�@��&�R4@��>�ΐ!?� QqX��@��9�ٿ���cp�@��&�R4@��>�ΐ!?� QqX��@��9�ٿ���cp�@��&�R4@��>�ΐ!?� QqX��@�nfF͑ٿk�|�!�@cܭ4@���͐!?�p�Q���@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@⍎��ٿJdJxAg�@p�!v4@�%��!?��9�� �@c�
��ٿ��s�+��@��R.4@ U�b��!?0�ūd�@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�t|�{�ٿ�(�â�@�Ѣ�84@x!���!?[g���@�I����ٿ�a���@�nq��4@	�;�ѐ!?��|#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@7ݍ�Z�ٿb�!O��@ =��W4@�%Y�Đ!?�o�V�#�@P9����ٿi�,gNR�@O�R4@i� ~ڐ!?�eˏ�r�@P9����ٿi�,gNR�@O�R4@i� ~ڐ!?�eˏ�r�@P9����ٿi�,gNR�@O�R4@i� ~ڐ!?�eˏ�r�@P9����ٿi�,gNR�@O�R4@i� ~ڐ!?�eˏ�r�@P9����ٿi�,gNR�@O�R4@i� ~ڐ!?�eˏ�r�@+1�,4ٿ���VS�@y�U�4@�4��!?It��Y��@+1�,4ٿ���VS�@y�U�4@�4��!?It��Y��@�>�yxٿ+��[-�@��A"�4@�0-��!?K���@֋{�7}ٿ'+{��F�@94b�L4@N�����!?�{8���@֋{�7}ٿ'+{��F�@94b�L4@N�����!?�{8���@B�~Wiyٿ��8g���@`}���4@���l�!?OB�ӤZ�@B�~Wiyٿ��8g���@`}���4@���l�!?OB�ӤZ�@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@h�r\�ٿ�4�1X)�@�&�:W4@r�Ie��!?e�a����@x�'؀ٿ{������@Y���4@���.��!?੉Q(Q�@X.V��ٿR��)���@�G�
4@�x�VȐ!?^.sr�Q�@X.V��ٿR��)���@�G�
4@�x�VȐ!?^.sr�Q�@X.V��ٿR��)���@�G�
4@�x�VȐ!?^.sr�Q�@X.V��ٿR��)���@�G�
4@�x�VȐ!?^.sr�Q�@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@	�x��}ٿ�_3Ѧ�@P'���4@-�ߐ!?g�T�>��@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@� C[Ɔٿ�j�ɦ��@?}p	4@����|�!?윁���@�8Λٿc�c'�@w���<4@��'S�!?
��q��@�8Λٿc�c'�@w���<4@��'S�!?
��q��@�OL{�ٿ���'Qx�@��F�;4@Ey?�!?W��$�@�OL{�ٿ���'Qx�@��F�;4@Ey?�!?W��$�@�OL{�ٿ���'Qx�@��F�;4@Ey?�!?W��$�@P�"�ٿO�pB���@��R�74@����`�!?�m��}��@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@&�o�ٿG�>�A�@K�9��4@�����!?�����@��҆ٿ��#W/}�@��R�	4@n��1��!?�:�z�Z�@��҆ٿ��#W/}�@��R�	4@n��1��!?�:�z�Z�@��҆ٿ��#W/}�@��R�	4@n��1��!?�:�z�Z�@��҆ٿ��#W/}�@��R�	4@n��1��!?�:�z�Z�@��҆ٿ��#W/}�@��R�	4@n��1��!?�:�z�Z�@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@�R��D�ٿ���O�@��	4@0ܦʐ!?�{�b���@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@ǩ���ٿqy\��e�@�ɚ�k4@�Y����!?0�ns�y�@���ٿ�����@w�X�'4@�$t�Ґ!?[�o0-!�@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@����ٿ}�Y��@����4@����!?|J�ڗ��@���g�ٿs<hAz��@᫚�@4@�m�*�!?U艀��@���g�ٿs<hAz��@᫚�@4@�m�*�!?U艀��@���g�ٿs<hAz��@᫚�@4@�m�*�!?U艀��@�q|��ٿ�f��a��@���m4@X"�x�!?�/��}��@��	Q��ٿ+2��\��@u��W4@�2e���!?Wʒ���@��	Q��ٿ+2��\��@u��W4@�2e���!?Wʒ���@8��~�ٿg�<�β�@�%�	4@�- �!?��)��@8��~�ٿg�<�β�@�%�	4@�- �!?��)��@gS�b�ٿ�C�U*��@$���4@��	��!?���t`��@9���*}ٿ11Y]R�@�Ubn�4@�F�ߐ!?E��J8�@�t�Jٿsfy<@�@�J�#�4@:�Хѐ!?����ӻ�@�t�Jٿsfy<@�@�J�#�4@:�Хѐ!?����ӻ�@�t�Jٿsfy<@�@�J�#�4@:�Хѐ!?����ӻ�@�t�Jٿsfy<@�@�J�#�4@:�Хѐ!?����ӻ�@�t�Jٿsfy<@�@�J�#�4@:�Хѐ!?����ӻ�@8v'ʓ�ٿ���;x�@���o4@(���!?�
`>�k�@8v'ʓ�ٿ���;x�@���o4@(���!?�
`>�k�@8v'ʓ�ٿ���;x�@���o4@(���!?�
`>�k�@8v'ʓ�ٿ���;x�@���o4@(���!?�
`>�k�@8v'ʓ�ٿ���;x�@���o4@(���!?�
`>�k�@\���p�ٿ�{�v؀�@a��4@��k��!?$T3x5��@\���p�ٿ�{�v؀�@a��4@��k��!?$T3x5��@\���p�ٿ�{�v؀�@a��4@��k��!?$T3x5��@�^���~ٿ\��g}�@ⷂ�7	4@?�]�ݐ!?�Ħj��@�^���~ٿ\��g}�@ⷂ�7	4@?�]�ݐ!?�Ħj��@_�q�~�ٿl���)��@��4@w����!?s�ߗ��@_�q�~�ٿl���)��@��4@w����!?s�ߗ��@�R[��}ٿYR��)�@JY��4@���SА!?�i��Zv�@�R[��}ٿYR��)�@JY��4@���SА!?�i��Zv�@����ٿ��\}n�@O<�#4@����!?��-��@����ٿ��\}n�@O<�#4@����!?��-��@����ٿ��\}n�@O<�#4@����!?��-��@�DY�zٿh��7$�@���4@5��!?z�OЖ�@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@<t|��ٿXI����@3|p8p4@��d��!?me����@�e��T�ٿ������@��t�4@j_̓�!?��٬J�@�e��T�ٿ������@��t�4@j_̓�!?��٬J�@�e��T�ٿ������@��t�4@j_̓�!?��٬J�@�e��T�ٿ������@��t�4@j_̓�!?��٬J�@�e��T�ٿ������@��t�4@j_̓�!?��٬J�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@"r���ٿ�?E"�P�@?��*24@����t�!?�O\*�@.)3wp�ٿ⹡��@�ky�4@q��Ր!?m��܊Z�@.)3wp�ٿ⹡��@�ky�4@q��Ր!?m��܊Z�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@/���h�ٿ�kMՑD�@��8WP4@2����!?��󀩍�@MM��D�ٿ`A��/�@"ꧏ4@�S�4�!?�<��eP�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@�� ̆ٿ����v�@����n4@^(}��!?X?�l�U�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@T;'ׅٿ݉7#��@T�:߻4@���軐!?���'p�@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@ox�Ąٿ����n�@�8���3@�)���!?$̆��@#�޾u�ٿ.��5|z�@bΌ���3@��n���!?K��2�+�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@a�8�ٿu�����@�ۣ3�4@:Q�c�!?%yQP�'�@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@���ٿ5�h�s�@���|4@�B���!?X�{��@�L��ٿ����E�@�&��4@��+А!?e�U����@�L��ٿ����E�@�&��4@��+А!?e�U����@�vW��ٿ%D��C�@���vk4@a����!?��\��#�@�vW��ٿ%D��C�@���vk4@a����!?��\��#�@�vW��ٿ%D��C�@���vk4@a����!?��\��#�@u.��ٿ>�	!�@�Z�4@(C��!?YZq�Y�@���iՊٿ6,4P)��@֔~Ek4@H�����!?�����@���iՊٿ6,4P)��@֔~Ek4@H�����!?�����@���iՊٿ6,4P)��@֔~Ek4@H�����!?�����@���q^�ٿc~�k��@+�n�b4@k����!?�� �D�@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@��ϝ��ٿ?�H%r��@O�{E4@N	����!?�T��u��@�L砀ٿE@���*�@:��[!4@� V��!?.J���@�L砀ٿE@���*�@:��[!4@� V��!?.J���@�L砀ٿE@���*�@:��[!4@� V��!?.J���@�L砀ٿE@���*�@:��[!4@� V��!?.J���@�L砀ٿE@���*�@:��[!4@� V��!?.J���@c'��9ٿ]��"�-�@���4@��*��!?���S4m�@c'��9ٿ]��"�-�@���4@��*��!?���S4m�@{�]P�ٿ4|I��b�@�?�,�4@OP��!?��Ds@L�@{�]P�ٿ4|I��b�@�?�,�4@OP��!?��Ds@L�@{�]P�ٿ4|I��b�@�?�,�4@OP��!?��Ds@L�@{�]P�ٿ4|I��b�@�?�,�4@OP��!?��Ds@L�@��Ȃٿc=I�'��@�BJ[4@������!?��XQT�@��Ȃٿc=I�'��@�BJ[4@������!?��XQT�@��Ȃٿc=I�'��@�BJ[4@������!?��XQT�@��Ȃٿc=I�'��@�BJ[4@������!?��XQT�@��Ȃٿc=I�'��@�BJ[4@������!?��XQT�@H7��ٿ�h
�O��@��f�z4@~���u�!?{5��B��@H7��ٿ�h
�O��@��f�z4@~���u�!?{5��B��@�K�y}ٿ���5���@sNKa�	4@��M�v�!?R�zz�@p(��hzٿ�P�2\T�@=n4@c�Yb�!?>�f�,�@� 4}ٿw�.�k��@�
��%4@��L�&�!?��n��t�@� 4}ٿw�.�k��@�
��%4@��L�&�!?��n��t�@� 4}ٿw�.�k��@�
��%4@��L�&�!?��n��t�@� 4}ٿw�.�k��@�
��%4@��L�&�!?��n��t�@� 4}ٿw�.�k��@�
��%4@��L�&�!?��n��t�@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@)�����ٿV_$\��@![�4@5ܖd��!?�d�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@�$��чٿWGHF���@FT{{4@��]?�!?�����@��ׂ��ٿ��+@a��@�����4@���X�!?�]��s�@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@8��Z�ٿ�%Ϟ�/�@�SE�	4@� hJ�!?0�:@H��@f��}�ٿґ���.�@"�.R4@�:�j�!?Ԑ��}�@l-[.�ٿ|C�H��@�8��4@|�����!?2yh�K�@l-[.�ٿ|C�H��@�8��4@|�����!?2yh�K�@l-[.�ٿ|C�H��@�8��4@|�����!?2yh�K�@l-[.�ٿ|C�H��@�8��4@|�����!?2yh�K�@��X�.�ٿ؝o#J�@ŝ'�D4@�?�!?B�h�V��@��X�.�ٿ؝o#J�@ŝ'�D4@�?�!?B�h�V��@��X�.�ٿ؝o#J�@ŝ'�D4@�?�!?B�h�V��@:(�Q<�ٿ՗H?0�@�&��q4@�uj�Ґ!?����٥�@�ԣ��ٿ�� T���@��V�&4@��$;�!?,�����@�(���ٿ҃|@[�@2�[؃4@6/�B�!?.#�4��@�(���ٿ҃|@[�@2�[؃4@6/�B�!?.#�4��@�(���ٿ҃|@[�@2�[؃4@6/�B�!?.#�4��@�(���ٿ҃|@[�@2�[؃4@6/�B�!?.#�4��@�(���ٿ҃|@[�@2�[؃4@6/�B�!?.#�4��@��0ڞ�ٿl��'b�@����T4@����R�!?賆�(�@�֋�ٿ����7�@1����4@�c�}�!?bU.C��@Y�۶��ٿi,�Ԡ��@�����4@���!?^.�u��@Y�۶��ٿi,�Ԡ��@�����4@���!?^.�u��@Y�۶��ٿi,�Ԡ��@�����4@���!?^.�u��@Y�۶��ٿi,�Ԡ��@�����4@���!?^.�u��@@���ٿ�B7B�)�@��Võ4@�uS��!?�Ů�=�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@gD���ٿ��sw��@$H�Ҳ4@�|�֐!?����)�@��=��ٿ�9�d��@��)l 4@y*"%k�!?ztm� ��@�/����ٿ���d ��@�W]���3@].�&��!?�t�$�@X���ٿ�@c-.��@�z& 4@�3Wѣ�!?�Ϫ�c�@X���ٿ�@c-.��@�z& 4@�3Wѣ�!?�Ϫ�c�@X���ٿ�@c-.��@�z& 4@�3Wѣ�!?�Ϫ�c�@�S��ٿ.�XWaE�@6e��
4@�Yy��!?�tkT?��@�;L�ٿ㞕	�_�@�9�t4@�F8��!?4�
�v�@�;L�ٿ㞕	�_�@�9�t4@�F8��!?4�
�v�@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@+�!�9�ٿ�����@j�o4@ö���!?Y�/�P��@�R�ٿ���DK�@}~��4@hiO<�!?��O>
k�@VĠjE�ٿ`��_�@�D��F4@qs�8�!?b~���@VĠjE�ٿ`��_�@�D��F4@qs�8�!?b~���@VĠjE�ٿ`��_�@�D��F4@qs�8�!?b~���@VĠjE�ٿ`��_�@�D��F4@qs�8�!?b~���@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@	<�	b�ٿ_@�iC�@4����4@�yVG��!?���X,�@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�yHoψٿ"� k���@y�I�74@���ؐ!?a�����@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@�"c��ٿgAX��@=Fw�4@e�����!?��e�E�@���X�ٿ�5Tc�@WL��4@��k3%�!?�#kF!�@���X�ٿ�5Tc�@WL��4@��k3%�!?�#kF!�@���X�ٿ�5Tc�@WL��4@��k3%�!?�#kF!�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��ʙq�ٿN��e��@F��4@\����!?+�J�@��7tu�ٿ :e��%�@t�kI4@�� ��!?����@n�m=9�ٿ��-�@F���4@��x���!?��ف� �@n�m=9�ٿ��-�@F���4@��x���!?��ف� �@n�m=9�ٿ��-�@F���4@��x���!?��ف� �@n�m=9�ٿ��-�@F���4@��x���!?��ف� �@m��ǁٿHTO<��@���ry4@����!?h�{1��@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@(^^!�ٿ�Ҡyu��@��% c4@�n-��!?c��T�9�@��B�ٿ)��Y��@܍��4@箤��!?:�=q���@��B�ٿ)��Y��@܍��4@箤��!?:�=q���@��B�ٿ)��Y��@܍��4@箤��!?:�=q���@��B�ٿ)��Y��@܍��4@箤��!?:�=q���@� �ϙ�ٿ/�ٝ6&�@���4@��ː!?KN�fv��@� �ϙ�ٿ/�ٝ6&�@���4@��ː!?KN�fv��@0��b��ٿ�dI�c��@�ȧ4@7�;W̐!?pRX�J�@0��b��ٿ�dI�c��@�ȧ4@7�;W̐!?pRX�J�@0��b��ٿ�dI�c��@�ȧ4@7�;W̐!?pRX�J�@c��}ٿX �:�@D�vi84@��jь�!?ǉ;7x��@t��h�ٿk:�����@f&��4@�I��!?�ϿW�@t��h�ٿk:�����@f&��4@�I��!?�ϿW�@t��h�ٿk:�����@f&��4@�I��!?�ϿW�@t��h�ٿk:�����@f&��4@�I��!?�ϿW�@t��h�ٿk:�����@f&��4@�I��!?�ϿW�@J0���ٿ�_�;��@��*�� 4@���J"�!?�?�Jd�@J0���ٿ�_�;��@��*�� 4@���J"�!?�?�Jd�@J0���ٿ�_�;��@��*�� 4@���J"�!?�?�Jd�@o����~ٿ �\���@���\4@�SNgG�!?|��܈�@r�>�e|ٿΒ@�i�@�ٚ�}4@�R}5�!?M֊֊U�@r�>�e|ٿΒ@�i�@�ٚ�}4@�R}5�!?M֊֊U�@r�>�e|ٿΒ@�i�@�ٚ�}4@�R}5�!?M֊֊U�@r�>�e|ٿΒ@�i�@�ٚ�}4@�R}5�!?M֊֊U�@�{� H�ٿ6���8��@�EJ�4@��cݐ!?>K(�@	�@�{� H�ٿ6���8��@�EJ�4@��cݐ!?>K(�@	�@2ʰ���ٿ�2)ax4�@����Y4@�'�
ِ!?ei?f�O�@�� D{ٿ�Ԩ{��@�-4@�:=:q�!?)�*f���@�� D{ٿ�Ԩ{��@�-4@�:=:q�!?)�*f���@ ��s�ٿe7O�X�@�e~�v4@�M�2ʐ!?,̰;6H�@ ��s�ٿe7O�X�@�e~�v4@�M�2ʐ!?,̰;6H�@ ��s�ٿe7O�X�@�e~�v4@�M�2ʐ!?,̰;6H�@ ��s�ٿe7O�X�@�e~�v4@�M�2ʐ!?,̰;6H�@����ٿ��+�jz�@#�i��4@s���r�!?"a>���@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@�X�iG~ٿ��(59��@�ġn�4@(Hs��!?�	��G�@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@��W�ٿ�zJ��@��W!�4@��ۢ�!?%�����@T���ōٿO<����@��=14@�4D�!?�)t&�N�@��q���ٿ�	�}��@3�Uk4@��o[�!?��$p=�@��q���ٿ�	�}��@3�Uk4@��o[�!?��$p=�@��q���ٿ�	�}��@3�Uk4@��o[�!?��$p=�@��q���ٿ�	�}��@3�Uk4@��o[�!?��$p=�@��q���ٿ�	�}��@3�Uk4@��o[�!?��$p=�@��t�c�ٿ.鼰���@"�U6�4@;��2 �!?�Xr���@��t�c�ٿ.鼰���@"�U6�4@;��2 �!?�Xr���@��t�c�ٿ.鼰���@"�U6�4@;��2 �!?�Xr���@_��b�ٿ�.���S�@�c��U4@��'�!?d/�T'��@_��b�ٿ�.���S�@�c��U4@��'�!?d/�T'��@_��b�ٿ�.���S�@�c��U4@��'�!?d/�T'��@_��b�ٿ�.���S�@�c��U4@��'�!?d/�T'��@�2�h��ٿ�Q1ߢ��@�G|R�4@���r�!?�QM:��@�2�h��ٿ�Q1ߢ��@�G|R�4@���r�!?�QM:��@�2�h��ٿ�Q1ߢ��@�G|R�4@���r�!?�QM:��@�2�h��ٿ�Q1ߢ��@�G|R�4@���r�!?�QM:��@-'x�ٿ��3k�@|�1a�4@ª5U�!?�T��&��@���^�ٿ��͆�@��T4@�QGOv�!?C�����@¬�\�ٿg�C`��@ڤp @4@��[.��!?�0��u��@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�R�c��ٿ�&�΀�@f�!�|4@H�A���!?>|[�h�@�$�_�ٿ	DX���@��dM4@�K�;��!?�@-\��@�$�_�ٿ	DX���@��dM4@�K�;��!?�@-\��@\W˅ٿ��PsC�@]���4@q(���!?e�ͬ��@\W˅ٿ��PsC�@]���4@q(���!?e�ͬ��@\W˅ٿ��PsC�@]���4@q(���!?e�ͬ��@\W˅ٿ��PsC�@]���4@q(���!?e�ͬ��@��qU�|ٿm��8��@���B4@m�w��!?z������@��qU�|ٿm��8��@���B4@m�w��!?z������@��qU�|ٿm��8��@���B4@m�w��!?z������@��qU�|ٿm��8��@���B4@m�w��!?z������@��qU�|ٿm��8��@���B4@m�w��!?z������@{�`�n�ٿ���ˆ��@�CO��	4@�XF�9�!?�� x���@{�`�n�ٿ���ˆ��@�CO��	4@�XF�9�!?�� x���@{�`�n�ٿ���ˆ��@�CO��	4@�XF�9�!?�� x���@�����~ٿ��i��@�w�]�4@&��#
�!?�-<��@�����~ٿ��i��@�w�]�4@&��#
�!?�-<��@�����~ٿ��i��@�w�]�4@&��#
�!?�-<��@�����~ٿ��i��@�w�]�4@&��#
�!?�-<��@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@#��;��ٿ^�����@���aY4@�6�"�!?����N�@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@�$S�ٿ����w�@(ԑw�4@$�d�!?�tP+���@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@���,�ٿ�i����@W�Cq4@S�= �!?&f��]�@��}ɍٿ���)���@�u?�4@�"��4�!?�Љ���@��}ɍٿ���)���@�u?�4@�"��4�!?�Љ���@~���ٿ�2�T�@�&��	4@��W��!?�֬(d�@~���ٿ�2�T�@�&��	4@��W��!?�֬(d�@~���ٿ�2�T�@�&��	4@��W��!?�֬(d�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@��N�ٿ3d��/U�@�Q�/	4@"��!?R�?�<�@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@]i��3�ٿ(�רlJ�@�y㗕4@{�[��!?5�ؕ���@����ٿ��ɧH�@�-���4@B����!?bZկ-�@����ٿ��ɧH�@�-���4@B����!?bZկ-�@����ٿ��ɧH�@�-���4@B����!?bZկ-�@����ٿ��ɧH�@�-���4@B����!?bZկ-�@����ٿ��ɧH�@�-���4@B����!?bZկ-�@����ٿ��ɧH�@�-���4@B����!?bZկ-�@(M�)�ٿ��Л��@kT�J�4@��Ϩ��!?i�07��@(M�)�ٿ��Л��@kT�J�4@��Ϩ��!?i�07��@(M�)�ٿ��Л��@kT�J�4@��Ϩ��!?i�07��@$(�ށٿʸ�K��@l��H34@�|�V��!?����j��@$(�ށٿʸ�K��@l��H34@�|�V��!?����j��@$(�ށٿʸ�K��@l��H34@�|�V��!?����j��@$(�ށٿʸ�K��@l��H34@�|�V��!?����j��@m��`Z�ٿvlZ�@��@7��4@�/f���!?8A�MA5�@m��`Z�ٿvlZ�@��@7��4@�/f���!?8A�MA5�@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@�5��ٿ�X�B���@�ӒG4@ļ*��!?
�O����@в�۷�ٿ�%.����@���Hs4@��Ɛ!?�U���@f���T�ٿ�1��.��@Y,=�4@��ʜ�!?��m��@f���T�ٿ�1��.��@Y,=�4@��ʜ�!?��m��@f���T�ٿ�1��.��@Y,=�4@��ʜ�!?��m��@f���T�ٿ�1��.��@Y,=�4@��ʜ�!?��m��@-�?���ٿw���z^�@nc.).4@MO9%Ӑ!?������@-�?���ٿw���z^�@nc.).4@MO9%Ӑ!?������@�0�ȕٿC�����@C1�7z4@N&:ǐ!?۬�^8�@��<܀ٿE���I��@��g�p	4@�C?�ܐ!?�w����@��<܀ٿE���I��@��g�p	4@�C?�ܐ!?�w����@��<܀ٿE���I��@��g�p	4@�C?�ܐ!?�w����@��<܀ٿE���I��@��g�p	4@�C?�ܐ!?�w����@��<܀ٿE���I��@��g�p	4@�C?�ܐ!?�w����@m-H���ٿ��H�@	S9z4@:�W��!?�m�YT��@m-H���ٿ��H�@	S9z4@:�W��!?�m�YT��@+9_��ٿo��R(��@�t���4@j�|2��!?��Ϙ�@+9_��ٿo��R(��@�t���4@j�|2��!?��Ϙ�@+9_��ٿo��R(��@�t���4@j�|2��!?��Ϙ�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@���ٿ���8���@��.4@;�����!?�Y�N�p�@�j/ٿ�Y$��@�ɲr4@��l�!?#�`s���@�j/ٿ�Y$��@�ɲr4@��l�!?#�`s���@�j/ٿ�Y$��@�ɲr4@��l�!?#�`s���@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@�	��τٿ��f-���@�h�,4@�c�Y��!?�:��U��@W?F��ٿ�k��i��@{s���4@߂��ΐ!?6S�����@�+�g��ٿ�s�T�@�lo
�4@B��S�!?}B�p-�@�KLH��ٿ�������@�ik�N4@�؆��!?��sc���@�KLH��ٿ�������@�ik�N4@�؆��!?��sc���@�KLH��ٿ�������@�ik�N4@�؆��!?��sc���@%5�{ӈٿ�D^���@B�CE�4@��I�&�!?sx�>$�@�����ٿU��!M��@۞��4@f? ���!?�[L����@�����ٿU��!M��@۞��4@f? ���!?�[L����@�����ٿU��!M��@۞��4@f? ���!?�[L����@S�)R��ٿ�1W�<��@)��9g4@����y�!?��ö���@S�)R��ٿ�1W�<��@)��9g4@����y�!?��ö���@S�)R��ٿ�1W�<��@)��9g4@����y�!?��ö���@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@D팊ٿ��:����@�#'�4@;td��!?q�f^D��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@PO�Bۄٿ�0��W`�@��x;4@�yiu��!?TB?~2��@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@$���ٿ_[����@Jc�i	4@�+Zΐ!?F��+�!�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@ 5�t�ٿ%�����@�E�7�4@^z:��!?�)�A�+�@�d�w}ٿ����[��@�be^�4@�L3^�!?��$Ċp�@�d�w}ٿ����[��@�be^�4@�L3^�!?��$Ċp�@I�=���ٿ��0R�@.��J�4@�����!?�^���#�@I�=���ٿ��0R�@.��J�4@�����!?�^���#�@I�=���ٿ��0R�@.��J�4@�����!?�^���#�@I�=���ٿ��0R�@.��J�4@�����!?�^���#�@b����}ٿ�EҎ�.�@�&��&4@*纔�!?�z�����@b����}ٿ�EҎ�.�@�&��&4@*纔�!?�z�����@b����}ٿ�EҎ�.�@�&��&4@*纔�!?�z�����@b����}ٿ�EҎ�.�@�&��&4@*纔�!?�z�����@�����ٿn�G3��@[�%]	4@4#�Đ!? �OrH�@�����ٿn�G3��@[�%]	4@4#�Đ!? �OrH�@�����ٿn�G3��@[�%]	4@4#�Đ!? �OrH�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@>h5�w�ٿլkP��@ઠ+B
4@��!�Ð!?b"�@�Z��ٿI� ��B�@e��4@wKW��!?�fN��@�Z��ٿI� ��B�@e��4@wKW��!?�fN��@�o�4Z�ٿ����I��@{���4@���ߐ!?ݏ3���@�o�4Z�ٿ����I��@{���4@���ߐ!?ݏ3���@�o�4Z�ٿ����I��@{���4@���ߐ!?ݏ3���@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@�1V���ٿ�B���@�-EH�4@4�TԤ�!?F�[S�@=��.q�ٿp�)�@�)�;�4@h%�<��!?��c��@=��.q�ٿp�)�@�)�;�4@h%�<��!?��c��@=��.q�ٿp�)�@�)�;�4@h%�<��!?��c��@=��.q�ٿp�)�@�)�;�4@h%�<��!?��c��@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@I��V��ٿ�]2S��@���zx4@�+(���!?�0�a���@��ɇ�}ٿ'+�b���@N��B4@PJ�Ȑ!?��GIQ|�@��ɇ�}ٿ'+�b���@N��B4@PJ�Ȑ!?��GIQ|�@��ɇ�}ٿ'+�b���@N��B4@PJ�Ȑ!?��GIQ|�@��ɇ�}ٿ'+�b���@N��B4@PJ�Ȑ!?��GIQ|�@|f��ٿNN�<�@O�� 4@�����!?��ص�@|f��ٿNN�<�@O�� 4@�����!?��ص�@|f��ٿNN�<�@O�� 4@�����!?��ص�@|f��ٿNN�<�@O�� 4@�����!?��ص�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@�{cK�ٿ����#1�@I���%4@c��˝�!?� �(�G�@'�M0��ٿ���q�~�@�Up�4@��'��!?AAE���@'�M0��ٿ���q�~�@�Up�4@��'��!?AAE���@'�M0��ٿ���q�~�@�Up�4@��'��!?AAE���@'�M0��ٿ���q�~�@�Up�4@��'��!?AAE���@��
���ٿ��D���@Ӌ�C�	4@VAw���!?1ӳR*�@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@�bȃ�ٿ�Q�]-�@؉�D4@��Aʳ�!?��P���@.��Tb�ٿ�8(��9�@����4@��T4�!?�K����@.��Tb�ٿ�8(��9�@����4@��T4�!?�K����@.��Tb�ٿ�8(��9�@����4@��T4�!?�K����@.��Tb�ٿ�8(��9�@����4@��T4�!?�K����@.��Tb�ٿ�8(��9�@����4@��T4�!?�K����@m�0ᯊٿ�-i���@Qz�y�4@j�M��!?�;0�8�@m�0ᯊٿ�-i���@Qz�y�4@j�M��!?�;0�8�@m�0ᯊٿ�-i���@Qz�y�4@j�M��!?�;0�8�@m�0ᯊٿ�-i���@Qz�y�4@j�M��!?�;0�8�@!�,^؅ٿ��.�j5�@]k\4%4@(j�ϐ!?�+�|���@!�,^؅ٿ��.�j5�@]k\4%4@(j�ϐ!?�+�|���@!�,^؅ٿ��.�j5�@]k\4%4@(j�ϐ!?�+�|���@!�,^؅ٿ��.�j5�@]k\4%4@(j�ϐ!?�+�|���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@?x�Y��ٿ^I��R�@S��T�4@�z�s�!?	d�P���@� 1y�ٿ�Bͺ[t�@ڲD04@g���!?��	����@� 1y�ٿ�Bͺ[t�@ڲD04@g���!?��	����@� 1y�ٿ�Bͺ[t�@ڲD04@g���!?��	����@� 1y�ٿ�Bͺ[t�@ڲD04@g���!?��	����@� 1y�ٿ�Bͺ[t�@ڲD04@g���!?��	����@�Gd`��ٿ*	z<��@|��ͭ4@�TWʁ�!?t�[���@�Gd`��ٿ*	z<��@|��ͭ4@�TWʁ�!?t�[���@�Gd`��ٿ*	z<��@|��ͭ4@�TWʁ�!?t�[���@�$��ōٿ�/�g'��@6P:384@��@K�!?%�w��@�$��ōٿ�/�g'��@6P:384@��@K�!?%�w��@�$��ōٿ�/�g'��@6P:384@��@K�!?%�w��@�$��ōٿ�/�g'��@6P:384@��@K�!?%�w��@b�t�ٿ2ޮ)��@&�4@��`mb�!?-��G�@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@��ጌٿf��OY��@�Ƈ�4@@�|��!?!9��@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�ʮNڊٿ�&E�X�@��<4@��\��!?�Iʻ�T�@�)7��ٿ��P:n`�@6�.5� 4@�`DƐ!?ii�V5�@�)7��ٿ��P:n`�@6�.5� 4@�`DƐ!?ii�V5�@�)7��ٿ��P:n`�@6�.5� 4@�`DƐ!?ii�V5�@�)7��ٿ��P:n`�@6�.5� 4@�`DƐ!?ii�V5�@�)7��ٿ��P:n`�@6�.5� 4@�`DƐ!?ii�V5�@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@5@�j��ٿ����@��@[*�4@�N��ߐ!?�<��@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@�a,U�ٿ���Â�@�ذ9�4@�	��!?�k~���@��䆙�ٿ	��5f�@.��4@{�*"�!?�SA�+�@��䆙�ٿ	��5f�@.��4@{�*"�!?�SA�+�@L���ٿ�����@��4�^4@,���!?lkD����@L���ٿ�����@��4�^4@,���!?lkD����@L���ٿ�����@��4�^4@,���!?lkD����@l��&b�ٿ����:u�@��,
4@؛$͐!?6�œȧ�@��2f�ٿ��3���@���g	4@�*�Q��!?�(����@��2f�ٿ��3���@���g	4@�*�Q��!?�(����@��2f�ٿ��3���@���g	4@�*�Q��!?�(����@��2f�ٿ��3���@���g	4@�*�Q��!?�(����@r�A���ٿݩ�.�@K
��4@���!?[^!��@`�iW�ٿ��,�Ka�@��[�4@��`�!?�)��z�@�
8Qg{ٿ,'�k�@r�D$�4@�K����!?P�5��@�
8Qg{ٿ,'�k�@r�D$�4@�K����!?P�5��@�
8Qg{ٿ,'�k�@r�D$�4@�K����!?P�5��@�
8Qg{ٿ,'�k�@r�D$�4@�K����!?P�5��@���l'{ٿ׶�s��@Q�,^�4@?�ծܐ!?{�Q��@���l'{ٿ׶�s��@Q�,^�4@?�ծܐ!?{�Q��@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@u���Dxٿj�e��@�Dɪ�4@�8�%�!?+��Y�@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��R��}ٿz��n��@��9J4@h΅��!?�e@��@��*}ٿ��,�ib�@_)hf�4@�G ��!?�~�U;��@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@�ؿ#{ٿ|y�z>��@6��4@X�
��!?s�\ �@#~ٿ%<�;�@�`�=#4@�����!?qP�B~��@��ٿ>V$z��@ȕ_�4@�4W/��!?t�׮A��@��ٿ>V$z��@ȕ_�4@�4W/��!?t�׮A��@��ٿ>V$z��@ȕ_�4@�4W/��!?t�׮A��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@�ta]6�ٿ�d�
��@.~Y��4@����!?�n��"��@(��|Іٿ@JȔ�@�1���4@'�.y��!?t;�v��@(��|Іٿ@JȔ�@�1���4@'�.y��!?t;�v��@(��|Іٿ@JȔ�@�1���4@'�.y��!?t;�v��@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@P�d3j�ٿ��@r�5�@�{=�54@:7𝽐!?GQ�H�+�@����~�ٿ^!|J>�@����4@�z����!?d�>����@����~�ٿ^!|J>�@����4@�z����!?d�>����@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@w"�]�ٿ��#E�@�/E4@�P&Zϐ!?�1�i��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�M����ٿ������@��g�w4@��A��!?dr��@�Py�7�ٿ�v���b�@��9N4@2;Ӑ!?*�ܯ�Q�@�Py�7�ٿ�v���b�@��9N4@2;Ӑ!?*�ܯ�Q�@��С�ٿk��M{[�@�z܂�4@�[r��!?���h���@3Kܡ�ٿ�6P��@"C4@5����!?�98ns��@3Kܡ�ٿ�6P��@"C4@5����!?�98ns��@3Kܡ�ٿ�6P��@"C4@5����!?�98ns��@3Kܡ�ٿ�6P��@"C4@5����!?�98ns��@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@��F[�ٿ0 I�q��@X	N�4@TJ��!?�����@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@�@�ٿd��Y���@"i��4@��M,��!?�$:��-�@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@y#)�ٿ)P?��@�Ȣ��4@>�+���!?t|$���@��jV�ٿl�����@j��,94@|�y"{�!?$��K��@��jV�ٿl�����@j��,94@|�y"{�!?$��K��@��͉�ٿ�3�����@�ڣ4@c�[��!?;����@��͉�ٿ�3�����@�ڣ4@c�[��!?;����@w���ٿJ��-a�@�k�T4@�;Z.̐!?�����+�@w���ٿJ��-a�@�k�T4@�;Z.̐!?�����+�@�A3��ٿ�i�%Q@�@n7�?K4@�Y�Yp�!?1L�Qk��@�A3��ٿ�i�%Q@�@n7�?K4@�Y�Yp�!?1L�Qk��@�A3��ٿ�i�%Q@�@n7�?K4@�Y�Yp�!?1L�Qk��@�A3��ٿ�i�%Q@�@n7�?K4@�Y�Yp�!?1L�Qk��@�A3��ٿ�i�%Q@�@n7�?K4@�Y�Yp�!?1L�Qk��@�W(��ٿ9��-Zo�@���]�4@�}�sȐ!?�("���@���D��ٿ�MAC��@-��%4@���Ə�!?�� ����@���D��ٿ�MAC��@-��%4@���Ə�!?�� ����@>�j�ٿk�?zvk�@���� 4@<��:��!?y����@>�j�ٿk�?zvk�@���� 4@<��:��!?y����@���{�ٿ!��[�@�;���4@�NO;�!?5tN��@�.Lw�ٿ@�-��^�@����' 4@��~=�!??�96���@�q\�҈ٿ��
�1�@6��~�4@}�&8�!?�0��H�@�q\�҈ٿ��
�1�@6��~�4@}�&8�!?�0��H�@��;�Ŋٿ��q��@X�-��3@	�ֵm�!?{�#0l|�@��;�Ŋٿ��q��@X�-��3@	�ֵm�!?{�#0l|�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�?�a.�ٿ�)�h��@�&��� 4@�Z�A\�!?�?���S�@�p�Ǎٿ�� �@�4B�W 4@k��aw�!?x(���@�p�Ǎٿ�� �@�4B�W 4@k��aw�!?x(���@�p�Ǎٿ�� �@�4B�W 4@k��aw�!?x(���@�p�Ǎٿ�� �@�4B�W 4@k��aw�!?x(���@geʛ�ٿ|�|�p��@��Oy�4@�A����!?��?�q��@geʛ�ٿ|�|�p��@��Oy�4@�A����!?��?�q��@�>Ѹ��ٿ��V~P��@Q��4@/KpPE�!?����{��@##߃�ٿy:[�D��@0r��4@���J�!?�����@##߃�ٿy:[�D��@0r��4@���J�!?�����@##߃�ٿy:[�D��@0r��4@���J�!?�����@##߃�ٿy:[�D��@0r��4@���J�!?�����@�5���ٿ[�Mo��@�R^�44@�.$)��!?d�o�|h�@�5���ٿ[�Mo��@�R^�44@�.$)��!?d�o�|h�@�5���ٿ[�Mo��@�R^�44@�.$)��!?d�o�|h�@��Ћ�ٿ������@�XRv4@�%(Đ�!?iNɄ��@w���ٿY�7vb��@)]1}4@�GJ̐!?�3��@w���ٿY�7vb��@)]1}4@�GJ̐!?�3��@w���ٿY�7vb��@)]1}4@�GJ̐!?�3��@w���ٿY�7vb��@)]1}4@�GJ̐!?�3��@�^�yC�ٿ}��Jy�@����4@6�7��!?�}> ���@E5��b�ٿ�y���@�"WJ4@o�}G��!?c��(*=�@E5��b�ٿ�y���@�"WJ4@o�}G��!?c��(*=�@�K*�܈ٿ���a�@;�'7C4@o.T��!?U
��E3�@�K*�܈ٿ���a�@;�'7C4@o.T��!?U
��E3�@��9J�ٿ�h����@/���4@Q�q��!?�Q�Ae��@��9J�ٿ�h����@/���4@Q�q��!?�Q�Ae��@��9J�ٿ�h����@/���4@Q�q��!?�Q�Ae��@��@J�ٿZS=�;�@Y0�4@��p԰�!?N������@��@J�ٿZS=�;�@Y0�4@��p԰�!?N������@��@J�ٿZS=�;�@Y0�4@��p԰�!?N������@��@J�ٿZS=�;�@Y0�4@��p԰�!?N������@��@J�ٿZS=�;�@Y0�4@��p԰�!?N������@}mF,�ٿhN7k���@XJJ�4@z
���!?� �h��@R�{:�~ٿ�}7�Ċ�@��4@r��ܐ!?L�:�]�@R�{:�~ٿ�}7�Ċ�@��4@r��ܐ!?L�:�]�@R�{:�~ٿ�}7�Ċ�@��4@r��ܐ!?L�:�]�@R�{:�~ٿ�}7�Ċ�@��4@r��ܐ!?L�:�]�@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@-�ɤ{ٿ�[M�֨�@~�h��4@����ې!?)�Ń���@�F�q�ٿ �sM�0�@4���4@[�b�!?���nU�@\7JgۅٿL	�Ԭ��@�M���4@d��y�!?��6���@\7JgۅٿL	�Ԭ��@�M���4@d��y�!?��6���@\7JgۅٿL	�Ԭ��@�M���4@d��y�!?��6���@\7JgۅٿL	�Ԭ��@�M���4@d��y�!?��6���@\7JgۅٿL	�Ԭ��@�M���4@d��y�!?��6���@Z%鯅�ٿ���X��@40��4@1�%ȵ�!?�}(���@Z%鯅�ٿ���X��@40��4@1�%ȵ�!?�}(���@�����ٿ������@�ǜٳ4@����!?t)��JN�@�����ٿ������@�ǜٳ4@����!?t)��JN�@�V��ٿ�A����@��;��4@P뭁͐!?��3�@�V��ٿ�A����@��;��4@P뭁͐!?��3�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@����%ٿ<O���@Mk�#-4@�����!?rX��'�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�Y���ٿc��_��@b sg4@����R�!?����1�@�U�a��ٿ�O[�f�@'�gi.	4@Z:�{�!?L�wm^�@�Cp���ٿ���#��@�<��.4@�J\�!?9)mQj9�@z�
���ٿ@�l��@r���	4@�c繱�!?X$Qt|q�@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@x�)�/}ٿ�-,æ�@�,(4@��(��!?�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�:I�{ٿ��\«��@�T�4@� D��!?}�����@�A�p��ٿJh
��O�@�k�� 4@.+�pq�!?z�՟��@�A�p��ٿJh
��O�@�k�� 4@.+�pq�!?z�՟��@�A�p��ٿJh
��O�@�k�� 4@.+�pq�!?z�՟��@�A�p��ٿJh
��O�@�k�� 4@.+�pq�!?z�՟��@�A�p��ٿJh
��O�@�k�� 4@.+�pq�!?z�՟��@ߊǦ�ٿza_��@�"��-4@R7|#9�!?����O��@ߊǦ�ٿza_��@�"��-4@R7|#9�!?����O��@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@�wj�N�ٿ���Y�@�Nޡ� 4@�@�ِ!?��AB���@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@w����ٿ4[�h��@0' %E4@!�p��!?�����\�@����ٿV��]t�@B�P�4@��0��!?���R�>�@��E�ٿ��Id�@9�;~��3@v��א!?����ݜ�@7e�Foٿ̾���n�@�*��3@�� ���!?)@��� �@�A1�b�ٿL�|����@Y�<�4@9�	��!?m4����@�A1�b�ٿL�|����@Y�<�4@9�	��!?m4����@�A1�b�ٿL�|����@Y�<�4@9�	��!?m4����@�A1�b�ٿL�|����@Y�<�4@9�	��!?m4����@�A1�b�ٿL�|����@Y�<�4@9�	��!?m4����@�Z4�|ٿ���L~-�@8S�U=4@^��Ӑ!?���=@��@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@\����ٿ6�>��C�@E�W��4@���=�!?֍2�<�@e_`�ٿ��t���@�ggY4@��D��!?��mր+�@�w��c�ٿ�f)�a�@`|�!4@Rױ��!?�<�ن�@�w��c�ٿ�f)�a�@`|�!4@Rױ��!?�<�ن�@�w��c�ٿ�f)�a�@`|�!4@Rױ��!?�<�ن�@u���ٿt��2E��@R��O�4@�Ka���!?�32 0��@u���ٿt��2E��@R��O�4@�Ka���!?�32 0��@u���ٿt��2E��@R��O�4@�Ka���!?�32 0��@u���ٿt��2E��@R��O�4@�Ka���!?�32 0��@u���ٿt��2E��@R��O�4@�Ka���!?�32 0��@��56؅ٿ$�kL��@����a4@��?˼�!?�����f�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@qģ���ٿ`.����@h�k�4@�ǿ´�!?����W�@/��e}ٿ9����@�d��4@I�Y�Ɛ!?f�;�r�@/��e}ٿ9����@�d��4@I�Y�Ɛ!?f�;�r�@/��e}ٿ9����@�d��4@I�Y�Ɛ!?f�;�r�@/��e}ٿ9����@�d��4@I�Y�Ɛ!?f�;�r�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@�q��~ٿ��:���@j�ً�4@%z��!?�Պr�(�@j��㴀ٿ�NHE.�@�<��4@���ސ!?θ�	׆�@3'!M�}ٿ�}i�Z��@���lc4@�@���!?�����@3'!M�}ٿ�}i�Z��@���lc4@�@���!?�����@3'!M�}ٿ�}i�Z��@���lc4@�@���!?�����@˚oO{�ٿ
a-s���@�V34@��Q��!?�j#S*�@ݍP�ٿ�D̹���@+�6P4@�T/�!?�:�����@`��;�ٿ��%u���@���O\4@�O3�!?���ѫ��@`��;�ٿ��%u���@���O\4@�O3�!?���ѫ��@`��;�ٿ��%u���@���O\4@�O3�!?���ѫ��@`��;�ٿ��%u���@���O\4@�O3�!?���ѫ��@-��]e�ٿ���7���@��e��4@�iE�~�!?���J���@-��]e�ٿ���7���@��e��4@�iE�~�!?���J���@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@ǻC�:�ٿE�8e���@����	4@�C��D�!?���oId�@hT4D2�ٿM�+�j�@{#:�2
4@�aiN�!?���b'��@�щ�R�ٿu�\b���@���	4@,�<���!?c� .^m�@�щ�R�ٿu�\b���@���	4@,�<���!?c� .^m�@�щ�R�ٿu�\b���@���	4@,�<���!?c� .^m�@�щ�R�ٿu�\b���@���	4@,�<���!?c� .^m�@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@*�3/ىٿ���(?e�@`��4@�Ǵ1��!?����*��@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�;'8]~ٿ��Z=i}�@�ȃ�@4@����Ð!?\�����@�R��ٿcߢ�@׮�4@��(�!?�3����@���΃ٿ̷���@�@��4@�ȍK��!?��`H���@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@��@ �ٿThĥ��@����|4@Y�ܘ��!?��\�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@�y{ϊٿE�����@y:�4@W�2<l�!?����>�@(MN~ˊٿ�6E�@drd�g4@k�͐!?�
�p�@(MN~ˊٿ�6E�@drd�g4@k�͐!?�
�p�@(MN~ˊٿ�6E�@drd�g4@k�͐!?�
�p�@(MN~ˊٿ�6E�@drd�g4@k�͐!?�
�p�@(MN~ˊٿ�6E�@drd�g4@k�͐!?�
�p�@5�)�:�ٿ�'��W�@ūd2� 4@M��ΐ!?�
@t���@5�)�:�ٿ�'��W�@ūd2� 4@M��ΐ!?�
@t���@5�)�:�ٿ�'��W�@ūd2� 4@M��ΐ!?�
@t���@5�)�:�ٿ�'��W�@ūd2� 4@M��ΐ!?�
@t���@�����ٿ��Ǡ\�@�¾3�4@_�n�̐!?K'����@WnzD{ٿ��;��@���7�4@8]n*��!?�+�
]�@WnzD{ٿ��;��@���7�4@8]n*��!?�+�
]�@WnzD{ٿ��;��@���7�4@8]n*��!?�+�
]�@WnzD{ٿ��;��@���7�4@8]n*��!?�+�
]�@������ٿ�gK���@�b� 4@҇�~��!?���5�@������ٿ�gK���@�b� 4@҇�~��!?���5�@������ٿ�gK���@�b� 4@҇�~��!?���5�@������ٿ�gK���@�b� 4@҇�~��!?���5�@E���,�ٿ|`F��@�@/vB�4@�dӏɐ!?��#ӹ�@`hZ!�ٿ��+Y�d�@�T�"�4@�����!?ᬱ/5�@`hZ!�ٿ��+Y�d�@�T�"�4@�����!?ᬱ/5�@`hZ!�ٿ��+Y�d�@�T�"�4@�����!?ᬱ/5�@`hZ!�ٿ��+Y�d�@�T�"�4@�����!?ᬱ/5�@3��Rh�ٿY-q�5��@aZ��4@x�:���!?�:�m5�@3��Rh�ٿY-q�5��@aZ��4@x�:���!?�:�m5�@3��Rh�ٿY-q�5��@aZ��4@x�:���!?�:�m5�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@y@֣ �ٿ`&��H��@N����4@�/k��!?$!�ߚ�@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�n�XC�ٿq�\����@����4@kdb�!?��}��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�&ʊ�ٿ�5����@_#\�4@ؙ$���!?�e�c��@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@�x}H�ٿ&�E���@�ქ�4@�V�V�!?0����@$X��ٿdƌ}2�@���<v4@�-�ڐ!?�ˣ�0�@$X��ٿdƌ}2�@���<v4@�-�ڐ!?�ˣ�0�@$X��ٿdƌ}2�@���<v4@�-�ڐ!?�ˣ�0�@$X��ٿdƌ}2�@���<v4@�-�ڐ!?�ˣ�0�@"^�� �ٿ���Y�@?�LF4@���!?<��XA��@"^�� �ٿ���Y�@?�LF4@���!?<��XA��@"^�� �ٿ���Y�@?�LF4@���!?<��XA��@"^�� �ٿ���Y�@?�LF4@���!?<��XA��@��^�ٿd�n����@�b3�z4@9��3�!?�q��Do�@|�2��|ٿ�s�
���@b}�(4@~���.�!?��,���@|�2��|ٿ�s�
���@b}�(4@~���.�!?��,���@|�2��|ٿ�s�
���@b}�(4@~���.�!?��,���@|�2��|ٿ�s�
���@b}�(4@~���.�!?��,���@|�2��|ٿ�s�
���@b}�(4@~���.�!?��,���@
���ٿ�m�����@�w]��4@ 3>��!?J+�a�-�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@o�_ٿ��v.��@�+�m4@�]�-ܐ!?�V��<�@8vi/=�ٿjo=��@�w]	4@�[BKɐ!?!�i~<�@8vi/=�ٿjo=��@�w]	4@�[BKɐ!?!�i~<�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@`�;�Y�ٿ���	���@A�o�4@�x�얐!?�ٟ�6�@��;L�ٿֺ�a��@�AI
4@>_�>l�!?��	���@��;L�ٿֺ�a��@�AI
4@>_�>l�!?��	���@ � �ٿog+#��@L���4@)����!?f�!���@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@4��<�ٿ�;{���@�<�4@�{(w��!?u��9K�@��J	�ٿ,�����@��[)�4@=�)6��!?ϑӀ�`�@��7U�ٿ�yV�&��@S7:o4@��w�|�!?����!*�@��7U�ٿ�yV�&��@S7:o4@��w�|�!?����!*�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@�e���ٿX�x��0�@���4@r<Ƥ�!?s�P�r�@���s�ٿ	gw���@��� 4@�j>�!?R)�
���@���s�ٿ	gw���@��� 4@�j>�!?R)�
���@���s�ٿ	gw���@��� 4@�j>�!?R)�
���@���s�ٿ	gw���@��� 4@�j>�!?R)�
���@���s�ٿ	gw���@��� 4@�j>�!?R)�
���@#"��5�ٿ�����@<���4@��^��!?4pzk�@#"��5�ٿ�����@<���4@��^��!?4pzk�@#"��5�ٿ�����@<���4@��^��!?4pzk�@��;㤋ٿ!�#c2�@�#��4@:��Ʋ�!?@r��0�@��;㤋ٿ!�#c2�@�#��4@:��Ʋ�!?@r��0�@��;㤋ٿ!�#c2�@�#��4@:��Ʋ�!?@r��0�@��;㤋ٿ!�#c2�@�#��4@:��Ʋ�!?@r��0�@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@�$O�ׂٿ���C��@,���4@�����!?��`����@���M�ٿ��W�l�@�����4@p/ `��!?�����@���M�ٿ��W�l�@�����4@p/ `��!?�����@���M�ٿ��W�l�@�����4@p/ `��!?�����@���M�ٿ��W�l�@�����4@p/ `��!?�����@�@�V�ٿP)�@v��@���4@�6Qƿ�!?`�c*�L�@�@�V�ٿP)�@v��@���4@�6Qƿ�!?`�c*�L�@�T��ٿ�
S�?��@���w4@����̐!?�_����@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@j����ٿ�Q�2^��@���94@'Pk��!?�c�&��@\/���ٿ0�7�Z�@�a���4@��7��!?�+Ad���@X�?6)�ٿ/.��@���l4@y�DҐ!?_��˘<�@X�?6)�ٿ/.��@���l4@y�DҐ!?_��˘<�@uqN1��ٿQ�l|�@c��{�4@����ڐ!?�l ��h�@�����ٿ�����@�@5���j4@`��̐!?�����@�����ٿ�����@�@5���j4@`��̐!?�����@�z4-q�ٿC82��@"��4@�P�3��!?��I���@�z4-q�ٿC82��@"��4@�P�3��!?��I���@�z4-q�ٿC82��@"��4@�P�3��!?��I���@�z4-q�ٿC82��@"��4@�P�3��!?��I���@3�����ٿ&��[�F�@�z��4@�ckM�!?�mYe��@���I��ٿ1����@���Z`4@b�A�!?Zan�L`�@���I��ٿ1����@���Z`4@b�A�!?Zan�L`�@���I��ٿ1����@���Z`4@b�A�!?Zan�L`�@���&�ٿ��R��>�@s��l 4@_
0{T�!?͵v[�+�@���&�ٿ��R��>�@s��l 4@_
0{T�!?͵v[�+�@�v��]�ٿV�~{���@�zRHP4@VJ*n�!?�}Pý�@�v��]�ٿV�~{���@�zRHP4@VJ*n�!?�}Pý�@�v��]�ٿV�~{���@�zRHP4@VJ*n�!?�}Pý�@�v��]�ٿV�~{���@�zRHP4@VJ*n�!?�}Pý�@�v��]�ٿV�~{���@�zRHP4@VJ*n�!?�}Pý�@g����ٿa��J��@���'4@73�
�!?�+�!���@P�h~�ٿ�eL��=�@C��}4@�pf�,�!?�i����@P�h~�ٿ�eL��=�@C��}4@�pf�,�!?�i����@P�h~�ٿ�eL��=�@C��}4@�pf�,�!?�i����@P�h~�ٿ�eL��=�@C��}4@�pf�,�!?�i����@P�h~�ٿ�eL��=�@C��}4@�pf�,�!?�i����@����8ٿ<��9�@�O�.�4@}z�ِ!?t/1����@s�_�ٿL/�)��@"#9�"4@֤��t�!?jv'�+��@s�_�ٿL/�)��@"#9�"4@֤��t�!?jv'�+��@|���ٿ/+�*���@�K��� 4@�
�댐!?憎��F�@Dl�O~ٿL�v���@h�$4@.T7C��!?�m���@Dl�O~ٿL�v���@h�$4@.T7C��!?�m���@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�vrh�ٿ��G�@�|�� 4@��M���!?pWdm�+�@�$�!��ٿ3���E�@?�W
4@|N¨�!?��atg��@�$�!��ٿ3���E�@?�W
4@|N¨�!?��atg��@�g/K-�ٿ�O �׃�@�:k˜�3@ �tX�!?�;ST��@�g/K-�ٿ�O �׃�@�:k˜�3@ �tX�!?�;ST��@��)H܈ٿ�jb��`�@��-�N�3@(�X���!?�B�%���@��)H܈ٿ�jb��`�@��-�N�3@(�X���!?�B�%���@��)H܈ٿ�jb��`�@��-�N�3@(�X���!?�B�%���@��)H܈ٿ�jb��`�@��-�N�3@(�X���!?�B�%���@iඍ�ٿ��ZK1�@��k�4@(�Á��!?�c"m�7�@iඍ�ٿ��ZK1�@��k�4@(�Á��!?�c"m�7�@iඍ�ٿ��ZK1�@��k�4@(�Á��!?�c"m�7�@�Yи�ٿq�ԙ���@PC]w�4@i�Λ�!?1K�t�@(0KW<�ٿ����@�Ὁ4@w��Ӑ!?�g���@(0KW<�ٿ����@�Ὁ4@w��Ӑ!?�g���@(0KW<�ٿ����@�Ὁ4@w��Ӑ!?�g���@(0KW<�ٿ����@�Ὁ4@w��Ӑ!?�g���@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@���ٿ��(�@h�\{4@:�PT��!?��]�K��@:m�8�ٿ<�y!���@j|�"4@}��R�!?��M���@:m�8�ٿ<�y!���@j|�"4@}��R�!?��M���@:m�8�ٿ<�y!���@j|�"4@}��R�!?��M���@�+\a�ٿ�6A~�@\��4@���p�!?HJ���a�@���8x�ٿYGN��l�@t��4@�Y���!?�Cg
b�@���8x�ٿYGN��l�@t��4@�Y���!?�Cg
b�@���8x�ٿYGN��l�@t��4@�Y���!?�Cg
b�@{�w���ٿ������@^0�54@�3Xҍ�!?]Q��J�@{�w���ٿ������@^0�54@�3Xҍ�!?]Q��J�@{�w���ٿ������@^0�54@�3Xҍ�!?]Q��J�@{�w���ٿ������@^0�54@�3Xҍ�!?]Q��J�@a^0�d�ٿZ?��@ď[4<4@7�*dt�!?� lZ@�@a^0�d�ٿZ?��@ď[4<4@7�*dt�!?� lZ@�@a^0�d�ٿZ?��@ď[4<4@7�*dt�!?� lZ@�@a^0�d�ٿZ?��@ď[4<4@7�*dt�!?� lZ@�@E�hC��ٿ�r���@a&���4@n�����!?P�*�%�@E�hC��ٿ�r���@a&���4@n�����!?P�*�%�@E�hC��ٿ�r���@a&���4@n�����!?P�*�%�@E�hC��ٿ�r���@a&���4@n�����!?P�*�%�@cw8σٿ�7N
��@�xOE 4@���ې!?�~{k��@cw8σٿ�7N
��@�xOE 4@���ې!?�~{k��@�v.�ٿ �X3�"�@�����4@�\�!?����@B�y�zٿ�x����@�{Q���3@b�`��!?ZhrL=��@B�y�zٿ�x����@�{Q���3@b�`��!?ZhrL=��@B�y�zٿ�x����@�{Q���3@b�`��!?ZhrL=��@�o�#a{ٿc?��j�@���4@f���ΐ!?�����@�o�#a{ٿc?��j�@���4@f���ΐ!?�����@NZ�Ls�ٿ�q*PK�@V��.	4@�`s�ِ!?�ZN���@NZ�Ls�ٿ�q*PK�@V��.	4@�`s�ِ!?�ZN���@NZ�Ls�ٿ�q*PK�@V��.	4@�`s�ِ!?�ZN���@NZ�Ls�ٿ�q*PK�@V��.	4@�`s�ِ!?�ZN���@NZ�Ls�ٿ�q*PK�@V��.	4@�`s�ِ!?�ZN���@E��xČٿ,����@����z4@��J�!?��0C7�@�_�O�ٿ��!7���@�AcS�4@F�yp�!?�>��	�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@E�=Gx�ٿ/t��^�@��L�R	4@���u��!?J ݚ�@1���k}ٿdm��j��@���+4@�?��̐!??ֳ���@�VN�5yٿG��\r@�@ȋ쵫4@4�i4�!?�a��/��@�VN�5yٿG��\r@�@ȋ쵫4@4�i4�!?�a��/��@�VN�5yٿG��\r@�@ȋ쵫4@4�i4�!?�a��/��@�VN�5yٿG��\r@�@ȋ쵫4@4�i4�!?�a��/��@ȹp�lzٿbe/����@2+�?��3@�o� �!?цǇT��@ȹp�lzٿbe/����@2+�?��3@�o� �!?цǇT��@��`�yٿ�F��@�H���3@ަQǐ!?���*;�@��`�yٿ�F��@�H���3@ަQǐ!?���*;�@� ���ٿ}��~M��@����3@�MG/��!?�vn���@� ���ٿ}��~M��@����3@�MG/��!?�vn���@��V��ٿ+���*�@��� 4@b�U���!?���ԝ.�@��V��ٿ+���*�@��� 4@b�U���!?���ԝ.�@Pg��ٿ�v�I�@Y;�"�3@���K�!?�;	�7�@Pg��ٿ�v�I�@Y;�"�3@���K�!?�;	�7�@�>���ٿ��s��@m�@� 4@��^6I�!?�v[_o�@��\�ˇٿ"����@���~4@0�:Y�!?����@��\�ˇٿ"����@���~4@0�:Y�!?����@�@���ٿkcd���@{��3|4@"QD�T�!?}��
 ��@�@���ٿkcd���@{��3|4@"QD�T�!?}��
 ��@�Y }ٿ0�w��@;�R�M4@��g��!?��q����@Ow���ٿ�D�h��@��4@A "�D�!?�㏵�q�@Ow���ٿ�D�h��@��4@A "�D�!?�㏵�q�@��3�f�ٿ��y�0h�@V�6� 4@p��֐!?H�e��@��3�f�ٿ��y�0h�@V�6� 4@p��֐!?H�e��@��3�f�ٿ��y�0h�@V�6� 4@p��֐!?H�e��@��3�f�ٿ��y�0h�@V�6� 4@p��֐!?H�e��@l�jw��ٿ�B�~G�@*F�"4@	�E��!?v%O��@l�jw��ٿ�B�~G�@*F�"4@	�E��!?v%O��@l�jw��ٿ�B�~G�@*F�"4@	�E��!?v%O��@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@?���ٿ���o��@���z�4@j�N1ϐ!?.�t$`�@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�`�ÚٿG���n�@����4@H4�
�!?��Ɗ{��@�!e3�~ٿ��1cF��@�wt?�4@����!?�W)��@�@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@��9�ٿJ�VǺ�@��}4@�ఁ�!?��Ѣ1��@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@a �}��ٿ�[ ��@�5>�I4@�|��!?	T��p�@B�Ӣ\�ٿM� Ӥ��@U�N,	4@���d��!?Y��(t��@B�Ӣ\�ٿM� Ӥ��@U�N,	4@���d��!?Y��(t��@B�Ӣ\�ٿM� Ӥ��@U�N,	4@���d��!?Y��(t��@f��"��ٿ
�Ӷ,��@Û���4@���P�!?�b���@f��"��ٿ
�Ӷ,��@Û���4@���P�!?�b���@f��"��ٿ
�Ӷ,��@Û���4@���P�!?�b���@f��"��ٿ
�Ӷ,��@Û���4@���P�!?�b���@�	���ٿV㙅���@�L����3@�`p`Ր!?���ֻ��@��*��ٿ��}��@Y6F��3@C����!?М�V��@��*��ٿ��}��@Y6F��3@C����!?М�V��@��*��ٿ��}��@Y6F��3@C����!?М�V��@��*��ٿ��}��@Y6F��3@C����!?М�V��@��*��ٿ��}��@Y6F��3@C����!?М�V��@ոN��ٿ:lS��1�@T�A}	�3@طer��!?ݘ�o��@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@y��6ٿi�V.>��@�cs�4@Ø���!?���W�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�k����ٿ�C�x��@��	'4@�q5���!?WL�Q�@�����ٿ`�7�l)�@�GD4@s���!?��\Q�@�����ٿ`�7�l)�@�GD4@s���!?��\Q�@�����ٿ`�7�l)�@�GD4@s���!?��\Q�@�����ٿ`�7�l)�@�GD4@s���!?��\Q�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@�
�Q`�ٿBy�u���@�=�%4@����!?��U�1�@P��'�ٿ�	�����@�pKS4@��C���!?+��*eR�@P��'�ٿ�	�����@�pKS4@��C���!?+��*eR�@P��'�ٿ�	�����@�pKS4@��C���!?+��*eR�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@`�T	ϋٿ	<W��@�l��04@@b���!?F�JKg�@�0�ٿ��mfK�@�(��44@��62��!?ͻAGK�@�0�ٿ��mfK�@�(��44@��62��!?ͻAGK�@�0�ٿ��mfK�@�(��44@��62��!?ͻAGK�@�0�ٿ��mfK�@�(��44@��62��!?ͻAGK�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@#����ٿnS��2��@��	�4@���6��!?>>T�M�@>nv�ٿ���m)x�@�Ι��4@z��ҥ�!?�.)�L�@>nv�ٿ���m)x�@�Ι��4@z��ҥ�!?�.)�L�@>nv�ٿ���m)x�@�Ι��4@z��ҥ�!?�.)�L�@>nv�ٿ���m)x�@�Ι��4@z��ҥ�!?�.)�L�@>nv�ٿ���m)x�@�Ι��4@z��ҥ�!?�.)�L�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@N���ʈٿ��u;��@��"4@��;�Ȑ!?p=H��6�@Y�}|�ٿ	�����@�
��6	4@B���!?d�Z� ��@zq�ٿ�@�a��@m0�)
4@Ky�c��!?:t~�m�@zq�ٿ�@�a��@m0�)
4@Ky�c��!?:t~�m�@zq�ٿ�@�a��@m0�)
4@Ky�c��!?:t~�m�@zq�ٿ�@�a��@m0�)
4@Ky�c��!?:t~�m�@zq�ٿ�@�a��@m0�)
4@Ky�c��!?:t~�m�@B"אɂٿ�}xMɫ�@*ɻ{4@RU}���!?^�:��m�@B"אɂٿ�}xMɫ�@*ɻ{4@RU}���!?^�:��m�@+�arރٿ�����@>���4@]��!?�Z`�em�@+�arރٿ�����@>���4@]��!?�Z`�em�@+�arރٿ�����@>���4@]��!?�Z`�em�@�0(��ٿ�E����@���P4@� i ː!?W�T��@�0(��ٿ�E����@���P4@� i ː!?W�T��@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@�rx/��ٿ%��Q�@�;S��4@m�0b��!?��$I���@b/� %�ٿ�"9/T�@�R���4@����!?Q�����@e��T�ٿ4�r��@���f	4@V���!?oS#ߌ!�@�����ٿ�^O���@���k4@��h��!?����e��@vJ6���ٿ��y���@8vK�4@��3��!?��|q��@vJ6���ٿ��y���@8vK�4@��3��!?��|q��@vJ6���ٿ��y���@8vK�4@��3��!?��|q��@77f��ٿ9�����@���l�4@���X�!?̽6�_�@#0���ٿ�-?��@s�s�Z4@v8U�B�!?����Z�@�O΁ٿFBp$��@9I�R4@�6�k�!?9��M߻�@����~ٿ���=�J�@w��4A4@�k�ܐ!?@�[MLd�@����~ٿ���=�J�@w��4A4@�k�ܐ!?@�[MLd�@����~ٿ���=�J�@w��4A4@�k�ܐ!?@�[MLd�@����~ٿ���=�J�@w��4A4@�k�ܐ!?@�[MLd�@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@KA8d�|ٿշ=P&-�@P�,q4@�蟪�!?��Ԃ��@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@C�0�uٿ�\�ȓ�@5�0a�4@�-bf�!?�U~���@�^2�ٿ�9����@H�7�k4@.0[���!?-��o�]�@lD4�~�ٿ$EZH��@���	Q4@�]�V�!?�ӹRi#�@lD4�~�ٿ$EZH��@���	Q4@�]�V�!?�ӹRi#�@_�fǴ~ٿ�-�����@��>�R4@$�}�\�!?�����@2C�T�ٿD	���4�@cj���
4@=Bg��!?��$�@��@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@��	ʈٿK|1E �@��Ą�4@��Ԥ��!?�(�+�C�@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@���G�ٿ�4 ��@�v���4@V9y���!?Q+���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@}_�^ӈٿ��7�!�@��"!l4@'�lӐ!?�p(j���@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�+��:�ٿ5��b��@-o�Je4@�w����!?Lś�4�@�<�#�ٿ�ǥ���@�Y��4@��ggϐ!?��8	�@�<�#�ٿ�ǥ���@�Y��4@��ggϐ!?��8	�@�<�#�ٿ�ǥ���@�Y��4@��ggϐ!?��8	�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�玄�ٿ��<�&�@��H�4@�,���!?Y{P?m�@�B(p�ٿO ��@��U*�	4@֡�А!?F�Y2��@�B(p�ٿO ��@��U*�	4@֡�А!?F�Y2��@�B(p�ٿO ��@��U*�	4@֡�А!?F�Y2��@�B(p�ٿO ��@��U*�	4@֡�А!?F�Y2��@���O�|ٿ �բ��@�v�L4@t@�`��!?�P9��@���O�|ٿ �բ��@�v�L4@t@�`��!?�P9��@���O�|ٿ �բ��@�v�L4@t@�`��!?�P9��@���O�|ٿ �բ��@�v�L4@t@�`��!?�P9��@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�.�{zٿ��p�V(�@�`��4@��%���!?����Q+�@�eb�ކٿoYN �x�@���H�3@���#��!?�mݼ���@���ٿ�;�Q�h�@	���4@�����!?����@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@��a�ٿ�c~��@ֳ��4@�����!?��3Ƿ��@㋣��ٿ�؂�P��@����M4@uQ���!?%�5���@㋣��ٿ�؂�P��@����M4@uQ���!?%�5���@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@AA�\ٿҚWo�-�@��Q,�4@����ɐ!?PlA��G�@�A�5�ٿ"�(�[!�@<bd4@�L�ސ!?̦�H>��@�A�5�ٿ"�(�[!�@<bd4@�L�ސ!?̦�H>��@�A�5�ٿ"�(�[!�@<bd4@�L�ސ!?̦�H>��@�A�5�ٿ"�(�[!�@<bd4@�L�ސ!?̦�H>��@�A�5�ٿ"�(�[!�@<bd4@�L�ސ!?̦�H>��@�{�g��ٿC����0�@��Q�|4@��v��!?��*���@�{�g��ٿC����0�@��Q�|4@��v��!?��*���@�{�g��ٿC����0�@��Q�|4@��v��!?��*���@�{�g��ٿC����0�@��Q�|4@��v��!?��*���@�{�g��ٿC����0�@��Q�|4@��v��!?��*���@����̉ٿ1l���@����T4@x!�Đ!?�u����@����̉ٿ1l���@����T4@x!�Đ!?�u����@����̉ٿ1l���@����T4@x!�Đ!?�u����@A�+�j�ٿhm����@��x�4@`����!?��|@~��@�鯜��ٿu��(�@�k��4@O�y�!?��S;�U�@�鯜��ٿu��(�@�k��4@O�y�!?��S;�U�@�鯜��ٿu��(�@�k��4@O�y�!?��S;�U�@��~h�ٿn@|2f;�@8Y:�4@�����!?dl9���@��~h�ٿn@|2f;�@8Y:�4@�����!?dl9���@�Ƨq�ٿd��Х��@"�u1�4@����!?�s����@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���6�ٿ]%�L)��@�����4@��ש��!?���}��@���&!�ٿ��A���@9��E4@�,`�Ȑ!?�R�i��@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@z�)^�ٿ}c��@��	K4@���@ΐ!?A�>F�%�@%8×W�ٿ��qo}�@9��4@c����!?Vb����@%8×W�ٿ��qo}�@9��4@c����!?Vb����@%8×W�ٿ��qo}�@9��4@c����!?Vb����@��Lǃٿ�%�w���@��*��	4@�3��Ӑ!?�'��h�@�g �ٿ��I]N�@����o	4@�?|�!?��W��@�g �ٿ��I]N�@����o	4@�?|�!?��W��@Q,іw�ٿ�=+�`�@�09g�	4@0��o��!?�围��@Q,іw�ٿ�=+�`�@�09g�	4@0��o��!?�围��@Q,іw�ٿ�=+�`�@�09g�	4@0��o��!?�围��@Q,іw�ٿ�=+�`�@�09g�	4@0��o��!?�围��@]'� 8�ٿt~�[��@���4�4@��iѐ!?J�A��@���;�ٿ�VfG�@b�wP�4@��D	�!?�v����@���;�ٿ�VfG�@b�wP�4@��D	�!?�v����@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@㦏ˤ}ٿ덫6s��@G{��
4@/l'��!??�cv-�@F�����ٿj������@,�C�4@���͒�!?@�|7�v�@F�����ٿj������@,�C�4@���͒�!?@�|7�v�@F�����ٿj������@,�C�4@���͒�!?@�|7�v�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@(󾫂ٿ��A���@at�i4@���@ �!?x�Wx H�@�FPnȅٿ�,�]�@vp�UO4@[]У�!?�%Ζ��@�FPnȅٿ�,�]�@vp�UO4@[]У�!?�%Ζ��@�FPnȅٿ�,�]�@vp�UO4@[]У�!?�%Ζ��@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@	RG9�ٿ�GxT�@0=sC4@��$hϐ!?FW�����@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@�Y�R�ٿ��.M�N�@��o�4@a���!?;��m+o�@��+�ٿp������@���GB4@J�""�!?�r�AQ�@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�Kki�ٿ� ,��@��=�64@Q�V��!?G����@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@�UC��ٿn��TZ�@V� S4@�iob��!?�0�ۋ��@C�ʇٿ�RAa�f�@myZ:�4@8����!?3�%����@C�ʇٿ�RAa�f�@myZ:�4@8����!?3�%����@C�ʇٿ�RAa�f�@myZ:�4@8����!?3�%����@��Di��ٿ�^r��@���
 4@Sh��!?b�5��@��Di��ٿ�^r��@���
 4@Sh��!?b�5��@��Di��ٿ�^r��@���
 4@Sh��!?b�5��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@��u��ٿ�l��ȓ�@E!4@_v�dΐ!?���P��@Ϳ�0V�ٿyXQϷ�@Ph7�k4@�3�+��!?�H�fM��@Oe��T�ٿ�@�h�@���4@����!?05�ú�@Oe��T�ٿ�@�h�@���4@����!?05�ú�@Oe��T�ٿ�@�h�@���4@����!?05�ú�@��v�ٿq����H�@�M�J4@Y�@�!?��T�dD�@��v�ٿq����H�@�M�J4@Y�@�!?��T�dD�@��v�ٿq����H�@�M�J4@Y�@�!?��T�dD�@��v�ٿq����H�@�M�J4@Y�@�!?��T�dD�@��v�ٿq����H�@�M�J4@Y�@�!?��T�dD�@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@�M-5�ٿZ���˽�@�����4@&*DNې!?�!-N���@���LԀٿW+ig�Y�@�)݌4@���:�!?�F�W���@���LԀٿW+ig�Y�@�)݌4@���:�!?�F�W���@���LԀٿW+ig�Y�@�)݌4@���:�!?�F�W���@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@[���ٿ�6���@'�oA4@]	ߚ�!?�fY�c��@��5�ٿ@�\P��@���K�4@g���!?��6�,�@��5�ٿ@�\P��@���K�4@g���!?��6�,�@��5�ٿ@�\P��@���K�4@g���!?��6�,�@��5�ٿ@�\P��@���K�4@g���!?��6�,�@��5�ٿ@�\P��@���K�4@g���!?��6�,�@�]{�+�ٿ����@����A4@�E��!?�D�.��@�]{�+�ٿ����@����A4@�E��!?�D�.��@�]{�+�ٿ����@����A4@�E��!?�D�.��@�]{�+�ٿ����@����A4@�E��!?�D�.��@��ߛg�ٿ�ͣ�gB�@J���3@e].��!?p�)��@	\�}ٿB�J4���@���y4@����!?��#�2��@�X0M�ٿ�'��5�@~s�/4@#�����!?���@�@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@��r/R�ٿ$�{[���@Q	���3@��N��!?���P=��@"�Cd�ٿQ�@����@7�p��3@Ң �k�!?�d�oɼ�@"�Cd�ٿQ�@����@7�p��3@Ң �k�!?�d�oɼ�@"�Cd�ٿQ�@����@7�p��3@Ң �k�!?�d�oɼ�@"�Cd�ٿQ�@����@7�p��3@Ң �k�!?�d�oɼ�@"�Cd�ٿQ�@����@7�p��3@Ң �k�!?�d�oɼ�@�A�ӆٿN�/p
�@��2�� 4@��l̫�!?�\��8�@�A�ӆٿN�/p
�@��2�� 4@��l̫�!?�\��8�@�A�ӆٿN�/p
�@��2�� 4@��l̫�!?�\��8�@�A�ӆٿN�/p
�@��2�� 4@��l̫�!?�\��8�@E��#��ٿ{U�p���@��k�g4@Z�r���!?4&;�p�@���ٿ��̓�;�@��YU� 4@>]Z���!?�~�k���@���ٿ��̓�;�@��YU� 4@>]Z���!?�~�k���@���ٿ��̓�;�@��YU� 4@>]Z���!?�~�k���@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@9quj��ٿ�8.ͺ%�@x�[-+4@�w���!?{��Z��@X߯e��ٿ��[�#�@�аU�4@1� ��!??��<�@X߯e��ٿ��[�#�@�аU�4@1� ��!??��<�@X߯e��ٿ��[�#�@�аU�4@1� ��!??��<�@X߯e��ٿ��[�#�@�аU�4@1� ��!??��<�@X߯e��ٿ��[�#�@�аU�4@1� ��!??��<�@K{l1�ٿ �h���@���*�4@�B�\ɐ!?��&Pp��@�SЙ�ٿ8��kP�@���4@2;�t�!?i�?.�6�@ �t�ٿ�^�o��@	Z�Z4@�Q<֐!?�)+��|�@ �t�ٿ�^�o��@	Z�Z4@�Q<֐!?�)+��|�@�1>��ٿؓ�`��@��� 4@�d���!?mTb��@�1>��ٿؓ�`��@��� 4@�d���!?mTb��@�1>��ٿؓ�`��@��� 4@�d���!?mTb��@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@%O��C�ٿ�a�-���@���h�4@�e�嵐!?�h�o7�@�':�ٿ�4l�}��@�;�e4@μ��֐!?t\'pu<�@I�t��ٿ$@Rp�M�@[ϻ�4@[ű�͐!?~���@I�t��ٿ$@Rp�M�@[ϻ�4@[ű�͐!?~���@�����ٿi���@P Yڗ4@k�K��!?�|�I1�@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@�q�c~�ٿ�R_�� �@��]k4@�#N���!?�jQ�3��@>���ٿ��E �@�]G4@���6n�!?���=~�@>���ٿ��E �@�]G4@���6n�!?���=~�@>���ٿ��E �@�]G4@���6n�!?���=~�@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@c(���~ٿe�4]���@r�-�o4@Cߝ+x�!?|�vD��@�-��ٿ��<�_�@W��84@��v�s�!?������@�-��ٿ��<�_�@W��84@��v�s�!?������@�-��ٿ��<�_�@W��84@��v�s�!?������@�-��ٿ��<�_�@W��84@��v�s�!?������@s�R�{�ٿ[�8<�@i%�4@�
�Ӽ�!?�~j���@s�R�{�ٿ[�8<�@i%�4@�
�Ӽ�!?�~j���@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@>���s�ٿ�]�H�@D��4@6�.�ؐ!?�\ 
�;�@�� �y�ٿ��u�{	�@H�p��4@���א!?���.K��@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@o�,>��ٿ�M�p��@?yC4@����Ӑ!?k����@�iyU��ٿ+�w�'��@tJ�164@X<��"�!??z7�@�iyU��ٿ+�w�'��@tJ�164@X<��"�!??z7�@�iyU��ٿ+�w�'��@tJ�164@X<��"�!??z7�@�_�T\�ٿ;9h��@>�|� 4@k�8�!?*��~��@�_�T\�ٿ;9h��@>�|� 4@k�8�!?*��~��@�_�T\�ٿ;9h��@>�|� 4@k�8�!?*��~��@�_�T\�ٿ;9h��@>�|� 4@k�8�!?*��~��@�_�T\�ٿ;9h��@>�|� 4@k�8�!?*��~��@�[��8�ٿN[�� ��@6�,�4@[y�y�!?�k�O��@�[��8�ٿN[�� ��@6�,�4@[y�y�!?�k�O��@�[��8�ٿN[�� ��@6�,�4@[y�y�!?�k�O��@�[��8�ٿN[�� ��@6�,�4@[y�y�!?�k�O��@�[��8�ٿN[�� ��@6�,�4@[y�y�!?�k�O��@�~xt�ٿ��llV�@�L�4@�b�e�!?1R/<*J�@2V���ٿ��ڨ���@�\�x�4@��!?��o+Ҧ�@2V���ٿ��ڨ���@�\�x�4@��!?��o+Ҧ�@2V���ٿ��ڨ���@�\�x�4@��!?��o+Ҧ�@2V���ٿ��ڨ���@�\�x�4@��!?��o+Ҧ�@���#M�ٿ����@�5�K4@���.��!?�4'�߇�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@U�ޮ#ٿ�P�4��@��[�4@z,�=�!?�)�5;0�@��_Yyٿ⫉���@m� 4@�b�!? �Ewp%�@��_Yyٿ⫉���@m� 4@�b�!? �Ewp%�@!Щ�szٿ�`�Pѵ�@�j��'4@.HG��!?B�����@!Щ�szٿ�`�Pѵ�@�j��'4@.HG��!?B�����@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@U��+ׂٿD���wQ�@.A|ւ4@�'hݐ!?��)q��@%�����ٿ�`�m��@���2�
4@�^)��!?`#j��@%�����ٿ�`�m��@���2�
4@�^)��!?`#j��@%�����ٿ�`�m��@���2�
4@�^)��!?`#j��@%�����ٿ�`�m��@���2�
4@�^)��!?`#j��@%�����ٿ�`�m��@���2�
4@�^)��!?`#j��@�/��ٿ�gv�@o�RV	4@0Oop�!?�zmts�@�/��ٿ�gv�@o�RV	4@0Oop�!?�zmts�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@�X����ٿ��vƙg�@�w��7	4@y��'�!?`y��b�@��lq�ٿ���|�!�@F���S4@���C�!?���<��@�{��6�ٿQ=��@�2�Yb4@v��A�!?�e�^��@�{��6�ٿQ=��@�2�Yb4@v��A�!?�e�^��@�{��6�ٿQ=��@�2�Yb4@v��A�!?�e�^��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@o,�g͇ٿ3�1[pg�@��L�4@�L��!?9�	>��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@^P��w�ٿY�Eq���@l}�Y�4@�BN�!?}q*#��@X�F�׉ٿSw��~s�@,��	4@V�D��!?T[@R��@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@���ߙٿ�����@.洵��3@pz�2[�!?2���+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@�*әٿʾȕ���@bW&h��3@eda+�!?���v�+�@��e>��ٿ;����@{��U��3@!t�G�!?N|�w�+�@��e>��ٿ;����@{��U��3@!t�G�!?N|�w�+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@����ٿ��u���@��"���3@��|��!?�+���+�@7=t؛�ٿ��t���@�g��3@�3�xF�!?�c;�+�@7=t؛�ٿ��t���@�g��3@�3�xF�!?�c;�+�@ ̷Aʙٿ`
�w���@󡢐��3@{�'?�!?-�y��+�@ ̷Aʙٿ`
�w���@󡢐��3@{�'?�!?-�y��+�@B}���ٿ)_�]���@�-�|��3@~k�:�!?�!S��+�@�����ٿ�K�O���@�5H���3@a4�m�!?�����+�@� &ʙٿ�5,q���@�����3@��S��!?<����+�@� &ʙٿ�5,q���@�����3@��S��!?<����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@��H���ٿ*7����@�mݺ��3@%^�ʱ�!?�����+�@�a����ٿ��Y����@h �$��3@��uƐ!?��u��+�@�a����ٿ��Y����@h �$��3@��uƐ!?��u��+�@p/Ƿ�ٿ/3y���@5���3@<g����!?�:<��+�@p/Ƿ�ٿ/3y���@5���3@<g����!?�:<��+�@p/Ƿ�ٿ/3y���@5���3@<g����!?�:<��+�@p/Ƿ�ٿ/3y���@5���3@<g����!?�:<��+�@.68ęٿ&����@�V?/��3@?	���!?M�ź�+�@.68ęٿ&����@�V?/��3@?	���!?M�ź�+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@��Dٿ}�����@C p]��3@�;+1��!?Ő���+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@���M��ٿ-�L����@�N���3@&��K�!?lsV��+�@.�v��ٿ�z
����@��I���3@��>#�!?�Σ��+�@����ٿ�������@0fR��3@.F��!?O�\��+�@����ٿ�������@0fR��3@.F��!?O�\��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�l����ٿ�&�����@�5���3@�EK��!?� ��+�@�+o䭙ٿ�}�����@$���3@�Y5�!?E���+�@&$C��ٿV�j����@������3@�?{㨐!?G�f��+�@&$C��ٿV�j����@������3@�?{㨐!?G�f��+�@&$C��ٿV�j����@������3@�?{㨐!?G�f��+�@�|�%��ٿ������@3����3@R����!?t�q��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@wwc���ٿ��R����@n�Z���3@Ӓ*Ӑ!?Q�I��+�@���ú�ٿ��F����@̪�>��3@:�)��!?mly��+�@���ú�ٿ��F����@̪�>��3@:�)��!?mly��+�@���ú�ٿ��F����@̪�>��3@:�)��!?mly��+�@���ú�ٿ��F����@̪�>��3@:�)��!?mly��+�@��N���ٿ�yƜ���@)���3@�sT��!?�^��+�@��s���ٿ_�ʛ���@�ս���3@�	vr��!?x�̬�+�@�"�Ϧ�ٿ������@�/f���3@xCf��!?�?���+�@�"�Ϧ�ٿ������@�/f���3@xCf��!?�?���+�@�"�Ϧ�ٿ������@�/f���3@xCf��!?�?���+�@�;ۄ��ٿJ@����@
;>k��3@t��a�!?^H���+�@�;ۄ��ٿJ@����@
;>k��3@t��a�!?^H���+�@�;ۄ��ٿJ@����@
;>k��3@t��a�!?^H���+�@����ٿ�x�����@��9���3@�����!?�_��+�@�D��ٿ�
����@r����3@�|��!?.�0��+�@�D��ٿ�
����@r����3@�|��!?.�0��+�@6��+��ٿ��t����@֝v���3@�O��ː!?c��+�@6��+��ٿ��t����@֝v���3@�O��ː!?c��+�@rH��ٿ�h����@�����3@���"�!?c���+�@��䨙ٿ�������@���^��3@_��6�!?�;v��+�@K>�y��ٿ������@�+���3@&O��!?�~��+�@�nN+��ٿXZ#����@:��c��3@���!?�դ�+�@�nN+��ٿXZ#����@:��c��3@���!?�դ�+�@L�qç�ٿv�̳���@p���3@�>�<��!?��+�@hk���ٿ�[M����@+��3@�Co�!?OLe��+�@�i����ٿ����@�3���3@�U���!?��e��+�@�i����ٿ����@�3���3@�U���!?��e��+�@�㹙ٿ�������@�Rr���3@#�Vl��!?���+�@��ZN��ٿaw�����@�K����3@��~���!?J��+�@K
���ٿp�����@������3@Ըְ�!?�4���+�@K
���ٿp�����@������3@Ըְ�!?�4���+�@K
���ٿp�����@������3@Ըְ�!?�4���+�@K
���ٿp�����@������3@Ըְ�!?�4���+�@ ��t��ٿE������@�����3@�+ͷz�!?	���+�@ ��t��ٿE������@�����3@�+ͷz�!?	���+�@h��f��ٿE	�����@E(O��3@�+���!?k;��+�@��@ ��ٿ�J����@��j��3@�[���!?	E��+�@򯲙ٿE������@?�5I��3@��gF��!?�pK��+�@򯲙ٿE������@?�5I��3@��gF��!?�pK��+�@�1�S��ٿ��Ҩ���@Rl#9��3@01b/Ð!?]�.��+�@]����ٿ������@{H�l��3@� ٧��!?�=ͫ�+�@c�.��ٿ�����@�_x���3@�ۻ#�!?J�1��+�@ 2�q��ٿ�\����@�52}��3@����ې!?�hw��+�@ 2�q��ٿ�\����@�52}��3@����ې!?�hw��+�@ 2�q��ٿ�\����@�52}��3@����ې!?�hw��+�@����ٿ��%����@�����3@c݌���!?��3��+�@����ٿ��%����@�����3@c݌���!?��3��+�@q/o��ٿ<�k����@!mq��3@�ؑS��!?&eb��+�@h;"籙ٿ�#����@�'�#��3@Pu����!?5}ְ�+�@h;"籙ٿ�#����@�'�#��3@Pu����!?5}ְ�+�@h;"籙ٿ�#����@�'�#��3@Pu����!?5}ְ�+�@��fҲ�ٿ�k����@"�M���3@H�o�p�!?�{��+�@3jZH��ٿ$qa����@t2_��3@vg��!?�ų�+�@��A��ٿ�ť���@a�/��3@��V�!?
=���+�@��p��ٿM�N����@��#J��3@@����!?�����+�@��p��ٿM�N����@��#J��3@@����!?�����+�@�Z���ٿ�`�����@M�D_��3@�V���!?#�Ҷ�+�@jx����ٿ�b�����@������3@w���a�!?�@���+�@��ƶ�ٿ��ʐ���@mF���3@���s�!?7�e��+�@[	�岙ٿ�`����@ zaS��3@�7��Ր!?W�&��+�@[	�岙ٿ�`����@ zaS��3@�7��Ր!?W�&��+�@[	�岙ٿ�`����@ zaS��3@�7��Ր!?W�&��+�@SV��ٿ�qp����@hz ���3@�"�!?(λ��+�@SV��ٿ�qp����@hz ���3@�"�!?(λ��+�@�w���ٿ��J����@�8��3@cds��!?���+�@�s�2��ٿUU����@N�0���3@m�ƌ�!?p����+�@9�X��ٿA*����@6���3@fᬘ��!?7���+�@�$	L��ٿ�6�����@�����3@��>��!?�����+�@����ٿG�����@��B��3@c�H�ِ!?��:��+�@�iCƬ�ٿM�����@슌���3@>1�k�!?*郱�+�@Fw����ٿ'�ߥ���@60�u��3@��kސ!?TU���+�@�B�ѵ�ٿ������@�dp��3@u4А!?@���+�@aKd��ٿ)#D����@�.i��3@U8��!?��T��+�@aKd��ٿ)#D����@�.i��3@U8��!?��T��+�@%*d��ٿ������@�:���3@�ι��!?����+�@%*d��ٿ������@�:���3@�ι��!?����+�@�+4캙ٿ�}�����@�q���3@��US��!?{�2��+�@A߯��ٿe5�����@m� }��3@F��Ґ!?B�(��+�@��n}��ٿY6����@ʢϔ��3@�t���!?����+�@��n}��ٿY6����@ʢϔ��3@�t���!?����+�@�s�^��ٿB�=����@{����3@��vM�!?�]��+�@ �����ٿ+����@j����3@Fvr�=�!?�/-��+�@w>���ٿ7iJ���@�J����3@v�u&h�!?��ǵ�+�@�>���ٿ�n�z���@v����3@Ȓo<T�!?�aX��+�@	�B㹙ٿ�0v���@������3@ݺ�/`�!?m���+�@��F4��ٿC?pu���@l}����3@f����!?�y��+�@�u¼�ٿ�n.s���@�Q����3@�ᦢ�!?�n��+�@�u¼�ٿ�n.s���@�Q����3@�ᦢ�!?�n��+�@V�lؾ�ٿ؇Tt���@A����3@C��D��!?�ح�+�@ ��.��ٿ@pn���@'$�C��3@ތ�;��!?�_q��+�@ ��.��ٿ@pn���@'$�C��3@ތ�;��!?�_q��+�@�����ٿ��n���@�:���3@���]��!?�
f��+�@������ٿc��{���@ݮ���3@i�N��!?����+�@�4�͸�ٿ���p���@p%����3@r�U)�!?d���+�@?A���ٿW�.}���@�����3@'Z��!?.	��+�@?A���ٿW�.}���@�����3@'Z��!?.	��+�@��T%��ٿ������@/X����3@Z����!?�u���+�@�EZ��ٿV�����@�����3@~�����!?l�T��+�@�EZ��ٿV�����@�����3@~�����!?l�T��+�@�EZ��ٿV�����@�����3@~�����!?l�T��+�@'����ٿ������@I�q��3@~[��!?�V#��+�@���"��ٿ��ƚ���@$�Et��3@/��ِ!?�����+�@(����ٿ?����@s����3@���I��!?����+�@.�w��ٿz������@����3@奎K��!?�(��+�@�����ٿ�z�����@��J5��3@
ք�!?���+�@�����ٿ�z�����@��J5��3@
ք�!?���+�@C\򄪙ٿ�ګ����@P�q��3@d�q��!?�wQ��+�@�G�ª�ٿ�N����@�|]��3@n�'+��!?��`��+�@B��z��ٿ��t����@�u9���3@�eI ��!?�EC��+�@�	d���ٿƲͼ���@N�;���3@*NC�!?v��+�@�	d���ٿƲͼ���@N�;���3@*NC�!?v��+�@lrR��ٿ��~����@�}����3@�h�!?K�k��+�@j�{��ٿ������@ీ#��3@x
Hk�!?��n��+�@�L�9��ٿ}����@2�����3@�Q��!?�б��+�@��vw��ٿ'�����@&o/'��3@���EƐ!?̕	��+�@X�)K��ٿ�����@�q��3@T<����!?����+�@v#����ٿҨ����@K�6���3@�I�2w�!?_s��+�@��aU��ٿyM�����@S����3@�� ��!?{��+�@�7���ٿו����@����3@�X�>��!?��*��+�@��/��ٿ}غ����@q��{��3@=G�f��!?�1!��+�@��3��ٿic�����@_�����3@�~#��!?4W���+�@B�碙ٿu�����@A��}��3@щ�!?L%��+�@���ޛ�ٿ�ً����@ �����3@�	��!?�2"��+�@��ӷ��ٿ�-g����@�$���3@����j�!?�X��+�@��ӷ��ٿ�-g����@�$���3@����j�!?�X��+�@��Y��ٿ�x����@d�����3@��g���!?~;H��+�@;ol��ٿ��Ѻ���@�:�1��3@9�h���!?
���+�@% 9��ٿ7=����@���5��3@Z�-Nv�!?�)I��+�@�#����ٿ;S:����@�|�N��3@�}���!?ZT���+�@�#����ٿ;S:����@�|�N��3@�}���!?ZT���+�@1����ٿnZ�����@����3@,m��}�!?�d���+�@9wV��ٿ==E����@MI	��3@������!?��ޞ�+�@?�p�}�ٿ��N����@�{Zj��3@�1ߝ�!?_����+�@Y�/�ٿ������@U�[���3@�y�ͤ�!?��c��+�@K賅t�ٿ+�����@��V���3@a�ӝ��!?u2��+�@K賅t�ٿ+�����@��V���3@a�ӝ��!?u2��+�@^=��ٿi������@�џ���3@��Fpʐ!?��e��+�@��Oύ�ٿL�=����@�r���3@ASF�ݐ!?�/��+�@ם�a��ٿ������@�����3@�Z���!?��ې�+�@��p�ٿ�J�����@	��w��3@ �\DԐ!?:dH�+�@��p�ٿ�J�����@	��w��3@ �\DԐ!?:dH�+�@��p�ٿ�J�����@	��w��3@ �\DԐ!?:dH�+�@QxzIV�ٿ3_K ��@���^��3@!5�Ṑ!?v��l�+�@
f�Y�ٿ�n� ��@��w 4@��:8Ґ!?L"rf�+�@h~K�ٿXeF ��@���b��3@4���!?�Dvc�+�@!^��x�ٿ�z����@A.mt��3@�m�f�!?}i#��+�@��NY�ٿX9�! ��@��z  4@b���!?��Li�+�@��NY�ٿX9�! ��@��z  4@b���!?��Li�+�@��NY�ٿX9�! ��@��z  4@b���!?��Li�+�@��NY�ٿX9�! ��@��z  4@b���!?��Li�+�@���&��ٿN�6����@ ��3@�k@��!?OK���+�@�yLn��ٿ%&v����@'1���3@�^���!?��ω�+�@��[��ٿ�N�����@���b��3@
��O��!?����+�@��[��ٿ�N�����@���b��3@
��O��!?����+�@|U<�ٿN`�����@�"W��3@���B��!?�='��+�@ϫ8b��ٿGJ�����@��E��3@d��Đ!?��#��+�@]��ʙٿ�q?����@��a��3@���Ж�!?�	\��+�@�.u鯙ٿ�����@EOQ��3@z�O��!?]�p��+�@�.u鯙ٿ�����@EOQ��3@z�O��!?]�p��+�@�.u鯙ٿ�����@EOQ��3@z�O��!?]�p��+�@P��咙ٿ�@�����@����3@́뗐!?�f��+�@P��咙ٿ�@�����@����3@́뗐!?�f��+�@P��咙ٿ�@�����@����3@́뗐!?�f��+�@�~Vc�ٿ:�i����@rO����3@.��Ԑ!?��Bt�+�@GΕFU�ٿ�K	 ��@oO 4@A��L��!?��_�+�@�(Szf�ٿk�o����@-�n< 4@:�&沐!?uhs�+�@b��w�ٿҥ�����@���t 4@��٬�!?2Rz�+�@Y���P�ٿ#64  ��@�tQ� 4@2ŸD��!?�be�+�@��F�ٿ{�2 ��@�=& 4@v���!?ն Z�+�@8���t�ٿ1Ɉ����@�X���3@�����!?�G���+�@�h�i�ٿ��� ��@�6����3@���Ő!?��}��+�@޵���ٿ�V����@��+��3@i\;�ΐ!?�5���+�@u	ۺ��ٿ�g����@]��'��3@`��@ؐ!?�ș��+�@�e�u�ٿ��� ��@V�?0��3@_C
	��!?�}�+�@z5H�e�ٿ�< ��@	=����3@�;a<��!?��7{�+�@���yW�ٿ�V ��@��̂��3@ �g�!?A~Y}�+�@���yW�ٿ�V ��@��̂��3@ �g�!?A~Y}�+�@��Yg�ٿe�Z ��@��t4��3@�*�J�!?a�x�+�@${�p�ٿ������@�U���3@���|��!?�T5�+�@${�p�ٿ������@�U���3@���|��!?�T5�+�@M�
�p�ٿdɃ ��@dw��3@�Q�䃐!?A	z�+�@r�|v��ٿ�i�����@�QI���3@�R�y�!?[���+�@��u?��ٿ��\����@	U����3@_ۤ�{�!?�����+�@��u?��ٿ��\����@	U����3@_ۤ�{�!?�����+�@�.�	��ٿ�FS����@%�����3@�Qݿ�!?�]��+�@S~����ٿ3�����@0\����3@-q����!?�G}��+�@������ٿ������@^����3@��3|�!?]����+�@OEH^W�ٿ��`����@!f�o 4@sp�l�!?�xr�+�@>��$C�ٿ��:# ��@�<,���3@���!?ļ�f�+�@/�#)�ٿT��; ��@)�� 4@���ِ!?���L�+�@/�#)�ٿT��; ��@)�� 4@���ِ!?���L�+�@���':�ٿx@�" ��@��#_ 4@��g�!?��Z^�+�@"u0l8�ٿ�4� ��@�e=4 4@n-Ss,�!?!�U�+�@/�]Q�ٿ������@�/N 4@�殨��!?w��`�+�@�5�:�ٿaU ��@��u	 4@ m��!?��I�+�@�5�:�ٿaU ��@��u	 4@ m��!?��I�+�@��x$�ٿ_�. ��@H��� 4@B[�, �!?�}�J�+�@�;ϣ��ٿ�n�J ��@�8��	 4@-F��<�!?���+�@  ��,�ٿ<�� ��@�Y`A 4@��޾-�!?$x�6�+�@  ��,�ٿ<�� ��@�Y`A 4@��޾-�!?$x�6�+�@�?)�ٿ4� ��@X�Q 4@�%�5�!?:�K*�+�@#Gr���ٿ�� ��@��K� 4@[�,1�!?:���+�@#Gr���ٿ�� ��@��K� 4@[�,1�!?:���+�@#Gr���ٿ�� ��@��K� 4@[�,1�!?:���+�@#Gr���ٿ�� ��@��K� 4@[�,1�!?:���+�@#Gr���ٿ�� ��@��K� 4@[�,1�!?:���+�@�/�fؘٿ�� ��@¶��% 4@˻G�V�!?�����+�@�d[٘ٿ(T/7 ��@=�E 4@^v3�!�!?����+�@�)�З�ٿ��Q����@��u� 4@�=�ɛ�!?dJZ��+�@8��~�ٿP������@u�� 4@}����!?�0�n�+�@�=s���ٿnd����@�u� 4@�����!?�h[�+�@��4ؙٿ��'s���@�`=� 4@���Ő!?����+�@։D�P�ٿ_��J���@��B���3@�ҽ�L�!?k��+�@։D�P�ٿ_��J���@��B���3@�ҽ�L�!?k��+�@։D�P�ٿ_��J���@��B���3@�ҽ�L�!?k��+�@։D�P�ٿ_��J���@��B���3@�ҽ�L�!?k��+�@k5�<v�ٿ�u4����@x�� 4@��g2�!?�B{l�+�@k5�<v�ٿ�u4����@x�� 4@��g2�!?�B{l�+�@��r7��ٿ�VSd���@w��� 4@�P9�!?Ը��+�@�ufe?�ٿ��
���@��� 4@(��/��!?5��+�@�ufe?�ٿ��
���@��� 4@(��/��!?5��+�@�?Y�ʙٿ��_����@��  4@�g$��!?�p��+�@{󈲘ٿR�W ��@N�� 4@��l��!?�+�@{󈲘ٿR�W ��@N�� 4@��l��!?�+�@{󈲘ٿR�W ��@N�� 4@��l��!?�+�@{󈲘ٿR�W ��@N�� 4@��l��!?�+�@hM��$�ٿ�(����@��e� 4@��
���!?7T&X�+�@hM��$�ٿ�(����@��e� 4@��
���!?7T&X�+�@�u%|�ٿc�����@�oe���3@���֐!?(I���+�@�u%|�ٿc�����@�oe���3@���֐!?(I���+�@4:�庙ٿ@�by���@�χ 4@0RZ�Ր!?��$��+�@��%D	�ٿ�`
���@�-/U 4@�3�lא!?��G�+�@��%D	�ٿ�`
���@�-/U 4@�3�lא!?��G�+�@\>*|�ٿ�g[g���@/I 4@;F��̐!?S���+�@(+j~}�ٿ���F ��@��� 4@�c��!?����+�@�_�#N�ٿ��m ��@ȧx# 4@K��r�!?8����+�@��:�R�ٿ�e�5��@��1�5 4@.�P�c�!?qN�A�+�@��:�R�ٿ�e�5��@��1�5 4@.�P�c�!?qN�A�+�@��:�R�ٿ�e�5��@��1�5 4@.�P�c�!?qN�A�+�@��:�R�ٿ�e�5��@��1�5 4@.�P�c�!?qN�A�+�@:���ٿIk�� ��@|1�H 4@�Vh�Ő!?V�z�+�@]��ٿm�����@68��  4@�`���!?�3I�+�@��F���ٿ�w�h��@���Y 4@-�߽!?��j��+�@��F���ٿ�w�h��@���Y 4@-�߽!?��j��+�@��F���ٿ�w�h��@���Y 4@-�߽!?��j��+�@��F���ٿ�w�h��@���Y 4@-�߽!?��j��+�@��F���ٿ�w�h��@���Y 4@-�߽!?��j��+�@]wT���ٿ�؂� ��@�J�? 4@��KD��!?�j��+�@  �d�ٿ������@r�5� 4@��(ِ!?bg��+�@  �d�ٿ������@r�5� 4@��(ِ!?bg��+�@  �d�ٿ������@r�5� 4@��(ِ!?bg��+�@_���J�ٿ>Z����@�I 4@PD�۪�!?a����+�@�f}�ٿ�I�����@$9mc 4@{@Ґ!?��'o�+�@�f}�ٿ�I�����@$9mc 4@{@Ґ!?��'o�+�@�1�ܕٿy���@$�m 4@"TCB�!?�ݪ�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@*�(J��ٿ�����@��S� 4@�/�*!?�[m�+�@K����ٿ�k�K��@���"4@��\�6�!?�]&�+�@��k�ٿJ�L��@�+)4@J6��8�!?�*���+�@1Ѻ	�ٿ�^����@�l�VX4@D�)F�!?�T<�+�@���ٿ��S���@\���84@����!?�dV��+�@E��ōٿ��F��@�J��Z4@�����!?�Z���+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@'��E�ٿ�� ���@H-7)�4@<FO�!?�)�$�+�@8�#{wٿ"p���@r !��4@4/^ې!?�\���+�@��a���ٿ�m=��@*�/��4@�%��,�!?�ӆ�+�@��a���ٿ�m=��@*�/��4@�%��,�!?�ӆ�+�@��a���ٿ�m=��@*�/��4@�%��,�!?�ӆ�+�@��a���ٿ�m=��@*�/��4@�%��,�!?�ӆ�+�@��a���ٿ�m=��@*�/��4@�%��,�!?�ӆ�+�@��i�ٿ��C���@o�,S�4@�r��!?�⦁�+�@��i�ٿ��C���@o�,S�4@�r��!?�⦁�+�@|Ũ`q�ٿkQ�	��@�0#4@���!??q<Q�+�@|Ũ`q�ٿkQ�	��@�0#4@���!??q<Q�+�@�t���ٿ"D;���@D3�{�4@�B���!?e��s�+�@�t���ٿ"D;���@D3�{�4@�B���!?e��s�+�@�t���ٿ"D;���@D3�{�4@�B���!?e��s�+�@�t���ٿ"D;���@D3�{�4@�B���!?e��s�+�@�t���ٿ"D;���@D3�{�4@�B���!?e��s�+�@`��ڝ�ٿ�on
��@��VS4@�):R��!?rk~��+�@`��ڝ�ٿ�on
��@��VS4@�):R��!?rk~��+�@`��ڝ�ٿ�on
��@��VS4@�):R��!?rk~��+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@���M��ٿbL5	��@�H &4@��2ȅ�!?g����+�@|�1͇ٿ������@.�n*4@���!?V���+�@|�1͇ٿ������@.�n*4@���!?V���+�@�c�le�ٿ��	��@^�a�R4@�ll�ܐ!?��`�+�@�c�le�ٿ��	��@^�a�R4@�ll�ܐ!?��`�+�@�p�!��ٿ3����@؇Lؖ4@�#�:"�!?%�9��+�@��4�Ʉٿ�:[
��@t�BG�4@�O<��!?��}e�+�@��4�Ʉٿ�:[
��@t�BG�4@�O<��!?��}e�+�@��{|ٿ�����@�@Q�4@��x�Ȑ!?޺g�+�@��{|ٿ�����@�@Q�4@��x�Ȑ!?޺g�+�@���+�ٿ=cH� ��@�b�4@tJ�#��!?��l�+�@���+�ٿ=cH� ��@�b�4@tJ�#��!?��l�+�@���+�ٿ=cH� ��@�b�4@tJ�#��!?��l�+�@G�o��ٿ��[��@Y
�7U4@��Ͳ�!?�PX�+�@G�o��ٿ��[��@Y
�7U4@��Ͳ�!?�PX�+�@G�o��ٿ��[��@Y
�7U4@��Ͳ�!?�PX�+�@���Q�ٿ=��b��@sq�#�4@eP�*�!?d�j��+�@���Q�ٿ=��b��@sq�#�4@eP�*�!?d�j��+�@���Q�ٿ=��b��@sq�#�4@eP�*�!?d�j��+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@#��}ٿ�w�W��@��1�4@�{Xِ!?R,���+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@~�#Y��ٿ�>��@�x���4@NHXj�!?wo]��+�@�4J��yٿ��
��@�)F�4@�y1�А!?#���+�@�I���}ٿ��݉��@(�0��4@#~v�F�!?F).�+�@�I���}ٿ��݉��@(�0��4@#~v�F�!?F).�+�@�I���}ٿ��݉��@(�0��4@#~v�F�!?F).�+�@�I���}ٿ��݉��@(�0��4@#~v�F�!?F).�+�@(�i�ٿű'���@��i�4@�t�6(�!?;�Ch�+�@f�>��ٿ�c����@pŘ�4@s�1�!?<���+�@f�>��ٿ�c����@pŘ�4@s�1�!?<���+�@f�>��ٿ�c����@pŘ�4@s�1�!?<���+�@f�>��ٿ�c����@pŘ�4@s�1�!?<���+�@�����ٿ�?]d���@u�s�4@��I@�!?7[��+�@�;e곉ٿ��>m ��@��C4@	�K��!?d'iV�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@���{�ٿ�ra����@'	�4@�����!?�4�b�+�@Q}'��ٿ�
����@�M�4@��!?�$"5�+�@�'�� �ٿ�B>���@�\�ۉ4@�Ո�2�!?_���+�@����ٿ�zb����@���4@AO��2�!?�����+�@����ٿ�zb����@���4@AO��2�!?�����+�@����ٿ�zb����@���4@AO��2�!?�����+�@����ٿ�zb����@���4@AO��2�!?�����+�@�f�Cp�ٿ�%���@�Km4@F9r9L�!?+�l>�+�@EP���zٿ:. 8��@�D�.'4@eV�a2�!?����+�@EP���zٿ:. 8��@�D�.'4@eV�a2�!?����+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@:F�m�ٿ��Y��@<�O�4@g��ܐ!?1p��+�@T�𝶇ٿjU����@���-4@�z�ΐ!?��|�+�@�Tv�яٿ�͈�
��@l�!H 4@�$��ɐ!?�I)#�+�@�Tv�яٿ�͈�
��@l�!H 4@�$��ɐ!?�I)#�+�@=��.��ٿ���7���@���;4@L�%��!?Ik�+�@�PQ���ٿ�Ӈ���@�6��`4@���!?Ò��+�@�Vٿ"�����@�i�4@�f�@��!?N8��+�@�Vٿ"�����@�i�4@�f�@��!?N8��+�@�Vٿ"�����@�i�4@�f�@��!?N8��+�@�Vٿ"�����@�i�4@�f�@��!?N8��+�@�Vٿ"�����@�i�4@�f�@��!?N8��+�@|WR�{ٿ�����@�j_�a4@	�Xݐ!?�cNC�+�@|WR�{ٿ�����@�j_�a4@	�Xݐ!?�cNC�+�@|WR�{ٿ�����@�j_�a4@	�Xݐ!?�cNC�+�@|WR�{ٿ�����@�j_�a4@	�Xݐ!?�cNC�+�@|WR�{ٿ�����@�j_�a4@	�Xݐ!?�cNC�+�@��)�ٿ�nԟ��@iX��4@����!?��:�+�@�@z�'�ٿ>�;��@�����4@�J��!?8/���+�@�K<���ٿ��5P��@n~�}�4@��ΐ!?*�5�+�@�K<���ٿ��5P��@n~�}�4@��ΐ!?*�5�+�@�K<���ٿ��5P��@n~�}�4@��ΐ!?*�5�+�@�K<���ٿ��5P��@n~�}�4@��ΐ!?*�5�+�@�K<���ٿ��5P��@n~�}�4@��ΐ!?*�5�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@���ٿ�t���@,���4@⒃�ǐ!?ϐ�O�+�@HmL��ٿ}TN���@ݼ��64@Hb�{��!?�w�V�+�@HmL��ٿ}TN���@ݼ��64@Hb�{��!?�w�V�+�@HmL��ٿ}TN���@ݼ��64@Hb�{��!?�w�V�+�@HmL��ٿ}TN���@ݼ��64@Hb�{��!?�w�V�+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@7�]�ٿ��J��@<z��4@�7��!?TN4��+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@ ��)R�ٿ������@>I�4@�7��ː!?����+�@~�����ٿNE�����@�b�84@��iY�!?/F���+�@~�����ٿNE�����@�b�84@��iY�!?/F���+�@~�����ٿNE�����@�b�84@��iY�!?/F���+�@~�����ٿNE�����@�b�84@��iY�!?/F���+�@~�����ٿNE�����@�b�84@��iY�!?/F���+�@6h/���ٿ�/���@�#�`4@if����!?�f���+�@6h/���ٿ�/���@�#�`4@if����!?�f���+�@6h/���ٿ�/���@�#�`4@if����!?�f���+�@6h/���ٿ�/���@�#�`4@if����!?�f���+�@s�j��ٿ�uo����@�z��G4@Q�8�Đ!?Kz���+�@������ٿ��_+��@��s�4@�qd��!?��^��+�@������ٿ��_+��@��s�4@�qd��!?��^��+�@������ٿ��_+��@��s�4@�qd��!?��^��+�@������ٿ��_+��@��s�4@�qd��!?��^��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@pD8��ٿ>����@��=�4@MJ�!?�-I��+�@�禍�ٿ������@�f`4@Ĳ���!?J:Ə�+�@���e�ٿ`����@5ayu4@Ͼ���!?�|,�+�@���e�ٿ`����@5ayu4@Ͼ���!?�|,�+�@���e�ٿ`����@5ayu4@Ͼ���!?�|,�+�@X�1\��ٿ�.���@���ǩ4@��뫐!?�M���+�@X�1\��ٿ�.���@���ǩ4@��뫐!?�M���+�@X�1\��ٿ�.���@���ǩ4@��뫐!?�M���+�@e�ĩ~ٿ9�c���@/!��4@詝�!?�\[a�+�@e�ĩ~ٿ9�c���@/!��4@詝�!?�\[a�+�@\4����ٿ�U���@_u�8�4@	V).�!?��|��+�@\4����ٿ�U���@_u�8�4@	V).�!?��|��+�@�1�@�ٿmUcxՇ�@��^W54@S���U�!?�W�+�@�1�@�ٿmUcxՇ�@��^W54@S���U�!?�W�+�@�1�@�ٿmUcxՇ�@��^W54@S���U�!?�W�+�@ՠ�-4zٿ"��fه�@��)�	4@fi��@�!?g�<Q�+�@�C�4ٿ'�ɇ�@F4�w4@��+�!?==a,�@�C�4ٿ'�ɇ�@F4�w4@��+�!?==a,�@ZyO�R�ٿŕZ���@_��I�
4@�u�EB�!?�Zq�,�@ZyO�R�ٿŕZ���@_��I�
4@�u�EB�!?�Zq�,�@ZyO�R�ٿŕZ���@_��I�
4@�u�EB�!?�Zq�,�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@T����ٿ�.����@���pL4@�p7��!?�}��+�@���h��ٿ�y?��@D�QӘ4@T�}��!?��!��+�@���h��ٿ�y?��@D�QӘ4@T�}��!?��!��+�@!��c�ٿ�����@}��S4@W�O8�!?Q�N��+�@!��c�ٿ�����@}��S4@W�O8�!?Q�N��+�@!��c�ٿ�����@}��S4@W�O8�!?Q�N��+�@!��c�ٿ�����@}��S4@W�O8�!?Q�N��+�@6�9Ӊٿ�r�/��@��&Z�4@�B?���!?�:� �+�@6�9Ӊٿ�r�/��@��&Z�4@�B?���!?�:� �+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@PJ�V��ٿn]3$��@Ʈ&_4@�[b���!?��6g�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@���5�ٿe�"}���@LΓ��4@�í��!?��o�+�@��m�ٿm->sŇ�@��i��4@� ^r�!?�[�,�@��_ �ٿfl�7���@uL��g4@�\�8��!?��'�,�@��_ �ٿfl�7���@uL��g4@�\�8��!?��'�,�@��_ �ٿfl�7���@uL��g4@�\�8��!?��'�,�@��_ �ٿfl�7���@uL��g4@�\�8��!?��'�,�@��_ �ٿfl�7���@uL��g4@�\�8��!?��'�,�@��zrG�ٿ��q���@�ag.�4@� � ��!?EsIe�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@� ƪD�ٿ�k"I��@�~Sg�4@D���!?~�A�+�@}PH���ٿD��z��@k�Uo�4@7E��!?��L*�+�@}PH���ٿD��z��@k�Uo�4@7E��!?��L*�+�@}PH���ٿD��z��@k�Uo�4@7E��!?��L*�+�@-�~ٿ/�2(��@���j4@U�%��!?k����+�@���ٿy�ԃ��@/~2�4@�}QK�!?͑ �+�@���ٿy�ԃ��@/~2�4@�}QK�!?͑ �+�@���ٿy�ԃ��@/~2�4@�}QK�!?͑ �+�@giQF�ٿ��:��@х;�)4@͎����!?p�֜+�@� N���ٿ��bPӇ�@���4@5l�!?��7��+�@*�c(��ٿ #���@��՜4@S��x#�!?��y��+�@*�c(��ٿ #���@��՜4@S��x#�!?��y��+�@�}�#ڍٿo#E���@-z��g4@�ok�А!?d�$,�@�}�#ڍٿo#E���@-z��g4@�ok�А!?d�$,�@�}�#ڍٿo#E���@-z��g4@�ok�А!?d�$,�@�}�#ڍٿo#E���@-z��g4@�ok�А!?d�$,�@3��ܒٿm*9��@A� ��4@���<�!?��mu�+�@�e�v�zٿQ�l@��@1�)Q4@���!?Mw��\+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@A ��ٿ^�E��@S�5�4@���Q��!?�)}x�+�@�j��v�ٿ
%�� ��@i��4@U)a��!?_,p��+�@�Lٕ�ٿ���#}��@͡��4@�֌��!?gW\+�@�Lٕ�ٿ���#}��@͡��4@�֌��!?gW\+�@� jB��ٿԄ��k��@�Q�A4@��۠�!?�D�?f+�@� jB��ٿԄ��k��@�Q�A4@��۠�!?�D�?f+�@� jB��ٿԄ��k��@�Q�A4@��۠�!?�D�?f+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@�-��_�ٿ�&'���@|�� 4@���>��!?���.K+�@z�,�Y�ٿf�t! ��@x�a4@����!?F`af�+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@�&-�ٿ
�4r��@끍Y4@�2�_�!?(8�]+�@d�ܹ�ٿ�&~���@rQR->4@�řF��!?����;+�@d�ܹ�ٿ�&~���@rQR->4@�řF��!?����;+�@d�ܹ�ٿ�&~���@rQR->4@�řF��!?����;+�@d�ܹ�ٿ�&~���@rQR->4@�řF��!?����;+�@��"<�ٿy�����@�h>d4@2��T�!?[��I,�@��"<�ٿy�����@�h>d4@2��T�!?[��I,�@��"<�ٿy�����@�h>d4@2��T�!?[��I,�@��"<�ٿy�����@�h>d4@2��T�!?[��I,�@@�~H�ٿ0���y��@�gx=a4@�����!?0�KS-�@@�~H�ٿ0���y��@�gx=a4@�����!?0�KS-�@�AM�c�ٿ��詮��@R�3%4@Z�q��!?+E�P+-�@�AM�c�ٿ��詮��@R�3%4@Z�q��!?+E�P+-�@�AM�c�ٿ��詮��@R�3%4@Z�q��!?+E�P+-�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@#�]�ՃٿYP)��@?l��b4@I�^X��!?Bt�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@�K��ٿ>�1�:��@�!�4@@�1!?	��p�/�@��+Mzٿ>\Bj)��@����4@�.5��!?�n'�)�@��+Mzٿ>\Bj)��@����4@�.5��!?�n'�)�@��+Mzٿ>\Bj)��@����4@�.5��!?�n'�)�@��+Mzٿ>\Bj)��@����4@�.5��!?�n'�)�@��+Mzٿ>\Bj)��@����4@�.5��!?�n'�)�@n�>�g�ٿ5anB���@Q�v�4@���-ߐ!?�~R&6/�@n�>�g�ٿ5anB���@Q�v�4@���-ߐ!?�~R&6/�@�
�>o�ٿUs 3o��@$L3�;4@#����!?\Kp,�@�
�>o�ٿUs 3o��@$L3�;4@#����!?\Kp,�@�
�>o�ٿUs 3o��@$L3�;4@#����!?\Kp,�@{����ٿKq��Q��@���UX 4@���鐐!?��y�2�@{����ٿKq��Q��@���UX 4@���鐐!?��y�2�@�y��!�ٿ�ds҇�@��2X�4@-��!?��%Q�+�@:�*6��ٿ�,��ʇ�@}��f4@�^W��!?�� �,�@:�*6��ٿ�,��ʇ�@}��f4@�^W��!?�� �,�@:�*6��ٿ�,��ʇ�@}��f4@�^W��!?�� �,�@:�*6��ٿ�,��ʇ�@}��f4@�^W��!?�� �,�@:�*6��ٿ�,��ʇ�@}��f4@�^W��!?�� �,�@��J��ٿ�B ���@7Nؾ4@��֪��!?j��t'&�@��J��ٿ�B ���@7Nؾ4@��֪��!?j��t'&�@��J��ٿ�B ���@7Nؾ4@��֪��!?j��t'&�@��J��ٿ�B ���@7Nؾ4@��֪��!?j��t'&�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@*��ö�ٿ �/% ��@\���4@�sn`��!?���B�,�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@ހ�FƋٿK��P��@7~��`4@3��E�!?�d�~*�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@`9z8~�ٿ'�����@��q��4@�[[ː!?X1�.�@P$�ٿ:�n� ��@�z���4@�g��!?��J�+�@P$�ٿ:�n� ��@�z���4@�g��!?��J�+�@�U-�ٿ�\�f���@@j#*�4@�
-]N�!?��Rxm1�@�U-�ٿ�\�f���@@j#*�4@�
-]N�!?��Rxm1�@�U-�ٿ�\�f���@@j#*�4@�
-]N�!?��Rxm1�@�U-�ٿ�\�f���@@j#*�4@�
-]N�!?��Rxm1�@�U-�ٿ�\�f���@@j#*�4@�
-]N�!?��Rxm1�@����ٿ�j��C��@�e��4@w�"���!?��|�)�@����ٿ�j��C��@�e��4@w�"���!?��|�)�@`m�H�ٿa����@J���4@/{4O�!?�XĸB(�@`m�H�ٿa����@J���4@/{4O�!?�XĸB(�@`m�H�ٿa����@J���4@/{4O�!?�XĸB(�@$btU}ٿG�h����@�]6�4@Ag�$�!?���r��@�t��}ٿ17��
��@�bKR4@��燐!?���Ô!�@���jٿM�91Ӑ�@f뜭�4@ό5�|�!?��"�@���jٿM�91Ӑ�@f뜭�4@ό5�|�!?��"�@���jٿM�91Ӑ�@f뜭�4@ό5�|�!?��"�@����܁ٿ���J��@Q����4@�yŗ��!?��eY"�@����܁ٿ���J��@Q����4@�yŗ��!?��eY"�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@ޣν�ٿd�HJ8��@�m[U4@�^R˚�!?���&�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@d7ڵ��ٿ��%E��@�/M�4@s"�ϐ!?J��!�@�MU�ٿX����@e�>q�4@#�G�s�!?ӏ����@�MU�ٿX����@e�>q�4@#�G�s�!?ӏ����@�<�ٿ*��B��@�g$:�4@�N�!?#D�`6
�@�<�ٿ*��B��@�g$:�4@�N�!?#D�`6
�@~Q6x�}ٿ�3~�w��@0�F�m4@�s��!?�N͟Z��@~Q6x�}ٿ�3~�w��@0�F�m4@�s��!?�N͟Z��@K{��ٿ�FRo���@�@%-4@�ǘ�!?�po�&�@K{��ٿ�FRo���@�@%-4@�ǘ�!?�po�&�@K{��ٿ�FRo���@�@%-4@�ǘ�!?�po�&�@K{��ٿ�FRo���@�@%-4@�ǘ�!?�po�&�@�~��ٿ�������@D���4@p����!?�K�8��@�~��ٿ�������@D���4@p����!?�K�8��@�~��ٿ�������@D���4@p����!?�K�8��@�|��ٿ$����@���	4@�]9�ِ!?�,��k��@�|��ٿ$����@���	4@�]9�ِ!?�,��k��@�|��ٿ$����@���	4@�]9�ِ!?�,��k��@mdFr�ٿ���1��@�iv+P4@��R��!?�:)��@a�MSe�ٿ|וv���@j��4@"��]E�!?2�`;��@a�MSe�ٿ|וv���@j��4@"��]E�!?2�`;��@a�MSe�ٿ|וv���@j��4@"��]E�!?2�`;��@��t̉ٿ�9(Y/��@��E4@in.���!?����@��t̉ٿ�9(Y/��@��E4@in.���!?����@��t̉ٿ�9(Y/��@��E4@in.���!?����@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�N� �ٿ	3�����@Kq�1O4@%�N�!?<��G3��@�~,�A~ٿ��w�@���/I4@��-���!?*�>����@�~,�A~ٿ��w�@���/I4@��-���!?*�>����@�~,�A~ٿ��w�@���/I4@��-���!?*�>����@�~,�A~ٿ��w�@���/I4@��-���!?*�>����@Ү�/K�ٿ�fi �7�@æ~��4@E��{�!?J5��x�@Ү�/K�ٿ�fi �7�@æ~��4@E��{�!?J5��x�@Ү�/K�ٿ�fi �7�@æ~��4@E��{�!?J5��x�@��+��~ٿ$����?�@�4��4@��*7��!?�g��o�@��+��~ٿ$����?�@�4��4@��*7��!?�g��o�@��+��~ٿ$����?�@�4��4@��*7��!?�g��o�@�+iҠ�ٿ&.�Bq�@�(q^�4@��~��!? F�9��@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@U�rgX�ٿ&`��d�@HP[�4@܇nx&�!?�I�7�J�@�����ٿZ=�y`��@��?�74@���ې!?�dka,��@�����ٿZ=�y`��@��?�74@���ې!?�dka,��@�����ٿZ=�y`��@��?�74@���ې!?�dka,��@�����ٿZ=�y`��@��?�74@���ې!?�dka,��@�����ٿZ=�y`��@��?�74@���ې!?�dka,��@.�>=�ٿ�[dg�E�@��ș4@�Q��$�!?>,��j�@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@�tNh�ٿ�6�����@�rK�4@਷'�!?�������@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@����6�ٿ�Ů^���@^���44@�HUy��!?:�fl��@�=B,�ٿ�Tu�o �@4�U+4@�a���!?�"����@�7�K�ٿU�6���@6a��4@����ʐ!?�c_��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@�5
��ٿ��No��@u�7\@4@�Cރ��!?�� ��@p�{�ٿ.Fr�%��@y,3�4@�h�!?'ޗѸ��@p�{�ٿ.Fr�%��@y,3�4@�h�!?'ޗѸ��@p�{�ٿ.Fr�%��@y,3�4@�h�!?'ޗѸ��@��ZaD�ٿڈ�$���@mM�*4@kE���!?uk�h��@��ZaD�ٿڈ�$���@mM�*4@kE���!?uk�h��@��ZaD�ٿڈ�$���@mM�*4@kE���!?uk�h��@�~�o�ٿ�#g��@�'�Q4@0y s��!?�C�N��@�e ~�ٿ���?�@/����4@mV�	�!?��0Z�o�@�e ~�ٿ���?�@/����4@mV�	�!?��0Z�o�@�e ~�ٿ���?�@/����4@mV�	�!?��0Z�o�@�e ~�ٿ���?�@/����4@mV�	�!?��0Z�o�@�e ~�ٿ���?�@/����4@mV�	�!?��0Z�o�@���*��ٿ����>k�@1�L4@�S���!?ǬZXDI�@���*��ٿ����>k�@1�L4@�S���!?ǬZXDI�@5�=PƊٿ3(���@F�2�4@�`{IА!?�iK�#�@5�=PƊٿ3(���@F�2�4@�`{IА!?�iK�#�@5�=PƊٿ3(���@F�2�4@�`{IА!?�iK�#�@�vQ@�ٿ�(�o;��@(��V4@]��Ȑ!?a���@�vQ@�ٿ�(�o;��@(��V4@]��Ȑ!?a���@�vQ@�ٿ�(�o;��@(��V4@]��Ȑ!?a���@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@�)bW��ٿd�.9��@��VՈ4@�����!?�k�F;��@3b���ٿfT�QcU�@�gɕ4@C��g
�!?�G��Y�@B<ބٿ���H��@���:4@*�=�!?�]RLD�@B<ބٿ���H��@���:4@*�=�!?�]RLD�@B<ބٿ���H��@���:4@*�=�!?�]RLD�@B<ބٿ���H��@���:4@*�=�!?�]RLD�@B<ބٿ���H��@���:4@*�=�!?�]RLD�@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@ID�&��ٿ*~7��@���k?4@�Y] ��!?{�=ސ��@AtT��ٿ��QRQ �@�l�4@�C����!?�R";��@AtT��ٿ��QRQ �@�l�4@�C����!?�R";��@AtT��ٿ��QRQ �@�l�4@�C����!?�R";��@AtT��ٿ��QRQ �@�l�4@�C����!?�R";��@J�R��ٿ��U;��@����4@�U���!?S1mv[��@J�R��ٿ��U;��@����4@�U���!?S1mv[��@�-i�݃ٿ ��7��@l��E	4@#Z@=��!?+Sc����@�-i�݃ٿ ��7��@l��E	4@#Z@=��!?+Sc����@�-i�݃ٿ ��7��@l��E	4@#Z@=��!?+Sc����@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@��Q��ٿ�%§�@����E4@9R}�ؐ!?p�Z_K�@&n�%#�ٿ �l*9�@	�fU4@��{Oې!?�0��v�@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�qaF�ٿ���k��@qw�+d4@��p5��!?�s����@�9˂ٿ<����@͵��"4@3����!?�.S��@�9˂ٿ<����@͵��"4@3����!?�.S��@�9˂ٿ<����@͵��"4@3����!?�.S��@�9˂ٿ<����@͵��"4@3����!?�.S��@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@z��ۜ�ٿ4��Z�@Gάt�4@�'�5ϐ!?dP	LT�@TR��Ѓٿ:c�.C�@]&�	4@>���А!?���B&��@TR��Ѓٿ:c�.C�@]&�	4@>���А!?���B&��@TR��Ѓٿ:c�.C�@]&�	4@>���А!?���B&��@�l@��ٿ�N���@����4@[E�\x�!?�7���@�l@��ٿ�N���@����4@[E�\x�!?�7���@�l@��ٿ�N���@����4@[E�\x�!?�7���@�l@��ٿ�N���@����4@[E�\x�!?�7���@�#�H�~ٿ9��&�2�@�|�
4@M(��ʐ!?}� }�@q%��5�ٿ�[ ��7�@XϮU�	4@������!?M�`/�w�@q%��5�ٿ�[ ��7�@XϮU�	4@������!?M�`/�w�@���& ~ٿ�B�O�@����	4@�#Ő!?hS��@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@7��ź~ٿ�V�/P6�@��� 4@j68�!?[Hy�`y�@��h�9�ٿqa�Mo��@��C:4@vr����!?Cd¶+�@��D���ٿ�OB1��@��Y4@���ε�!?�����@��D���ٿ�OB1��@��Y4@���ε�!?�����@��D���ٿ�OB1��@��Y4@���ε�!?�����@��D���ٿ�OB1��@��Y4@���ε�!?�����@��D���ٿ�OB1��@��Y4@���ε�!?�����@��D���ٿ�OB1��@��Y4@���ε�!?�����@�n�_�ٿF8�:w��@ƺ`{s4@��)��!?8�{����@�n�_�ٿF8�:w��@ƺ`{s4@��)��!?8�{����@�n�_�ٿF8�:w��@ƺ`{s4@��)��!?8�{����@�n�_�ٿF8�:w��@ƺ`{s4@��)��!?8�{����@�n�_�ٿF8�:w��@ƺ`{s4@��)��!?8�{����@Z��ߌٿL
����@b���4@�Ns���!?�[����@Z��ߌٿL
����@b���4@�Ns���!?�[����@Z��ߌٿL
����@b���4@�Ns���!?�[����@8��jԏٿ@�ڳ���@h��24@;N����!?�P�E���@8��jԏٿ@�ڳ���@h��24@;N����!?�P�E���@��&���ٿit{����@�F��g�3@3��聐!?���q���@��&���ٿit{����@�F��g�3@3��聐!?���q���@.zjȅٿ�$���@~�I!d4@�^6��!?#�=) �@.zjȅٿ�$���@~�I!d4@�^6��!?#�=) �@�v�z�ٿ�v"�@�-&f�	4@4��Yǐ!?��b"1��@���ٿ����.�@���e4@�UՐ!?0�+I���@���ٿ����.�@���e4@�UՐ!?0�+I���@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@�4w\�ٿKoU�9l�@�C�4@_�W��!?<<��B�@����0�ٿ�R��"��@9�ɴ�4@F����!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@����ٿ�����@��V��4@�hmݐ!?������@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�)c��ٿ8I1���@$�)��4@���!?��1ǣ�@�Q���ٿ�#�����@�~i4@%A#^ސ!?��0N0��@"�8�ٿ���w0�@��c�e4@���c��!? �{a��@"�8�ٿ���w0�@��c�e4@���c��!? �{a��@;�v���ٿq�(���@m�>�4@����!?���
x��@;�v���ٿq�(���@m�>�4@����!?���
x��@;�v���ٿq�(���@m�>�4@����!?���
x��@;�v���ٿq�(���@m�>�4@����!?���
x��@�λ�#�ٿ@��AI��@�'���4@|�󜄐!?�&����@|�dN��ٿ��M�p��@�;/3�4@_�\�\�!?}����@|�dN��ٿ��M�p��@�;/3�4@_�\�\�!?}����@|�dN��ٿ��M�p��@�;/3�4@_�\�\�!?}����@�+f��ٿ�ۏ��z�@���k4@ۗ�^��!?S�-�9�@�+f��ٿ�ۏ��z�@���k4@ۗ�^��!?S�-�9�@�+f��ٿ�ۏ��z�@���k4@ۗ�^��!?S�-�9�@�+f��ٿ�ۏ��z�@���k4@ۗ�^��!?S�-�9�@�+f��ٿ�ۏ��z�@���k4@ۗ�^��!?S�-�9�@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@�(�pE�ٿ$�*���@�Y�4@+ӆu��!?8�'���@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@x`ڤ��ٿ,G��1�@~[�4@��OLÐ!?	,Źb��@e��sH�ٿ1��A��@L��vq4@���,��!?q�K���@e��sH�ٿ1��A��@L��vq4@���,��!?q�K���@�7b�ٿ���̾$�@����04@��˽�!?���E��@�7b�ٿ���̾$�@����04@��˽�!?���E��@�7b�ٿ���̾$�@����04@��˽�!?���E��@�@�]�ٿ�M�����@�n��4@��O�!?��~���@�@�]�ٿ�M�����@�n��4@��O�!?��~���@�@�]�ٿ�M�����@�n��4@��O�!?��~���@�@�]�ٿ�M�����@�n��4@��O�!?��~���@�=��ٿ��
�#�@��c��4@6�8��!?���d��@�~��ٿ�ߝ�V�@���*4@��N��!?����[�@�~��ٿ�ߝ�V�@���*4@��N��!?����[�@�~��ٿ�ߝ�V�@���*4@��N��!?����[�@�~��ٿ�ߝ�V�@���*4@��N��!?����[�@�3����ٿ����Y�@ hl�?4@xR�~��!?��:��W�@�3����ٿ����Y�@ hl�?4@xR�~��!?��:��W�@2����ٿJ���C��@���4@�_�h��!?���J��@2����ٿJ���C��@���4@�_�h��!?���J��@2����ٿJ���C��@���4@�_�h��!?���J��@2����ٿJ���C��@���4@�_�h��!?���J��@�o��ނٿ@�����@QY��	4@��΄�!?�Uƻ^��@�o��ނٿ@�����@QY��	4@��΄�!?�Uƻ^��@�o��ނٿ@�����@QY��	4@��΄�!?�Uƻ^��@�o��ނٿ@�����@QY��	4@��΄�!?�Uƻ^��@�o��ނٿ@�����@QY��	4@��΄�!?�Uƻ^��@�u�' �ٿ|_��en�@7~�
/
4@�Fs8��!?�|H�E�@�u�' �ٿ|_��en�@7~�
/
4@�Fs8��!?�|H�E�@�*�XL�ٿ̻B���@�c�	4@}9ږސ!?MdNl��@@��{ٿ�l�^���@-���4@���ؐ!?tq�'�@@��{ٿ�l�^���@-���4@���ؐ!?tq�'�@@��{ٿ�l�^���@-���4@���ؐ!?tq�'�@@��{ٿ�l�^���@-���4@���ؐ!?tq�'�@���iلٿ�
RѪB�@em�s�4@3��xĐ!?�3�h�@���iلٿ�
RѪB�@em�s�4@3��xĐ!?�3�h�@���iلٿ�
RѪB�@em�s�4@3��xĐ!?�3�h�@���iلٿ�
RѪB�@em�s�4@3��xĐ!?�3�h�@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@��сDٿ�`�e���@U!d'4@�b8R �!?��?zY��@3iWVWٿhӭ�Q�@��m��4@v� =�!?l��?H�@3iWVWٿhӭ�Q�@��m��4@v� =�!?l��?H�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@���x(ٿ+��G�@�f�X4@�z�sː!?u�:)o�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@}�(��~ٿ��4��@�n��4@e��ei�!?=B���c�@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@�DzI �ٿ+�����@��e�C4@'�͋�!?h ����@]g��ٿ�kڈ���@ճ9�s4@�EAᑐ!?O�v�x��@]g��ٿ�kڈ���@ճ9�s4@�EAᑐ!?O�v�x��@]g��ٿ�kڈ���@ճ9�s4@�EAᑐ!?O�v�x��@��#�ٿ
�J�<�@b��m�4@�T�	�!?f���@��#�ٿ
�J�<�@b��m�4@�T�	�!?f���@��#�ٿ
�J�<�@b��m�4@�T�	�!?f���@��#�ٿ
�J�<�@b��m�4@�T�	�!?f���@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@|&�/X�ٿ�@�8�@a���A4@DDP�4�!?����nx�@��h��ٿ)�M,�^�@),�4@>���Z�!?)��4�@��h��ٿ)�M,�^�@),�4@>���Z�!?)��4�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@U{
jօٿ`���*�@>�`�
4@,C�6��!?���N�E�@�c�y�ٿBv%M���@7E�T4@��o�ؐ!?58TW)��@�c�y�ٿBv%M���@7E�T4@��o�ؐ!?58TW)��@�c�y�ٿBv%M���@7E�T4@��o�ؐ!?58TW)��@�c�y�ٿBv%M���@7E�T4@��o�ؐ!?58TW)��@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@��
P҆ٿ����QZ�@�ے)	4@�z��!?;�	�@�H�g��ٿ,߉���@�^��a4@Z��!?�f?��@�H�g��ٿ,߉���@�^��a4@Z��!?�f?��@�H�g��ٿ,߉���@�^��a4@Z��!?�f?��@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@f�!�Áٿ�.yf��@&a��4@�ZH���!?�#�Jn\�@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@GL]�ٿ�<#�'��@��_�4@c��>Ր!?D�~��@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@*��ٿ�&�
�@{�>4@����/�!?�i����@W���ٿ1?�i( �@u��&4@v��婐!?q�ȴ?
�@�� ˑٿ&��^&�@{zW�4@ފ�ʬ�!?p"�@�W�@�� ˑٿ&��^&�@{zW�4@ފ�ʬ�!?p"�@�W�@�� ˑٿ&��^&�@{zW�4@ފ�ʬ�!?p"�@�W�@�� ˑٿ&��^&�@{zW�4@ފ�ʬ�!?p"�@�W�@�� ˑٿ&��^&�@{zW�4@ފ�ʬ�!?p"�@�W�@�X��ٿ"�-&o��@���4@�zJ#��!?��C�:�@�X��ٿ"�-&o��@���4@�zJ#��!?��C�:�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@��-�ٿ�ؑ���@}���
4@n!�Xǐ!?<�2F�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@M�_t��ٿ&R <�A�@�\��V4@.�~�!?�2Nߣ�@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@���Ѝٿ��)�l(�@�9��(4@����!?R0\B	��@N����ٿ�PI:!��@�`$�
4@Z��0�!?��Z؟�@N����ٿ�PI:!��@�`$�
4@Z��0�!?��Z؟�@N����ٿ�PI:!��@�`$�
4@Z��0�!?��Z؟�@N����ٿ�PI:!��@�`$�
4@Z��0�!?��Z؟�@+�M�ٿL%�'��@�n�94@V˧�%�!?���#��@+�M�ٿL%�'��@�n�94@V˧�%�!?���#��@+�M�ٿL%�'��@�n�94@V˧�%�!?���#��@+�M�ٿL%�'��@�n�94@V˧�%�!?���#��@�P)!�ٿha��Q�@�q6�
4@P4SȺ�!?�6'�~��@�P)!�ٿha��Q�@�q6�
4@P4SȺ�!?�6'�~��@�P)!�ٿha��Q�@�q6�
4@P4SȺ�!?�6'�~��@Q��"G�ٿ�<�V�@��	��4@N�戀!?����T�@Q��"G�ٿ�<�V�@��	��4@N�戀!?����T�@���J�ٿĨ�O�L�@$kt4@�j�$,�!?tc�yc�@���J�ٿĨ�O�L�@$kt4@�j�$,�!?tc�yc�@���J�ٿĨ�O�L�@$kt4@�j�$,�!?tc�yc�@���J�ٿĨ�O�L�@$kt4@�j�$,�!?tc�yc�@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�d����ٿH7"�@��	�T4@ݹx�%�!? 񎪛��@�쟅ٿ�e	�
�@eg�Ѣ4@�%��ِ!?�	o���@�쟅ٿ�e	�
�@eg�Ѣ4@�%��ِ!?�	o���@�쟅ٿ�e	�
�@eg�Ѣ4@�%��ِ!?�	o���@�쟅ٿ�e	�
�@eg�Ѣ4@�%��ِ!?�	o���@�쟅ٿ�e	�
�@eg�Ѣ4@�%��ِ!?�	o���@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@'���ٿ� �g��@����4@iqHҚ�!?N1�s��@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@�}�C�ٿ�,(�C�@Rŧ84@E��:��!?�W`7�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@K�z�"�ٿ��I=*�@^.�w�4@Ξ[,~�!?w�!�"�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�0���ٿ���|P�@����4@/I^d�!?..��K�@�����}ٿsa´f��@��5��4@��m홐!?��OG'�@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@��dL��ٿ��W$��@�t��4@�#Ş�!?��F��@�b���ٿ+����@&/�<�4@x��ew�!?�Vƹ`��@�b���ٿ+����@&/�<�4@x��ew�!?�Vƹ`��@��	�ٿ�ŔYF��@b�-�!4@^ـ���!?�θ~���@��	�ٿ�ŔYF��@b�-�!4@^ـ���!?�θ~���@��	�ٿ�ŔYF��@b�-�!4@^ـ���!?�θ~���@��	�ٿ�ŔYF��@b�-�!4@^ـ���!?�θ~���@��<ԇٿH�Y�)_�@�2�;�4@��ᾐ!?�a�곖�@��<ԇٿH�Y�)_�@�2�;�4@��ᾐ!?�a�곖�@��<ԇٿH�Y�)_�@�2�;�4@��ᾐ!?�a�곖�@��<ԇٿH�Y�)_�@�2�;�4@��ᾐ!?�a�곖�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@� 3lk�ٿ��ufV��@kh}��4@���!?�t�6�r�@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@w	���ٿs.5-��@u�#`�4@�K�=��!?�u>���@�n$�1�ٿ���%4�@{fN�.4@�Q�ǐ!?0D�6��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@�;{��ٿ3WO�"+�@�u��g4@ת����!?�H̱��@����ٿT��.$�@`���&4@�G6��!?�2�#�@����ٿT��.$�@`���&4@�G6��!?�2�#�@����ٿT��.$�@`���&4@�G6��!?�2�#�@����ٿT��.$�@`���&4@�G6��!?�2�#�@����ٿT��.$�@`���&4@�G6��!?�2�#�@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@������ٿ8d
���@�y_4@{*�hK�!?2�����@�7c)c�ٿ?������@���oY4@y�*�Ԑ!? �a�3g�@�A��Ɇٿ�q���i�@4�>F4@���H��!?�"�f���@'*?-�ٿ��oۘ��@K�K�O4@s)��!?�Kb s�@'*?-�ٿ��oۘ��@K�K�O4@s)��!?�Kb s�@'*?-�ٿ��oۘ��@K�K�O4@s)��!?�Kb s�@&�-ۆٿQn���@�'o��4@ďw���!?q�x���@���~ٿ^���=�@�����	4@�ʺ��!?�u��)�@���~ٿ^���=�@�����	4@�ʺ��!?�u��)�@���~ٿ^���=�@�����	4@�ʺ��!?�u��)�@���~ٿ^���=�@�����	4@�ʺ��!?�u��)�@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@��<﯀ٿэ8�?�@�c��4@�IJ�ܐ!?�j���@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@���ʄٿ��9E�X�@z���E4@��i��!?��,<��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@N`c�ٿd������@��O4@~�!��!?/\�=��@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@#<g��ٿ��ka�a�@q�&�"4@^�ϐ!?Y��=~.�@�F��ٿh��j���@���K4@ǘSՐ!?��ڞ�@�F��ٿh��j���@���K4@ǘSՐ!?��ڞ�@�F��ٿh��j���@���K4@ǘSՐ!?��ڞ�@�F��ٿh��j���@���K4@ǘSՐ!?��ڞ�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@ou��ٿ��ad���@Ψ��d4@�L��ߐ!?�FB>m|�@�3flM�ٿ�8=�5�@�*�w4@��<�!?�UViG�@�3flM�ٿ�8=�5�@�*�w4@��<�!?�UViG�@�3flM�ٿ�8=�5�@�*�w4@��<�!?�UViG�@�0]r�ٿ.}��@B���4@dq�!?$X��$�@ͬ�߰�ٿ�o���=�@ޛ�i�4@?��(�!?�Z��]�@ͬ�߰�ٿ�o���=�@ޛ�i�4@?��(�!?�Z��]�@ͬ�߰�ٿ�o���=�@ޛ�i�4@?��(�!?�Z��]�@�4@ۇٿBH�yK4�@���"4@�G
|��!?ek?�6��@�4@ۇٿBH�yK4�@���"4@�G
|��!?ek?�6��@�4@ۇٿBH�yK4�@���"4@�G
|��!?ek?�6��@�4@ۇٿBH�yK4�@���"4@�G
|��!?ek?�6��@���L�ٿ��|x�q�@���2�4@*�ѽ�!?�
rbo�@���L�ٿ��|x�q�@���2�4@*�ѽ�!?�
rbo�@���L�ٿ��|x�q�@���2�4@*�ѽ�!?�
rbo�@���L�ٿ��|x�q�@���2�4@*�ѽ�!?�
rbo�@3&ϼ�ٿ����C�@hI�NL4@�"��!?b�n�;��@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@m��*��ٿM���$�@�>��4@��(�ڐ!?�[#�y�@�c�o�ٿsPz���@Ǌ�<�4@'fҍ��!?��S ���@lmD��ٿ����	��@���474@ ��d�!?�aH�<��@lmD��ٿ����	��@���474@ ��d�!?�aH�<��@lmD��ٿ����	��@���474@ ��d�!?�aH�<��@lmD��ٿ����	��@���474@ ��d�!?�aH�<��@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@T�ô��ٿp��Rx�@�>��4@�X�A�!?`�M�[�@��;�ٿV�c5~��@9��4@�C6�m�!?Y��+��@��;�ٿV�c5~��@9��4@�C6�m�!?Y��+��@��;�ٿV�c5~��@9��4@�C6�m�!?Y��+��@��Z��ٿ�瀆��@SNg�4@�VdJ�!?J�	 
��@��Z��ٿ�瀆��@SNg�4@�VdJ�!?J�	 
��@1�����ٿJB�K"��@��?��4@��lꖐ!?����[-�@Wz�FS�ٿ�w|�b�@p�hm4@ԊD��!?w���I�@Wz�FS�ٿ�w|�b�@p�hm4@ԊD��!?w���I�@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@)�wA}ٿ�)k��@tX�4@�W��Ր!?p��t��@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@i��ui�ٿ�Wl2T�@_�B�'4@/X�'��!?4��]:�@�5+C�ٿ<!^�@��@���h�3@�C����!?r;d�w�@�_}�ٿ�K��9�@	���3@Q��Đ!?)�H��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@�[v�\�ٿPEΔx�@ib��S4@�]"�ǐ!?6��#��@HMv(��ٿ�`���@�U��4@���.Ő!?yc���@HMv(��ٿ�`���@�U��4@���.Ő!?yc���@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@���A/�ٿ��2�o��@�J�t�4@s<#��!?/P'�՚�@�c�ٿd�NG��@r0(��	4@'�lE��!?����}�@�c�ٿd�NG��@r0(��	4@'�lE��!?����}�@�c�ٿd�NG��@r0(��	4@'�lE��!?����}�@�-�Áٿ�V����@qׁ��4@ؿ[wŐ!?Ez���@�-�Áٿ�V����@qׁ��4@ؿ[wŐ!?Ez���@I ��ٿ����@j�@<�)��4@�� ��!?T�J^�R�@I ��ٿ����@j�@<�)��4@�� ��!?T�J^�R�@I ��ٿ����@j�@<�)��4@�� ��!?T�J^�R�@I ��ٿ����@j�@<�)��4@�� ��!?T�J^�R�@I ��ٿ����@j�@<�)��4@�� ��!?T�J^�R�@�!P��ٿͤH/��@h$s	4@�x�^��!?������@϶��ыٿ���G��@�F�wE4@TI��!?���$4��@϶��ыٿ���G��@�F�wE4@TI��!?���$4��@϶��ыٿ���G��@�F�wE4@TI��!?���$4��@ !�ٿUV�����@����>4@ZƮ�2�!?�p��:7�@ !�ٿUV�����@����>4@ZƮ�2�!?�p��:7�@ !�ٿUV�����@����>4@ZƮ�2�!?�p��:7�@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@�sAU˃ٿXS`��@@����4@݄5�s�!?��.��@��?,�ٿ�Q�7t�@yQ6�4@�)�Ú�!?uE���N�@��?,�ٿ�Q�7t�@yQ6�4@�)�Ú�!?uE���N�@��?,�ٿ�Q�7t�@yQ6�4@�)�Ú�!?uE���N�@��?,�ٿ�Q�7t�@yQ6�4@�)�Ú�!?uE���N�@��?,�ٿ�Q�7t�@yQ6�4@�)�Ú�!?uE���N�@�����ٿ�6W����@�6Ʊ4@gSI���!?Q��	z��@�����ٿ�6W����@�6Ʊ4@gSI���!?Q��	z��@�e�h��ٿ��`�A.�@�]� 4@I�yՐ!?_�7�u2�@�e�h��ٿ��`�A.�@�]� 4@I�yՐ!?_�7�u2�@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@\@B�	�ٿ��� ��@2�!�/4@[v^`N�!?.u�����@�T8�E�ٿuj�&�@�w��4@��_�!?ĸ��N�@�T8�E�ٿuj�&�@�w��4@��_�!?ĸ��N�@�T8�E�ٿuj�&�@�w��4@��_�!?ĸ��N�@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@�n>I�ٿb"Q�A�@�*4@���!?l��}��@��F�ٿ%����3�@{Bm�4@_M���!?N,sIS
�@��F�ٿ%����3�@{Bm�4@_M���!?N,sIS
�@��F�ٿ%����3�@{Bm�4@_M���!?N,sIS
�@��F�ٿ%����3�@{Bm�4@_M���!?N,sIS
�@��F�ٿ%����3�@{Bm�4@_M���!?N,sIS
�@>xŏٿg��
���@�,�)n 4@aÞx��!?-K�]:��@>xŏٿg��
���@�,�)n 4@aÞx��!?-K�]:��@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�9�A��ٿ{������@ �.:�4@���Ԑ!?ڏ�V�P�@�����ٿ�Y�h(��@�
aX;4@�x����!?p@�#�S�@�����ٿ�Y�h(��@�
aX;4@�x����!?p@�#�S�@FzP���ٿ��F���@f�=·4@�0`]`�!?އY����@FzP���ٿ��F���@f�=·4@�0`]`�!?އY����@�_�	�ٿ��h�iJ�@EO�	4@���a��!?ct]zU��@X�6 z�ٿ�)�W��@7ht��4@F7��!?��i �@X�6 z�ٿ�)�W��@7ht��4@F7��!?��i �@X�6 z�ٿ�)�W��@7ht��4@F7��!?��i �@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@M T��ٿ�(��0�@�[:4@b����!?����z��@����}}ٿ���`�@�@I2f��4@��Ր!?�9K]�.�@����}}ٿ���`�@�@I2f��4@��Ր!?�9K]�.�@����}}ٿ���`�@�@I2f��4@��Ր!?�9K]�.�@����}}ٿ���`�@�@I2f��4@��Ր!?�9K]�.�@����}}ٿ���`�@�@I2f��4@��Ր!?�9K]�.�@#g��I�ٿW��5��@����b4@�יyw�!?N��VUu�@#g��I�ٿW��5��@����b4@�יyw�!?N��VUu�@#g��I�ٿW��5��@����b4@�יyw�!?N��VUu�@#g��I�ٿW��5��@����b4@�יyw�!?N��VUu�@��%L�ٿs �]���@SK�[�4@�,8g�!?������@��%L�ٿs �]���@SK�[�4@�,8g�!?������@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@����ٿ�À��@��u��4@j,;�Ӑ!?�$졮f�@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@d�)�ٿ;J�^ ��@���Y	4@?<H��!?�-���@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@��͋ٿ|

�o�@�%.[�4@�[��!?$�rd��@���ЎٿP����@�=���4@r���ǐ!?�ֶ�;��@���ЎٿP����@�=���4@r���ǐ!?�ֶ�;��@���ЎٿP����@�=���4@r���ǐ!?�ֶ�;��@���ЎٿP����@�=���4@r���ǐ!?�ֶ�;��@���ЎٿP����@�=���4@r���ǐ!?�ֶ�;��@��Rٿ���V�@�@���4@i4mې!?Ns g��@��Rٿ���V�@�@���4@i4mې!?Ns g��@��Rٿ���V�@�@���4@i4mې!?Ns g��@��Rٿ���V�@�@���4@i4mې!?Ns g��@�mB�ٿ�t�@�C�44@�;�i@�!?��M>9�@�mB�ٿ�t�@�C�44@�;�i@�!?��M>9�@�E�c�ٿ�!r:�k�@��)4@a��0�!?a�����@�E�c�ٿ�!r:�k�@��)4@a��0�!?a�����@�E�c�ٿ�!r:�k�@��)4@a��0�!?a�����@�u�v��ٿR�6�>��@d+$j4@B���6�!?{k* ^��@�u�v��ٿR�6�>��@d+$j4@B���6�!?{k* ^��@��b>��ٿn+�ìd�@%7� � 4@�c�!?��@��b>��ٿn+�ìd�@%7� � 4@�c�!?��@��b>��ٿn+�ìd�@%7� � 4@�c�!?��@��b>��ٿn+�ìd�@%7� � 4@�c�!?��@���z�ٿu�X�e=�@Z8^. 4@H�#�!?��Z�9�@���z�ٿu�X�e=�@Z8^. 4@H�#�!?��Z�9�@M~r���ٿ`Vk��%�@ܛ�_L4@��Ei��!?�.4�T��@�gH��ٿbs��@�����4@��3L��!?�=j��@�gH��ٿbs��@�����4@��3L��!?�=j��@7#"�6�ٿ��9-��@$sG�4@C��!?�$Y}���@7#"�6�ٿ��9-��@$sG�4@C��!?�$Y}���@7#"�6�ٿ��9-��@$sG�4@C��!?�$Y}���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@��M�ٿ[8ѷ,��@���4@q%���!?�#z���@�͒̍ٿ�2uo=�@)�84@N����!?�/�~]�@��_B��ٿE�g$��@m,d�4@�l���!?ZM�����@��_B��ٿE�g$��@m,d�4@�l���!?ZM�����@��_B��ٿE�g$��@m,d�4@�l���!?ZM�����@��_B��ٿE�g$��@m,d�4@�l���!?ZM�����@��_B��ٿE�g$��@m,d�4@�l���!?ZM�����@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@��p���ٿx!���@"�l�4@7�@j�!?���Trx�@�c.(�ٿ5q��]��@/���4@�r�Ѐ�!?d���m�@��Nύ�ٿI ����@��I�4@�bVS�!?�D:�y�@��Nύ�ٿI ����@��I�4@�bVS�!?�D:�y�@��Nύ�ٿI ����@��I�4@�bVS�!?�D:�y�@��Nύ�ٿI ����@��I�4@�bVS�!?�D:�y�@��Nύ�ٿI ����@��I�4@�bVS�!?�D:�y�@��C��ٿ_�ϔ�@KMܼ�4@m
��7�!?qo�q�@����ٿ���i8�@�7�4@0[�7�!?2+A$���@����ٿ���i8�@�7�4@0[�7�!?2+A$���@	2���ٿ��v�C�@�z�׿4@�&{!�!?�B��|��@	2���ٿ��v�C�@�z�׿4@�&{!�!?�B��|��@	2���ٿ��v�C�@�z�׿4@�&{!�!?�B��|��@*��V��ٿy����8�@�э��4@Q\p��!?���O�@�t��ٿ��X���@�h�?4@�����!?����z�@�t��ٿ��X���@�h�?4@�����!?����z�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�&򸶋ٿ��L�2I�@��ԬN4@V����!?} }:g�@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@�н��ٿ!"ׂM�@�̆4@�2{k��!?����@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@G�:W~�ٿ@�9��@�(^�4@�X 	��!?,���_�@2$��҉ٿ��D_m�@X����4@`?���!?M����]�@2$��҉ٿ��D_m�@X����4@`?���!?M����]�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@�D�2��ٿ�	����@�:p�4@{�4��!?�@�m�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@Fb5.2�ٿ�[����@��8v4@+NtԐ!?��J�@j�H.��ٿ0è�n��@�C�2�4@}����!?�v�t�@j�H.��ٿ0è�n��@�C�2�4@}����!?�v�t�@j�H.��ٿ0è�n��@�C�2�4@}����!?�v�t�@�B���ٿ��-��@c��]4@��Ő!?BkB���@�B���ٿ��-��@c��]4@��Ő!?BkB���@�B���ٿ��-��@c��]4@��Ő!?BkB���@�M��U�ٿ��~���@et�r4@�}�ى�!?�2��@�M��U�ٿ��~���@et�r4@�}�ى�!?�2��@o�Wo�ٿ��=PaZ�@ȋ诘4@��E賐!?�bWR~1�@o�Wo�ٿ��=PaZ�@ȋ诘4@��E賐!?�bWR~1�@o�Wo�ٿ��=PaZ�@ȋ诘4@��E賐!?�bWR~1�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�R:ٿQ��+���@�$�Q4@��c�M�!?�W]QSv�@�}{i-�ٿ
R�D���@�˗��4@_��
>�!?%�PgL��@R�!S�ٿ����=�@�x�4@8����!?�;�7
^�@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@,x�	}�ٿx���O�@qu�`�4@����!?բ-t��@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�3y��ٿ��F�t�@��4@�5��!?�x�� �@�6���ٿ��(@��@^�W[� 4@�E���!?*�eT�@d�R6�ٿu��A��@2 4@CC�đ�!?vs��.�@d�R6�ٿu��A��@2 4@CC�đ�!?vs��.�@d�R6�ٿu��A��@2 4@CC�đ�!?vs��.�@d�R6�ٿu��A��@2 4@CC�đ�!?vs��.�@d�R6�ٿu��A��@2 4@CC�đ�!?vs��.�@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@e�(�ٿ��A����@
�>�4@,�~��!?�Vu�2��@n/n�:�ٿ���[�@�,1��4@�p���!?Tx9{�*�@�T��]�ٿ<����@8XaIR4@��ڲ��!?�n�6Y�@��q��ٿZ��N$@�@���r4@u�O�Ȑ!?G��~�@��q��ٿZ��N$@�@���r4@u�O�Ȑ!?G��~�@���� �ٿ6V}��&�@͎�+4@�%�bb�!?��P��@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@;��TT�ٿŦ�����@l]O4@�'|⦐!?>6�i�~�@U|g�ٿdqe'��@�_��4@��V��!?�IO�s�@U|g�ٿdqe'��@�_��4@��V��!?�IO�s�@U|g�ٿdqe'��@�_��4@��V��!?�IO�s�@�ϟ���ٿ'�Xg��@�����3@�3�c�!?Sϛi���@�ϟ���ٿ'�Xg��@�����3@�3�c�!?Sϛi���@�ϟ���ٿ'�Xg��@�����3@�3�c�!?Sϛi���@�O'�M�ٿ|�=n�@�\/4@8�]��!?�������@�O'�M�ٿ|�=n�@�\/4@8�]��!?�������@�O'�M�ٿ|�=n�@�\/4@8�]��!?�������@I�ߊٿ�O6���@C|N�4@���o��!?���q:��@I�ߊٿ�O6���@C|N�4@���o��!?���q:��@I�ߊٿ�O6���@C|N�4@���o��!?���q:��@I�ߊٿ�O6���@C|N�4@���o��!?���q:��@I�ߊٿ�O6���@C|N�4@���o��!?���q:��@D�[B�ٿyc^��@�j���4@`�~��!?��*.�@D�[B�ٿyc^��@�j���4@`�~��!?��*.�@��Vq��ٿR�x��@��1Qi4@�����!?�w���P�@��Vq��ٿR�x��@��1Qi4@�����!?�w���P�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@S�ׇ��ٿqh'�0�@\�4@�6���!?��;��c�@v�p��ٿ���	��@?�YK>4@���!?�R{����@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@�>�Ř�ٿd� I��@1�n
,4@�Wf,�!?;�<Fm��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@]�.k�ٿ���5/�@�|��4@W_?�!?�JK��@$��N�ٿ+emT���@mu�/�4@�ѠC�!?�B��;l�@m}��ٿK��Rc��@����� 4@�;'�!?���ۃ�@m}��ٿK��Rc��@����� 4@�;'�!?���ۃ�@m}��ٿK��Rc��@����� 4@�;'�!?���ۃ�@m}��ٿK��Rc��@����� 4@�;'�!?���ۃ�@m}��ٿK��Rc��@����� 4@�;'�!?���ۃ�@FG����ٿYyx���@<���3@	q�? �!?�n5N��@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@�X�ٿ;�W���@˓8�3@$
���!?����I-�@��/��ٿO0����@���gZ4@�Q���!?�?����@��/��ٿO0����@���gZ4@�Q���!?�?����@��/��ٿO0����@���gZ4@�Q���!?�?����@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@ �E��ٿ�b9���@�dE� 4@D"`k��!?!o`W���@��c�{ٿ�6�|��@���4@>���!?bA���@��c�{ٿ�6�|��@���4@>���!?bA���@ZI���ٿ�ꬓJ��@]\�4@:�9��!?��j]���@ZI���ٿ�ꬓJ��@]\�4@:�9��!?��j]���@ZI���ٿ�ꬓJ��@]\�4@:�9��!?��j]���@ZI���ٿ�ꬓJ��@]\�4@:�9��!?��j]���@ZI���ٿ�ꬓJ��@]\�4@:�9��!?��j]���@�[x}ٿϊ�C�j�@E�ԕ4@��볽�!?� ԧ��@�[x}ٿϊ�C�j�@E�ԕ4@��볽�!?� ԧ��@�[x}ٿϊ�C�j�@E�ԕ4@��볽�!?� ԧ��@�[x}ٿϊ�C�j�@E�ԕ4@��볽�!?� ԧ��@�鐶~ٿV�����@��LQd4@�G�*!?J�՞�@�鐶~ٿV�����@��LQd4@�G�*!?J�՞�@�鐶~ٿV�����@��LQd4@�G�*!?J�՞�@�鐶~ٿV�����@��LQd4@�G�*!?J�՞�@�鐶~ٿV�����@��LQd4@�G�*!?J�՞�@M'�⋃ٿ�{�K�@��⁊4@NAov�!?����@��ﴹ�ٿB�9>�@�t�z4@"�	�!?��F�x��@��ﴹ�ٿB�9>�@�t�z4@"�	�!?��F�x��@��ﴹ�ٿB�9>�@�t�z4@"�	�!?��F�x��@�g�֐}ٿnʛN��@]�E4@̯�L��!?3�9��z�@�9�Q�ٿ��Z1��@]C��4@@[�p�!?֭�0�!�@�9�Q�ٿ��Z1��@]C��4@@[�p�!?֭�0�!�@�9�Q�ٿ��Z1��@]C��4@@[�p�!?֭�0�!�@��@��ٿ�+M���@����4@�X�!?�4*8���@��@��ٿ�+M���@����4@�X�!?�4*8���@��@��ٿ�+M���@����4@�X�!?�4*8���@��@��ٿ�+M���@����4@�X�!?�4*8���@��@��ٿ�+M���@����4@�X�!?�4*8���@��@��ٿ�+M���@����4@�X�!?�4*8���@<�᫹�ٿ���)|�@��X��4@���Ր!?�|9`+�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@���l��ٿm�_��@IjR�4@>�Hj�!?���4^�@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@��h�v�ٿ���p�@�5��q4@�S���!?c�k���@c�bQ�ٿh|�v8�@�����4@!�����!?��S)�@c�bQ�ٿh|�v8�@�����4@!�����!?��S)�@V�Q�!�ٿd��.�n�@ۄY;�4@r�C���!?9���@V�Q�!�ٿd��.�n�@ۄY;�4@r�C���!?9���@V�Q�!�ٿd��.�n�@ۄY;�4@r�C���!?9���@V�Q�!�ٿd��.�n�@ۄY;�4@r�C���!?9���@p��n�ٿ׈��
^�@~K<H44@)&2ِ!?x<\&4��@S�~/m�ٿ��9�`�@:��X;4@�\�(��!?`wp�3��@S�~/m�ٿ��9�`�@:��X;4@�\�(��!?`wp�3��@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@B�9���ٿ�#��b�@���҃4@��L��!?7ך���@Q�(��ٿ˶6��@��Z�� 4@�)x�ϐ!?|����w�@Q�(��ٿ˶6��@��Z�� 4@�)x�ϐ!?|����w�@Q�(��ٿ˶6��@��Z�� 4@�)x�ϐ!?|����w�@��O�4�ٿx�S�a�@M
�l4@K�!>$�!?.쏂 ��@�>g�ٿz5��YQ�@E�qUD4@�a��ې!?���HNe�@�>g�ٿz5��YQ�@E�qUD4@�a��ې!?���HNe�@�>g�ٿz5��YQ�@E�qUD4@�a��ې!?���HNe�@�>g�ٿz5��YQ�@E�qUD4@�a��ې!?���HNe�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�/詃ٿ���먻�@�).4@}Ot.��!?dJ��e�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@�G���ٿ��a��@�E���4@#�ك��!?��XaY�@��F��ٿxOC�Xz�@�aU�4@��H�ː!?�u���<�@��F��ٿxOC�Xz�@�aU�4@��H�ː!?�u���<�@��F��ٿxOC�Xz�@�aU�4@��H�ː!?�u���<�@2�JqP�ٿaE��#�@k��R4@�1$��!?�
���E�@�rF.�|ٿ��"�,�@nD��4@S\�W��!?-�����@�rF.�|ٿ��"�,�@nD��4@S\�W��!?-�����@�rF.�|ٿ��"�,�@nD��4@S\�W��!?-�����@�rF.�|ٿ��"�,�@nD��4@S\�W��!?-�����@�rF.�|ٿ��"�,�@nD��4@S\�W��!?-�����@3A`\!�ٿ����=P�@�	m�4@�'a�!?�d0����@f�8�v�ٿl�0��}�@K�y,4@��5#{�!?90�д��@f�8�v�ٿl�0��}�@K�y,4@��5#{�!?90�д��@�Qܙ��ٿ��l� ��@*[��4@ٚ�tn�!?	��Ob�@�Qܙ��ٿ��l� ��@*[��4@ٚ�tn�!?	��Ob�@TT0��ٿ5�����@� @4@�d&�x�!?yȂ�Vj�@TT0��ٿ5�����@� @4@�d&�x�!?yȂ�Vj�@TT0��ٿ5�����@� @4@�d&�x�!?yȂ�Vj�@TT0��ٿ5�����@� @4@�d&�x�!?yȂ�Vj�@TT0��ٿ5�����@� @4@�d&�x�!?yȂ�Vj�@�~��rٿ��"s7o�@���}4@F8����!??V�_��@�~��rٿ��"s7o�@���}4@F8����!??V�_��@,�'g�ٿ��x����@S�k4@��K��!?�x�A��@,�'g�ٿ��x����@S�k4@��K��!?�x�A��@��u�A�ٿ\���s��@ǆ�e:4@�e��!?ufWE��@��u�A�ٿ\���s��@ǆ�e:4@�e��!?ufWE��@��u�A�ٿ\���s��@ǆ�e:4@�e��!?ufWE��@��u�A�ٿ\���s��@ǆ�e:4@�e��!?ufWE��@��u�A�ٿ\���s��@ǆ�e:4@�e��!?ufWE��@y��:�ٿ�+V�n�@�
v�4@4���Ð!?*:
��@y��:�ٿ�+V�n�@�
v�4@4���Ð!?*:
��@y��:�ٿ�+V�n�@�
v�4@4���Ð!?*:
��@y��:�ٿ�+V�n�@�
v�4@4���Ð!?*:
��@y��:�ٿ�+V�n�@�
v�4@4���Ð!?*:
��@T& =d�ٿB��Y��@eKVb4@~�~�!?[7���@T& =d�ٿB��Y��@eKVb4@~�~�!?[7���@h��_I�ٿ:[Q̐F�@�.ٹ4@k;����!?��3���@h��_I�ٿ:[Q̐F�@�.ٹ4@k;����!?��3���@h��_I�ٿ:[Q̐F�@�.ٹ4@k;����!?��3���@h��_I�ٿ:[Q̐F�@�.ٹ4@k;����!?��3���@h��_I�ٿ:[Q̐F�@�.ٹ4@k;����!?��3���@�V	�ٿ
�����@�,;S�4@����!?�h���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@�J?�ٿĝ�n�@�;�C4@O�	g�!?.�M���@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��}/�ٿ�&�V��@�&SB�4@Â��!?Ǵ�o�8�@��2%�ٿ�H��%Q�@�����4@1
ӟk�!?�9���8�@��2%�ٿ�H��%Q�@�����4@1
ӟk�!?�9���8�@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@�y�Gp�ٿ�:��W�@�d��4@�@���!?�pU���@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@e�)��ٿ��|
ͫ�@���w4@�|����!?V�r�?�@�&�B�ٿ���ؕ��@\���4@z*Y��!?�>�]/�@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@��AH�ٿV���@��Ǣ\4@J�𨿐!?"M^l��@�U�$�ٿ�\>�t�@��{�4@=c��!?b =ID�@�U�$�ٿ�\>�t�@��{�4@=c��!?b =ID�@�
��\�ٿ�4X����@{4��4@]h�Κ�!?%�L���@�
��\�ٿ�4X����@{4��4@]h�Κ�!?%�L���@�
��\�ٿ�4X����@{4��4@]h�Κ�!?%�L���@�
��\�ٿ�4X����@{4��4@]h�Κ�!?%�L���@�
��\�ٿ�4X����@{4��4@]h�Κ�!?%�L���@A�y�~ٿk��頏�@h��4@�Ѥf��!?��3����@A�y�~ٿk��頏�@h��4@�Ѥf��!?��3����@A�y�~ٿk��頏�@h��4@�Ѥf��!?��3����@A�y�~ٿk��頏�@h��4@�Ѥf��!?��3����@w�S�ٿ?ձ�u�@��` 4@��$v�!?Z��5��@�c�f�ٿ�R`��@���4@�dٟ��!?݅B��m�@�c�f�ٿ�R`��@���4@�dٟ��!?݅B��m�@�c�f�ٿ�R`��@���4@�dٟ��!?݅B��m�@�c�f�ٿ�R`��@���4@�dٟ��!?݅B��m�@b1>^�ٿ�}8i���@�#Iݭ4@�O�\�!?����D�@b1>^�ٿ�}8i���@�#Iݭ4@�O�\�!?����D�@b1>^�ٿ�}8i���@�#Iݭ4@�O�\�!?����D�@b1>^�ٿ�}8i���@�#Iݭ4@�O�\�!?����D�@b1>^�ٿ�}8i���@�#Iݭ4@�O�\�!?����D�@��R���ٿ��r��@p��4@�E�Ր!?��an���@��R���ٿ��r��@p��4@�E�Ր!?��an���@3��ЇٿҺ���@�9��4@�\�7�!?�L���4�@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@L?i��ٿ�}�8� �@0��4@z
��!?���Y��@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@")m�ٿ'��J ��@e����4@A���!?���/�@�l�4�ٿ��8��@Y�?x�4@�NAߡ�!?fx$���@�l�4�ٿ��8��@Y�?x�4@�NAߡ�!?fx$���@�l�4�ٿ��8��@Y�?x�4@�NAߡ�!?fx$���@�l�4�ٿ��8��@Y�?x�4@�NAߡ�!?fx$���@�l�4�ٿ��8��@Y�?x�4@�NAߡ�!?fx$���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@i��z%�ٿ^'`ˏ�@{ Jj4@�Fmg�!?�)�f���@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@�+e�ٿ�u�*kl�@����:4@�����!?���)�Q�@=D�@=�ٿU�˒v�@zD4@ܻx�w�!?���v��@=D�@=�ٿU�˒v�@zD4@ܻx�w�!?���v��@=D�@=�ٿU�˒v�@zD4@ܻx�w�!?���v��@S���~ٿhe��@�m[�4@��Q��!?QM���I�@S���~ٿhe��@�m[�4@��Q��!?QM���I�@S���~ٿhe��@�m[�4@��Q��!?QM���I�@=W��ٿv���\�@�f	�4@C/͐!?3�j����@=W��ٿv���\�@�f	�4@C/͐!?3�j����@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@II�]�zٿF��B�E�@�a�=4@�4K��!?D������@�8�G�ٿ{Y�����@saq�d4@U�Ɨ�!?�]k#��@�8�G�ٿ{Y�����@saq�d4@U�Ɨ�!?�]k#��@��	���ٿ��	h ��@�E=!s4@!yԜ�!?�Y�m�@�F`׋ٿ}Dj�w��@)��9�4@�P�͐!?�����@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@�b	��ٿ:y�hl��@7�Lv4@�l�%�!?�t���@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���1�ٿ����@F""�4@(%�6��!?0 �_��@���6�ٿd�w%���@�d}��4@l�H���!?�a~́��@0Ѥ�ŏٿD��\��@tf^��4@[^COb�!?���3��@� �ΊٿR6b
��@��>CT4@��x�N�!?�-s;�@� �ΊٿR6b
��@��>CT4@��x�N�!?�-s;�@� �ΊٿR6b
��@��>CT4@��x�N�!?�-s;�@� �ΊٿR6b
��@��>CT4@��x�N�!?�-s;�@� �ΊٿR6b
��@��>CT4@��x�N�!?�-s;�@[�3���ٿ���d��@ڱw;4@\�AW�!?S�Z���@[�3���ٿ���d��@ڱw;4@\�AW�!?S�Z���@.u}/��ٿHX�r�@#N��S4@k���r�!?�G5�5�@.u}/��ٿHX�r�@#N��S4@k���r�!?�G5�5�@.u}/��ٿHX�r�@#N��S4@k���r�!?�G5�5�@.u}/��ٿHX�r�@#N��S4@k���r�!?�G5�5�@��E΍ٿ	��]��@ ��4@@����!?;�9N��@B;���ٿ��*j�@vC9�^4@���\]�!?�Aͥ*�@B;���ٿ��*j�@vC9�^4@���\]�!?�Aͥ*�@��/@�ٿ��}�֍�@s���f4@X���|�!?�
^�_�@��/@�ٿ��}�֍�@s���f4@X���|�!?�
^�_�@��/@�ٿ��}�֍�@s���f4@X���|�!?�
^�_�@�V�Hj�ٿm�[%4��@����
4@��-�!?�v_J���@�V�Hj�ٿm�[%4��@����
4@��-�!?�v_J���@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@/�r#�ٿ�^כ�@R����4@wb@��!?�Cl��@�8�_Ȍٿ��7w��@|��ه4@��AV��!?���U�@�8�_Ȍٿ��7w��@|��ه4@��AV��!?���U�@��9b��ٿ�lu���@hk!*4@�o��!?o4<�D�@��9b��ٿ�lu���@hk!*4@�o��!?o4<�D�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@>����ٿg�'��G�@jH�/a4@�&e$��!?�\1�sL�@+�5��ٿd�_��@��x��4@���Nڐ!?�1�p��@+�5��ٿd�_��@��x��4@���Nڐ!?�1�p��@+�5��ٿd�_��@��x��4@���Nڐ!?�1�p��@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@��w�ٿ�Q0+��@���~�4@�t�ΐ!?��U�t�@t�7.(�ٿpGKq��@�v_�4@�)�!��!?P�ɒ$P�@t�7.(�ٿpGKq��@�v_�4@�)�!��!?P�ɒ$P�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@�ϼ���ٿ��E�`9�@��L��4@�Ȼ`�!?����s�@��D��ٿM�� J��@`��4@2���!?���5��@��D��ٿM�� J��@`��4@2���!?���5��@��D��ٿM�� J��@`��4@2���!?���5��@<�NDN�ٿZS����@�K;r4@��7��!?���7H��@<�NDN�ٿZS����@�K;r4@��7��!?���7H��@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@$s�N�ٿ��.%��@��E�4@��8�!? ���5�@���HA�ٿ�����@�dE4@qS����!?l��YH��@���HA�ٿ�����@�dE4@qS����!?l��YH��@���HA�ٿ�����@�dE4@qS����!?l��YH��@���HA�ٿ�����@�dE4@qS����!?l��YH��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@�z
��ٿƚŬ�C�@�d9�4@�)o���!?�?#��@?GV�}ٿ$��w��@�3p7�4@�-7��!?�<��9��@OS��{ٿb]6a���@�:բ�4@}Hu�!?��i���@OS��{ٿb]6a���@�:բ�4@}Hu�!?��i���@OS��{ٿb]6a���@�:բ�4@}Hu�!?��i���@2R#Q�ٿ?%	W|��@���$�4@D3�N�!?F�(��4�@2R#Q�ٿ?%	W|��@���$�4@D3�N�!?F�(��4�@2R#Q�ٿ?%	W|��@���$�4@D3�N�!?F�(��4�@1Fr��ٿ��h�sf�@�Mc&4@��^��!?
F�>���@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@jn���ٿ�C�w}�@ε^!E4@GZ�`ʐ!?�,-w�F�@s!Jc��ٿr��n*�@Oڀ[4@G6G�ސ!?Ș�"�@s!Jc��ٿr��n*�@Oڀ[4@G6G�ސ!?Ș�"�@s!Jc��ٿr��n*�@Oڀ[4@G6G�ސ!?Ș�"�@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@kS}3�ٿFNfY׼�@hJ�HU�3@�2��e�!?�f���@�^e��ٿ K~�	�@��O�q4@�x��!?�����@��x�}ٿφ�W�@����{4@A-A>��!?#������@C�	�ٿ�!�4�@���$4@��1�!?<����@C�	�ٿ�!�4�@���$4@��1�!?<����@C�	�ٿ�!�4�@���$4@��1�!?<����@�mnU��ٿ"�Y�Ĭ�@�|ת�4@/%ݫ��!?X��z��@�mnU��ٿ"�Y�Ĭ�@�|ת�4@/%ݫ��!?X��z��@�mnU��ٿ"�Y�Ĭ�@�|ת�4@/%ݫ��!?X��z��@�mnU��ٿ"�Y�Ĭ�@�|ת�4@/%ݫ��!?X��z��@�mnU��ٿ"�Y�Ĭ�@�|ת�4@/%ݫ��!?X��z��@7�Xօٿѝq���@�O 4@�5�ސ!?H~uʒ�@7�Xօٿѝq���@�O 4@�5�ސ!?H~uʒ�@7�Xօٿѝq���@�O 4@�5�ސ!?H~uʒ�@7�Xօٿѝq���@�O 4@�5�ސ!?H~uʒ�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@m�,O�}ٿ��`��@A��(4@-qΐ!?�t�vEH�@��ӖG�ٿ<�`�[.�@chL��4@��*�!?��#9�@��ӖG�ٿ<�`�[.�@chL��4@��*�!?��#9�@��ӖG�ٿ<�`�[.�@chL��4@��*�!?��#9�@��ӖG�ٿ<�`�[.�@chL��4@��*�!?��#9�@��ӖG�ٿ<�`�[.�@chL��4@��*�!?��#9�@��7�ٿS�3*��@�Ci�4@�b��4�!?�/��#C�@�W�-�ٿ0���Y�@�;O�4@ܓ���!?�� ؔ�@5U�n�{ٿhA���@7�CZ4@�����!?�xf;Q��@5U�n�{ٿhA���@7�CZ4@�����!?�xf;Q��@�>vw�ٿ���@D�㝸4@��-	�!?򻽵@5�@����ٿ%���v�@q{>rV4@+�hI�!?3,芆�@����ٿ%���v�@q{>rV4@+�hI�!?3,芆�@����ٿ%���v�@q{>rV4@+�hI�!?3,芆�@�)�a��ٿ�*�9�t�@^��wf4@~�^�!?v9"��
�@V�e�	�ٿW��r)�@�g"�4@g�聐!?���rщ�@9O���ٿ $�B�@/�y>4@j��7�!?����,G�@9O���ٿ $�B�@/�y>4@j��7�!?����,G�@9O���ٿ $�B�@/�y>4@j��7�!?����,G�@>A\��ٿ
��$���@b�N�m4@��Bm��!?���q��@��{�ٿ7fG���@���9.4@�����!?�ԓ�]��@��{�ٿ7fG���@���9.4@�����!?�ԓ�]��@��{�ٿ7fG���@���9.4@�����!?�ԓ�]��@3�z�F�ٿ.X���'�@KQ�O4@u�9��!?�64J=��@3�z�F�ٿ.X���'�@KQ�O4@u�9��!?�64J=��@3�z�F�ٿ.X���'�@KQ�O4@u�9��!?�64J=��@3�z�F�ٿ.X���'�@KQ�O4@u�9��!?�64J=��@x<�n�ٿf���~s�@e[n4@ry땐!?�e{���@x<�n�ٿf���~s�@e[n4@ry땐!?�e{���@x<�n�ٿf���~s�@e[n4@ry땐!?�e{���@�弽�ٿԑ��0��@�#� <4@�0̲�!?��hA�`�@�弽�ٿԑ��0��@�#� <4@�0̲�!?��hA�`�@�弽�ٿԑ��0��@�#� <4@�0̲�!?��hA�`�@�弽�ٿԑ��0��@�#� <4@�0̲�!?��hA�`�@�ar��ٿIlTF���@ Oy �4@������!?|0����@�ar��ٿIlTF���@ Oy �4@������!?|0����@�ar��ٿIlTF���@ Oy �4@������!?|0����@��B�ٿd���.�@�Y�y4@�T	鵐!?�#��@��@��B�ٿd���.�@�Y�y4@�T	鵐!?�#��@��@��B�ٿd���.�@�Y�y4@�T	鵐!?�#��@��@����4�ٿK�V�?\�@
R��#4@��Y(ݐ!?o	'�Y	�@U���ωٿB�#���@h�Ad�4@0�e_א!?d_Q�׹�@U���ωٿB�#���@h�Ad�4@0�e_א!?d_Q�׹�@U���ωٿB�#���@h�Ad�4@0�e_א!?d_Q�׹�@U���ωٿB�#���@h�Ad�4@0�e_א!?d_Q�׹�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@Y���b�ٿ�	����@Q6� �4@�4�Ő!?ڹ ZH%�@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�J*��ٿ�yy���@�����4@��y�͐!?��n!���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�ՙc�ٿ��"��B�@G�o)4@�қ�ؐ!?�u�q���@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@�g���ٿ!����@��H�X4@�g{�Ő!?lEk#G�@`�A�ٿ��c��@��4@���K��!?�8Y���@`�A�ٿ��c��@��4@���K��!?�8Y���@����zٿ�)b���@R��4@��eB �!?��׵�@�@����zٿ�)b���@R��4@��eB �!?��׵�@�@����zٿ�)b���@R��4@��eB �!?��׵�@�@����zٿ�)b���@R��4@��eB �!?��׵�@�@/h\_�ٿ	|��l�@͒�x�4@�����!?���F�F�@/h\_�ٿ	|��l�@͒�x�4@�����!?���F�F�@/h\_�ٿ	|��l�@͒�x�4@�����!?���F�F�@/h\_�ٿ	|��l�@͒�x�4@�����!?���F�F�@Nɚ���ٿ���V�l�@^_�VM4@��,Đ!?Z�����@Nɚ���ٿ���V�l�@^_�VM4@��,Đ!?Z�����@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@�;׆�ٿQ'��1��@����4@��W��!?��n��E�@��&��ٿ颐����@�����4@��'��!?L�c���@��&��ٿ颐����@�����4@��'��!?L�c���@l���ٿIf�B��@�7s ��3@r��ZА!?hÿ"g�@l���ٿIf�B��@�7s ��3@r��ZА!?hÿ"g�@l���ٿIf�B��@�7s ��3@r��ZА!?hÿ"g�@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@������ٿJ꿱���@P;�~�4@��{ћ�!?��7��@��Q��ٿ/�����@ƕ�r4@I&���!?�G=`F��@��Q��ٿ/�����@ƕ�r4@I&���!?�G=`F��@��Q��ٿ/�����@ƕ�r4@I&���!?�G=`F��@�s#\"�ٿ���f��@e���4@���ΐ!?R����j�@�s#\"�ٿ���f��@e���4@���ΐ!?R����j�@�s#\"�ٿ���f��@e���4@���ΐ!?R����j�@�s#\"�ٿ���f��@e���4@���ΐ!?R����j�@�s#\"�ٿ���f��@e���4@���ΐ!?R����j�@��ԉٿ��|���@����4@a![��!?�0�m#�@��ԉٿ��|���@����4@a![��!?�0�m#�@��kgŋٿ�<�ii[�@�Y�74@	�{�!?W^d��`�@��l��ٿ��Jr>)�@7��j�4@�e����!?���V���@��l��ٿ��Jr>)�@7��j�4@�e����!?���V���@��U{�ٿ(-|k�4�@:X�}Z4@2�@��!?PBy����@b�7pl�ٿ��R����@��Js4@���@��!?(͖�aA�@b�7pl�ٿ��R����@��Js4@���@��!?(͖�aA�@QƠ2}�ٿS�Mf���@{3p�|4@�[�K��!?���w��@QƠ2}�ٿS�Mf���@{3p�|4@�[�K��!?���w��@QƠ2}�ٿS�Mf���@{3p�|4@�[�K��!?���w��@QƠ2}�ٿS�Mf���@{3p�|4@�[�K��!?���w��@QƠ2}�ٿS�Mf���@{3p�|4@�[�K��!?���w��@��8��ٿ�b/}���@��=4@�ݿ�!?#����@��8��ٿ�b/}���@��=4@�ݿ�!?#����@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@~�R
ٿ텘O��@�R���4@�n���!?�c�ѠN�@�;���ٿ���� �@�8�uG4@�-~��!?p�,_|�@�;���ٿ���� �@�8�uG4@�-~��!?p�,_|�@�;���ٿ���� �@�8�uG4@�-~��!?p�,_|�@�;���ٿ���� �@�8�uG4@�-~��!?p�,_|�@d5s��ٿ�e�ذ[�@9�
6 4@���(��!?R^.�\�@d5s��ٿ�e�ذ[�@9�
6 4@���(��!?R^.�\�@d5s��ٿ�e�ذ[�@9�
6 4@���(��!?R^.�\�@d5s��ٿ�e�ذ[�@9�
6 4@���(��!?R^.�\�@ �3�ٿh�	��7�@;�}3� 4@�o���!?���&��@ �3�ٿh�	��7�@;�}3� 4@�o���!?���&��@ �3�ٿh�	��7�@;�}3� 4@�o���!?���&��@ �3�ٿh�	��7�@;�}3� 4@�o���!?���&��@ �3�ٿh�	��7�@;�}3� 4@�o���!?���&��@k�1��ٿ@F��-}�@O��4@����!?b��,i��@k�1��ٿ@F��-}�@O��4@����!?b��,i��@k�1��ٿ@F��-}�@O��4@����!?b��,i��@k�1��ٿ@F��-}�@O��4@����!?b��,i��@�t-�$�ٿ痁���@�����4@qtު�!?\�X{�x�@�t-�$�ٿ痁���@�����4@qtު�!?\�X{�x�@P��Ìٿ2�M���@H���4@�&v�P�!?�%�*�]�@�q���ٿU�]Q��@W���4@7����!?�_��U��@�q���ٿU�]Q��@W���4@7����!?�_��U��@�q���ٿU�]Q��@W���4@7����!?�_��U��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@7�W���ٿ�#�UQq�@�yiMf4@]�鱐!?��$r��@X2eކٿ ��8��@}�gH4@�z�֐!?ٌ���@X2eކٿ ��8��@}�gH4@�z�֐!?ٌ���@X2eކٿ ��8��@}�gH4@�z�֐!?ٌ���@X2eކٿ ��8��@}�gH4@�z�֐!?ٌ���@�"FV�ٿ��ըQ0�@ o�R4@��!�Ӑ!?�lqZY�@�"FV�ٿ��ըQ0�@ o�R4@��!�Ӑ!?�lqZY�@���Fl�ٿ�\ -�)�@M�@�4@���	��!?�������@���Fl�ٿ�\ -�)�@M�@�4@���	��!?�������@���Fl�ٿ�\ -�)�@M�@�4@���	��!?�������@���Fl�ٿ�\ -�)�@M�@�4@���	��!?�������@���Fl�ٿ�\ -�)�@M�@�4@���	��!?�������@���酆ٿ:ݣ�=��@73��4@F�vĐ!?0?p_S�@���酆ٿ:ݣ�=��@73��4@F�vĐ!?0?p_S�@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@]pB� �ٿc+C]'�@e���K4@�/j�̐!?#�����@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@�?�C�ٿ� N4��@�o �$4@'OCʐ!?ˌv�w@�@`�Y�ٿ5�t7���@#E�44@QZ��!?:�~Le��@`�Y�ٿ5�t7���@#E�44@QZ��!?:�~Le��@`�Y�ٿ5�t7���@#E�44@QZ��!?:�~Le��@��&aA�ٿ�z�|���@F�Ot4@a|��%�!??���@��&aA�ٿ�z�|���@F�Ot4@a|��%�!??���@��&aA�ٿ�z�|���@F�Ot4@a|��%�!??���@��&aA�ٿ�z�|���@F�Ot4@a|��%�!??���@tG���ٿ�m�Q���@��ؼ�4@J�Y��!?�j=�w�@tG���ٿ�m�Q���@��ؼ�4@J�Y��!?�j=�w�@tG���ٿ�m�Q���@��ؼ�4@J�Y��!?�j=�w�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@[���ٿ3��+�@��l 4@�l��!?L�rX�@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@�y��ٿ-���.�@iD���4@w��N�!?m�m��@q:�T�ٿ��
��@���ji4@h����!?2ŀ.�m�@q:�T�ٿ��
��@���ji4@h����!?2ŀ.�m�@q:�T�ٿ��
��@���ji4@h����!?2ŀ.�m�@z��Q�ٿMvMR��@f�Ͳ4@~���А!?7�xn�_�@z��Q�ٿMvMR��@f�Ͳ4@~���А!?7�xn�_�@z��Q�ٿMvMR��@f�Ͳ4@~���А!?7�xn�_�@�}-��ٿ�	���@���p4@�gz��!?Y�[�@�@�}-��ٿ�	���@���p4@�gz��!?Y�[�@�@�}-��ٿ�	���@���p4@�gz��!?Y�[�@�@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@Y�=�ӆٿ�@��{��@���d 4@�sH�.�!?�"�=��@H\ʨZ�ٿ�Z����@:��4@E�u�ڐ!?������@�┖o�ٿ�>��H9�@��
>4@�����!?��.�A��@�┖o�ٿ�>��H9�@��
>4@�����!?��.�A��@�┖o�ٿ�>��H9�@��
>4@�����!?��.�A��@�┖o�ٿ�>��H9�@��
>4@�����!?��.�A��@%�h���ٿیb���@_�y�� 4@E�ٮ�!?�O� �@%�h���ٿیb���@_�y�� 4@E�ٮ�!?�O� �@%�h���ٿیb���@_�y�� 4@E�ٮ�!?�O� �@%�h���ٿیb���@_�y�� 4@E�ٮ�!?�O� �@%�h���ٿیb���@_�y�� 4@E�ٮ�!?�O� �@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@Y)k�ٿW}��a��@���/j4@���T�!?�%����@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@,�-�g�ٿ3��?"�@��#��4@�u�Td�!?$��+���@G��f��ٿۋKc_N�@�=0}4@����!?�(�1��@G��f��ٿۋKc_N�@�=0}4@����!?�(�1��@G��f��ٿۋKc_N�@�=0}4@����!?�(�1��@��-g�ٿw���,�@�)m�{4@��Ԑ!?���4eN�@��-g�ٿw���,�@�)m�{4@��Ԑ!?���4eN�@���n�ٿ 6���@3J�/4@^��7�!?�a��/�@���n�ٿ 6���@3J�/4@^��7�!?�a��/�@���n�ٿ 6���@3J�/4@^��7�!?�a��/�@�4m�ٿ7�B����@ :�4@�8='�!?�'w��@܃0���ٿ ڙnG��@0��%I4@����!?�i
(�v�@܃0���ٿ ڙnG��@0��%I4@����!?�i
(�v�@܃0���ٿ ڙnG��@0��%I4@����!?�i
(�v�@܃0���ٿ ڙnG��@0��%I4@����!?�i
(�v�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@��3�L�ٿ�$�K	�@}����3@��\��!?|Y��g�@g��!��ٿ�&��@m��/4@$�Ә��!?���Z�@g��!��ٿ�&��@m��/4@$�Ә��!?���Z�@g��!��ٿ�&��@m��/4@$�Ә��!?���Z�@!7�ٿ���s/�@��L�4@l
9���!?���H��@!7�ٿ���s/�@��L�4@l
9���!?���H��@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�K]���ٿjh`�x=�@m��z4@���%��!?Ƿ%�.�@�1Ap��ٿ��Yٞ$�@�>k 4@W�lNĐ!?�B����@�}�ٿ�a(/���@k��*4@h!0%j�!?6j�W�y�@�}�ٿ�a(/���@k��*4@h!0%j�!?6j�W�y�@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@4�o��ٿ���g�@�R�&d4@��H3��!?�_˄��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@��%b�ٿ�^�E���@K��74@_�%��!?U�.-m��@5D�W�ٿ޳��ߝ�@�Fx��4@4��ː!?�BS+��@5D�W�ٿ޳��ߝ�@�Fx��4@4��ː!?�BS+��@5D�W�ٿ޳��ߝ�@�Fx��4@4��ː!?�BS+��@5D�W�ٿ޳��ߝ�@�Fx��4@4��ː!?�BS+��@5D�W�ٿ޳��ߝ�@�Fx��4@4��ː!?�BS+��@U���&|ٿ�W����@�c��4@�痡Ӑ!?�4�oq�@�_�;{ٿ��~���@�1�ޛ4@��i��!?����US�@�_�;{ٿ��~���@�1�ޛ4@��i��!?����US�@�_�;{ٿ��~���@�1�ޛ4@��i��!?����US�@�_�;{ٿ��~���@�1�ޛ4@��i��!?����US�@���b�ٿ'r�����@�]�:!4@���
��!?c���uf�@j�t �ٿur(k���@�)D��4@��	�!?�j��V��@j�t �ٿur(k���@�)D��4@��	�!?�j��V��@j�t �ٿur(k���@�)D��4@��	�!?�j��V��@j�t �ٿur(k���@�)D��4@��	�!?�j��V��@v�@>a�ٿ��'E���@b�J�K4@���Ő!?Ճj�j��@v�@>a�ٿ��'E���@b�J�K4@���Ő!?Ճj�j��@v�@>a�ٿ��'E���@b�J�K4@���Ő!?Ճj�j��@v�@>a�ٿ��'E���@b�J�K4@���Ő!?Ճj�j��@v�@>a�ٿ��'E���@b�J�K4@���Ő!?Ճj�j��@���6�ٿ;]T��7�@(�B�4@x��ߐ!?͝���i�@C_���ٿ�~����@�Mǘ|	4@Z�C�!?0��=m8�@C_���ٿ�~����@�Mǘ|	4@Z�C�!?0��=m8�@C_���ٿ�~����@�Mǘ|	4@Z�C�!?0��=m8�@�J�~ٿ������@gc6�4@��a���!?X�Es��@����1�ٿ��\S*��@�G���4@���J�!?̶dA0p�@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@��Uz��ٿ}�E���@+�sx�4@{ ux�!?g8K�b��@#�����ٿ	H�Lt%�@_mn4@;�
җ�!?'�Ӡ�@#�����ٿ	H�Lt%�@_mn4@;�
җ�!?'�Ӡ�@��2�4�ٿ�bc�f�@�$ĝ4@D	mb��!?Uf�J	��@ޑ][��ٿRG鮠�@O0GL�4@h����!?ܖ�)��@ޑ][��ٿRG鮠�@O0GL�4@h����!?ܖ�)��@ޑ][��ٿRG鮠�@O0GL�4@h����!?ܖ�)��@r�:~ٿ,���Nq�@8wC�4@�Wq]�!?�s�E���@r�:~ٿ,���Nq�@8wC�4@�Wq]�!?�s�E���@r�:~ٿ,���Nq�@8wC�4@�Wq]�!?�s�E���@F�2N�ٿ(y���@Q�ϴ4@���!?.���G��@F�2N�ٿ(y���@Q�ϴ4@���!?.���G��@F�2N�ٿ(y���@Q�ϴ4@���!?.���G��@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@&B����ٿ!G0��@��YY� 4@�h拻�!?��M����@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��Qトٿk�I�#��@E\,;4@)�
��!?�!� �^�@��\E�ٿ�Tm]�@֐�4@n����!?C;�t�@��\E�ٿ�Tm]�@֐�4@n����!?C;�t�@��\E�ٿ�Tm]�@֐�4@n����!?C;�t�@��\E�ٿ�Tm]�@֐�4@n����!?C;�t�@��\E�ٿ�Tm]�@֐�4@n����!?C;�t�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@��M�ٿ���&��@Z�pj�4@܏�VĐ!?ƿ�΄x�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@7�s.ٿ&,e���@;���4@+� ���!?)�1�?L�@��R�ٿ�>����@��8�'4@cF����!?�xt$��@��R�ٿ�>����@��8�'4@cF����!?�xt$��@��R�ٿ�>����@��8�'4@cF����!?�xt$��@>�g��ٿY�����@�X�(4@�\G��!?>�U���@>�g��ٿY�����@�X�(4@�\G��!?>�U���@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@�.�孃ٿ�g��+��@��P�4@Q��!?�9�'m�@r	u�<�ٿ��0Z��@��Ja4@Ȗ�֐!?@�HsmT�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�oK��ٿ�F0�L��@ڂOC�4@
�Ȑ!?R6�K�u�@�����ٿ4����@�S>׼4@9�!?���jZ�@�����ٿ4����@�S>׼4@9�!?���jZ�@�ASԈٿC�a"�^�@��d��4@��B���!?����]&�@�ASԈٿC�a"�^�@��d��4@��B���!?����]&�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@d��{��ٿb�I���@�-y�4@��(���!?>����k�@�Z]�w�ٿ!9�h��@���h4@u�j�!?
z��@R���ٿԌj���@Z~��v 4@�M��Ȑ!?/o���b�@R���ٿԌj���@Z~��v 4@�M��Ȑ!?/o���b�@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@���ٿ�/���@Yҍ"k4@�n@',�!?�o����@�3TE�ٿ:���X��@�k9jM4@@�򯡐!?ğ~���@�3TE�ٿ:���X��@�k9jM4@@�򯡐!?ğ~���@���?�ٿ˩c-��@�ި�4@�~��Ɛ!?1J���v�@���?�ٿ˩c-��@�ި�4@�~��Ɛ!?1J���v�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@���%�ٿ`�\��@ш�x4@͡�Ő!?��/�v(�@uҚ�ˇٿ�=C�>�@��Jk%4@�*k��!?[piA��@���t��ٿa��y^�@�κj�4@�w�/�!?�_�9Ld�@���t��ٿa��y^�@�κj�4@�w�/�!?�_�9Ld�@Lg���ٿ�F��!�@�2Z6�4@���V�!?�`P���@:��Ȕ�ٿ��o��@��f4@c�Ae.�!?&��Pg��@:��Ȕ�ٿ��o��@��f4@c�Ae.�!?&��Pg��@0V��{�ٿۃ/S�*�@��[4@�-�!?�1����@0\�O|ٿ�I��@�"a|�4@�����!?V�B-��@0\�O|ٿ�I��@�"a|�4@�����!?V�B-��@�>Ҳ��ٿP��	.��@/Ï��4@��t��!?v�֊�G�@��w6�ٿȠ')�u�@�\+LA4@�t��!?,�{��@B�
�ׁٿ"��f��@6
�dS4@�{s��!?/m��,�@u�a��ٿ�k�٥��@���VA4@F��Ȑ!?{��B�x�@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@p��5�ٿ�8�w��@[��xE4@�O��!?Z�ץ���@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@��7�ٿ�4J�9��@n�L4@+��/w�!?��瘰K�@B���J�ٿ| :Ի�@<�h��4@�eY�v�!?��Mx�\�@B���J�ٿ| :Ի�@<�h��4@�eY�v�!?��Mx�\�@��pA4�ٿz�t��@�0��}4@�!F��!?�~f[�@�����ٿ��瑑��@�>s�64@ ��L��!?P���?�@��S|ٿ��B�T��@��Y��4@����!?C����@ T+�s}ٿA��z�|�@�X"R4@x���!?A���8�@ T+�s}ٿA��z�|�@�X"R4@x���!?A���8�@ T+�s}ٿA��z�|�@�X"R4@x���!?A���8�@ T+�s}ٿA��z�|�@�X"R4@x���!?A���8�@ T+�s}ٿA��z�|�@�X"R4@x���!?A���8�@�	�]$|ٿ�\S��@���?4@;8���!?D�=�˅�@ٟ%A-�ٿ�+*����@Zqs64@FR�֓�!?�u�U�@ٟ%A-�ٿ�+*����@Zqs64@FR�֓�!?�u�U�@ٟ%A-�ٿ�+*����@Zqs64@FR�֓�!?�u�U�@ٟ%A-�ٿ�+*����@Zqs64@FR�֓�!?�u�U�@�t�_��ٿ��̺;%�@*��n�4@�U;���!?��W��}�@�t�_��ٿ��̺;%�@*��n�4@�U;���!?��W��}�@�t�_��ٿ��̺;%�@*��n�4@�U;���!?��W��}�@�t�_��ٿ��̺;%�@*��n�4@�U;���!?��W��}�@Y����ٿt�6ʂ�@_³ԙ4@ۀAz�!?>rb��R�@�����ٿexVٌ�@�I�;4@W��!?�
	��@;�=�r�ٿJ��ߠ��@�M �24@����!?~��.N�@̟��ٿ*k�J�n�@Q9B�!4@u��-��!?�Rn�G�@̟��ٿ*k�J�n�@Q9B�!4@u��-��!?�Rn�G�@̟��ٿ*k�J�n�@Q9B�!4@u��-��!?�Rn�G�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@Qw��ٿ�@�6K��@�p(�4@��ʹ�!?�?�S	�@�dCi��ٿW���·�@ �X
4@Eg� ��!?�S��*��@�dCi��ٿW���·�@ �X
4@Eg� ��!?�S��*��@�dCi��ٿW���·�@ �X
4@Eg� ��!?�S��*��@�dCi��ٿW���·�@ �X
4@Eg� ��!?�S��*��@�'���ٿ�]���@�G���4@�q0�s�!?҄߸`�@�'���ٿ�]���@�G���4@�q0�s�!?҄߸`�@�'���ٿ�]���@�G���4@�q0�s�!?҄߸`�@.�Z��ٿz6W��U�@��Q�4@�pAۭ�!?�0��@.�Z��ٿz6W��U�@��Q�4@�pAۭ�!?�0��@_�R7z�ٿ��z�-�@p���y4@�|	�А!?C���Gl�@_�R7z�ٿ��z�-�@p���y4@�|	�А!?C���Gl�@_�R7z�ٿ��z�-�@p���y4@�|	�А!?C���Gl�@_�R7z�ٿ��z�-�@p���y4@�|	�А!?C���Gl�@_�R7z�ٿ��z�-�@p���y4@�|	�А!?C���Gl�@a��އٿ4��w�@��h��4@�F�ઐ!?�hv)�(�@a��އٿ4��w�@��h��4@�F�ઐ!?�hv)�(�@ޢ��Y�ٿ�B�2�
�@8gtE4@��Z���!??m���@ޢ��Y�ٿ�B�2�
�@8gtE4@��Z���!??m���@ޢ��Y�ٿ�B�2�
�@8gtE4@��Z���!??m���@n1�I݁ٿϊ���@��
14@�ʙ�!?������@n1�I݁ٿϊ���@��
14@�ʙ�!?������@n1�I݁ٿϊ���@��
14@�ʙ�!?������@n1�I݁ٿϊ���@��
14@�ʙ�!?������@n1�I݁ٿϊ���@��
14@�ʙ�!?������@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@#7H��ٿ�v)���@_� �e4@M���!?|j��b�@���O��ٿ]Ye�a�@pot��4@.;T���!?V-�S��@�K�&~�ٿ#�i��@j�mk�4@��H��!?h����@^�V�r�ٿ�߀l���@���)4@�t.[�!?��-"���@^�V�r�ٿ�߀l���@���)4@�t.[�!?��-"���@9��%�ٿ�ކ����@�g4@`����!?��P��@9��%�ٿ�ކ����@�g4@`����!?��P��@9��%�ٿ�ކ����@�g4@`����!?��P��@�bP�ٿ��rܸ�@����4@���n�!?��Ri.�@�� oٿ�6ny&�@��&�V4@��"���!?��WU]�@��lt/�ٿ\��;��@�R��4@v����!?�c����@��lt/�ٿ\��;��@�R��4@v����!?�c����@��lt/�ٿ\��;��@�R��4@v����!?�c����@��lt/�ٿ\��;��@�R��4@v����!?�c����@��lt/�ٿ\��;��@�R��4@v����!?�c����@�w�Pxٿ�"D)C�@�ɸ�4@��^��!?�v��v�@�p��zٿ����!��@��{\4@T�e���!?Ec��A�@ݚ\�ٿ�������@ g�7v
4@;�Ϭ�!?�&���@ݚ\�ٿ�������@ g�7v
4@;�Ϭ�!?�&���@���Mٿ��L	l6�@j�Ǳ
4@�8=��!?���E��@���Mٿ��L	l6�@j�Ǳ
4@�8=��!?���E��@ k��xٿ��&�Z�@1y[\4@}�z��!?�7��`��@g�yaxٿ�pI��>�@0I�{�	4@�%���!?����O��@g�yaxٿ�pI��>�@0I�{�	4@�%���!?����O��@g�yaxٿ�pI��>�@0I�{�	4@�%���!?����O��@z�vʻuٿn�4�Z^�@}�T�4@�M���!?ί�I�6�@z�vʻuٿn�4�Z^�@}�T�4@�M���!?ί�I�6�@z�vʻuٿn�4�Z^�@}�T�4@�M���!?ί�I�6�@z�vʻuٿn�4�Z^�@}�T�4@�M���!?ί�I�6�@�˨�yٿ�y8���@�xR74@�^Y�!?�G����@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@-�V�ٿ`�v��@�;P�4@O�Wm�!?�2T���@�E�q�ٿN7$��@��hN[4@Ӟ� �!?W�nr���@�E�q�ٿN7$��@��hN[4@Ӟ� �!?W�nr���@�E�q�ٿN7$��@��hN[4@Ӟ� �!?W�nr���@�E�q�ٿN7$��@��hN[4@Ӟ� �!?W�nr���@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@�3zqB�ٿĻ�I��@����4@�H� �!?�V�c�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@u7�8,�ٿ/�pn��@��~�4@p���!?C�
��k�@�5���ٿ؝�����@��h�Y 4@��ڳ��!?K���~��@�5���ٿ؝�����@��h�Y 4@��ڳ��!?K���~��@�5���ٿ؝�����@��h�Y 4@��ڳ��!?K���~��@�5���ٿ؝�����@��h�Y 4@��ڳ��!?K���~��@�5���ٿ؝�����@��h�Y 4@��ڳ��!?K���~��@��)f�ٿ+�M�02�@��o��3@�}3���!?s&��@��)f�ٿ+�M�02�@��o��3@�}3���!?s&��@��)f�ٿ+�M�02�@��o��3@�}3���!?s&��@��)f�ٿ+�M�02�@��o��3@�}3���!?s&��@��Vٿ7��:t�@��ӭ�4@]�1+�!?� yP��@��Vٿ7��:t�@��ӭ�4@]�1+�!?� yP��@�*�˃ٿ�x�\1&�@fI� 4@V�tX�!?��4�@�\&&މٿ�/(�@F��H� 4@��ŝ�!?���Ι��@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@�Zp�}�ٿ:Y���N�@�eY� 4@hF#�!?��mL�@)�$�ٿ'Y ����@@o��4@���ڐ!?o^��@)�$�ٿ'Y ����@@o��4@���ڐ!?o^��@)�$�ٿ'Y ����@@o��4@���ڐ!?o^��@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@^=źt�ٿ���	1-�@i�>�4@\��
�!?�Rk�%{�@�=a��ٿLS1��@��@<�4@�I��ǐ!?hQ=F��@�=a��ٿLS1��@��@<�4@�I��ǐ!?hQ=F��@!
��S�ٿd����@��@oV4@��=h��!?m�g ��@!
��S�ٿd����@��@oV4@��=h��!?m�g ��@!
��S�ٿd����@��@oV4@��=h��!?m�g ��@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@f�����ٿ���\�@����4@�����!?��(�@N�QF�ٿ��]`n�@z�4@�4@�����!?�� =��@N�QF�ٿ��]`n�@z�4@�4@�����!?�� =��@N�QF�ٿ��]`n�@z�4@�4@�����!?�� =��@N�QF�ٿ��]`n�@z�4@�4@�����!?�� =��@N�QF�ٿ��]`n�@z�4@�4@�����!?�� =��@�a�ٿ�њ��@���k�4@́Z���!?p�C�/�@���>�ٿc�q,�w�@yF�I4@�5���!?�eC�Gs�@���>�ٿc�q,�w�@yF�I4@�5���!?�eC�Gs�@���>�ٿc�q,�w�@yF�I4@�5���!?�eC�Gs�@�_i`Q�ٿ��7���@��kd4@�m���!?t����;�@��\u��ٿ3R�֤�@DK(� 4@��ِ!?*ȡ�I�@��\u��ٿ3R�֤�@DK(� 4@��ِ!?*ȡ�I�@�uK!�ٿ��aE9�@�A`� 4@K_!�!?Wq�����@�uK!�ٿ��aE9�@�A`� 4@K_!�!?Wq�����@�uK!�ٿ��aE9�@�A`� 4@K_!�!?Wq�����@(��_�ٿ�f�#���@JSt� 4@��h��!?����@(��_�ٿ�f�#���@JSt� 4@��h��!?����@(��_�ٿ�f�#���@JSt� 4@��h��!?����@(��_�ٿ�f�#���@JSt� 4@��h��!?����@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@�y�,ٿKzD|���@N$�?4@��L�ߐ!?�;
sG�@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@����ٿ�ēm��@��x4@�ʺ5��!?�+� ��@QE6���ٿ�+���@���(�4@D7 �!?�-5����@QE6���ٿ�+���@���(�4@D7 �!?�-5����@W����ٿ���(��@�丑84@��M�!?����?��@W����ٿ���(��@�丑84@��M�!?����?��@W����ٿ���(��@�丑84@��M�!?����?��@W����ٿ���(��@�丑84@��M�!?����?��@���s�ٿմ����@� j�?4@kZM� �!?`y 73e�@���s�ٿմ����@� j�?4@kZM� �!?`y 73e�@���s�ٿմ����@� j�?4@kZM� �!?`y 73e�@���s�ٿմ����@� j�?4@kZM� �!?`y 73e�@���s�ٿմ����@� j�?4@kZM� �!?`y 73e�@��s�ٿ�P��=��@�:�+4@���_ɐ!?�G�&&]�@��s�ٿ�P��=��@�:�+4@���_ɐ!?�G�&&]�@��s�ٿ�P��=��@�:�+4@���_ɐ!?�G�&&]�@U�vrY�ٿε�t��@��ϗe4@y�ɷ+�!?,��7�d�@x�4�y�ٿ�����@B��lQ 4@����!?� ��@x�4�y�ٿ�����@B��lQ 4@����!?� ��@x�4�y�ٿ�����@B��lQ 4@����!?� ��@x�4�y�ٿ�����@B��lQ 4@����!?� ��@x�4�y�ٿ�����@B��lQ 4@����!?� ��@x�4�y�ٿ�����@B��lQ 4@����!?� ��@���Z��ٿ��	%~!�@��p�,4@� $��!?���d��@���Z��ٿ��	%~!�@��p�,4@� $��!?���d��@���Z��ٿ��	%~!�@��p�,4@� $��!?���d��@���Z��ٿ��	%~!�@��p�,4@� $��!?���d��@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@	V(=v�ٿυR��@��034@�ϵ*W�!?9ʙT�U�@p:I�ٿo�$��b�@��$1� 4@)�
��!?^g34��@p:I�ٿo�$��b�@��$1� 4@)�
��!?^g34��@k��ٿ���l�;�@\ѽ�r4@�y�6��!?��ZL|H�@k��ٿ���l�;�@\ѽ�r4@�y�6��!?��ZL|H�@�>�⸂ٿ�V_�@�g_�4@,��Ɛ!?�w혤�@�>�⸂ٿ�V_�@�g_�4@,��Ɛ!?�w혤�@�Z�~ٿ� ���@�S8�4@���Ő!?�I��i�@�Z�~ٿ� ���@�S8�4@���Ő!?�I��i�@�Z�~ٿ� ���@�S8�4@���Ő!?�I��i�@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@�8GЇٿ��V��@] �N�4@��ٜ�!?��ˉ��@$�ty��ٿ�B9�1�@��A~4@Tp����!?��c*��@$�ty��ٿ�B9�1�@��A~4@Tp����!?��c*��@$�ty��ٿ�B9�1�@��A~4@Tp����!?��c*��@$�ty��ٿ�B9�1�@��A~4@Tp����!?��c*��@�b��L�ٿ!���>�@M�Z�4@�~0虐!?���y�U�@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@\�٨i�ٿ�g�3�@l�=y4@���b�!?<(l$X��@*ے�1�ٿ�8�֝�@���e�4@��ʈ�!?��\B��@*ے�1�ٿ�8�֝�@���e�4@��ʈ�!?��\B��@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@V�X"܊ٿ��Q`��@*\�mO4@���|��!?D_�\�W�@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@�?�%p�ٿa��אy�@�<�{( 4@̽I�א!?k�o4'��@zŜ,X�ٿ�,I ��@}���'4@4�|�7�!?���l٠�@zŜ,X�ٿ�,I ��@}���'4@4�|�7�!?���l٠�@?�+�{�ٿ�	I�@�O00�4@�L�Zh�!?��I��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@%R�!j�ٿ\/���@�Th�.4@������!?"�\��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@j8u�ٿt[�E�+�@� �4@@8m^�!?P���l��@�2'e�ٿ�C``�?�@��I44@�����!?ڽ��s%�@�2'e�ٿ�C``�?�@��I44@�����!?ڽ��s%�@�$�>�ٿה�
O�@C"럈4@���_Ր!?��X�`�@�D>|@�ٿ�vO[��@��O�4@�抐!?�n�av��@�1G8��ٿ�Bh���@̹SJ@4@�]�z��!?{&�$j�@�1G8��ٿ�Bh���@̹SJ@4@�]�z��!?{&�$j�@�1G8��ٿ�Bh���@̹SJ@4@�]�z��!?{&�$j�@�1G8��ٿ�Bh���@̹SJ@4@�]�z��!?{&�$j�@F�Y�ٿ��!G��@���`4@���|ѐ!?8��v�|�@F�Y�ٿ��!G��@���`4@���|ѐ!?8��v�|�@F�Y�ٿ��!G��@���`4@���|ѐ!?8��v�|�@�e�c�ٿ������@�u�P 4@�KS�!?�p	�P�@�e�c�ٿ������@�u�P 4@�KS�!?�p	�P�@�e�c�ٿ������@�u�P 4@�KS�!?�p	�P�@;*z�3zٿ�׻��@��xle4@~����!?	$e�cv�@;*z�3zٿ�׻��@��xle4@~����!?	$e�cv�@;*z�3zٿ�׻��@��xle4@~����!?	$e�cv�@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@�\'łٿaX��{��@����4@�j<��!?��e��@��:��ٿ�=���<�@<��H4@�x1��!?Dv�e$�@��:��ٿ�=���<�@<��H4@�x1��!?Dv�e$�@��:��ٿ�=���<�@<��H4@�x1��!?Dv�e$�@��:��ٿ�=���<�@<��H4@�x1��!?Dv�e$�@��:��ٿ�=���<�@<��H4@�x1��!?Dv�e$�@�CX3�ٿ`�D ��@7Y�4@�KW�!?I��{���@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@jj�[��ٿŘ���y�@ҽ2�4@2E�`��!?��CA��@�E3Ҹ�ٿ�fh���@X��4@�JYrА!?��e�@�E3Ҹ�ٿ�fh���@X��4@�JYrА!?��e�@^��_�ٿ���G��@�\+m3	4@X����!?l1��@^��_�ٿ���G��@�\+m3	4@X����!?l1��@^��_�ٿ���G��@�\+m3	4@X����!?l1��@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@��ٿ�I��@�@��0�4@�l���!?�7�C�@p��bZ�ٿf �@
!34@F��1��!?��!w�+�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@�`f�m�ٿ�M�Q/�@M`4@���x�!?d�Q�w�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@`x�޲�ٿؗLN��@��A�4@!�
�!?\����_�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@��`�ـٿx�<���@��TNL4@�L��͐!?��ܿ�3�@�/��0�ٿp]j݇��@]<:�4@|���ِ!?��߈��@�/��0�ٿp]j݇��@]<:�4@|���ِ!?��߈��@؉�;Ѓٿ���l��@�.��4@���֐!?��n`��@؉�;Ѓٿ���l��@�.��4@���֐!?��n`��@؉�;Ѓٿ���l��@�.��4@���֐!?��n`��@؉�;Ѓٿ���l��@�.��4@���֐!?��n`��@�/�c�ٿN��]-��@� VsE4@8�3���!?�R���@�/�c�ٿN��]-��@� VsE4@8�3���!?�R���@�/�c�ٿN��]-��@� VsE4@8�3���!?�R���@�/�c�ٿN��]-��@� VsE4@8�3���!?�R���@��ZȉٿUw���@���߫4@�_��!?pM����@��ZȉٿUw���@���߫4@�_��!?pM����@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�)��ٿ�?!����@����� 4@�fj�!?&�g��@�i �يٿǢ��_��@R��� 4@g����!?�{	���@���"هٿYQ3~LN�@���4@llx���!?����y�@���"هٿYQ3~LN�@���4@llx���!?����y�@���"هٿYQ3~LN�@���4@llx���!?����y�@GI����ٿ�q'~�@+���\4@��ߛϐ!?ܦQ4�@GI����ٿ�q'~�@+���\4@��ߛϐ!?ܦQ4�@GI����ٿ�q'~�@+���\4@��ߛϐ!?ܦQ4�@GI����ٿ�q'~�@+���\4@��ߛϐ!?ܦQ4�@GI����ٿ�q'~�@+���\4@��ߛϐ!?ܦQ4�@��i�҆ٿ?^�^a�@�^z�4@6%�-��!?�����@��i�҆ٿ?^�^a�@�^z�4@6%�-��!?�����@��i�҆ٿ?^�^a�@�^z�4@6%�-��!?�����@Q����ٿ"7|D';�@~���q4@�����!?m�P�B%�@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��rM%�ٿ@<[��8�@��p54@]�]��!?�
թt��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��|��ٿ��R�C�@��<ū4@�	h��!?AF�y��@��9yV�ٿ"�t�y�@��e��4@����ߐ!?Y1KJy�@��9yV�ٿ"�t�y�@��e��4@����ߐ!?Y1KJy�@��9yV�ٿ"�t�y�@��e��4@����ߐ!?Y1KJy�@����ٿ�N�@�\I��4@��Ʉ�!?����@����ٿ�N�@�\I��4@��Ʉ�!?����@����ٿ�N�@�\I��4@��Ʉ�!?����@����ٿ�N�@�\I��4@��Ʉ�!?����@����ٿ�N�@�\I��4@��Ʉ�!?����@f���؆ٿs6L��f�@�u^d4@A#/sc�!?ݙ�{9��@f���؆ٿs6L��f�@�u^d4@A#/sc�!?ݙ�{9��@f���؆ٿs6L��f�@�u^d4@A#/sc�!?ݙ�{9��@f���؆ٿs6L��f�@�u^d4@A#/sc�!?ݙ�{9��@f���؆ٿs6L��f�@�u^d4@A#/sc�!?ݙ�{9��@�$�:��ٿ���!��@��IB�4@��b�!?���[���@�$�:��ٿ���!��@��IB�4@��b�!?���[���@�$�:��ٿ���!��@��IB�4@��b�!?���[���@�%xN�ٿ�E9Il�@[��K4@NJ+V]�!?���b[�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@�BO�t�ٿ�����@Wm���4@�g#�2�!?��Y�%�@��~7�ٿ��p+�@vO_�4@��%~�!?S�r=��@��`ׄٿ		r��@��4@����!?�y�Ž��@��`ׄٿ		r��@��4@����!?�y�Ž��@3���Շٿ6 �D��@�Qq�4@�H���!?9�My�@3���Շٿ6 �D��@�Qq�4@�H���!?9�My�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@�y�X݌ٿ�^�H+�@��44@q���4�!?7����$�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@:�	O�ٿx��Б�@�2a�4@��D��!?��?�;�@����X�ٿ��N9���@�D}�4@��Fb�!?�h�}��@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@ߍa�o�ٿߣ�����@́�]�4@.sGM�!?��6���@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@�;�O�ٿ���]�@Z�U4x4@��2!Ӑ!?J6�+�@Q�oٿ�ֶ0���@����<4@��v���!?4�&Ձ��@Q�oٿ�ֶ0���@����<4@��v���!?4�&Ձ��@Q�oٿ�ֶ0���@����<4@��v���!?4�&Ձ��@Q�oٿ�ֶ0���@����<4@��v���!?4�&Ձ��@�ߨ���ٿ1l���@��ݽ4@E�1��!?�y�u�D�@�ߨ���ٿ1l���@��ݽ4@E�1��!?�y�u�D�@�ߨ���ٿ1l���@��ݽ4@E�1��!?�y�u�D�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@L����ٿ��ІA�@PW���4@4���Ґ!?<$�b�9�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@����ٿ�0��x��@�����4@	�Q��!?�f8x�@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@s�t,�ٿ̨@����@�̙�4@�����!?Aٌ `��@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���QO�ٿa�SZ�l�@rq���4@��xmސ!?�� }�O�@���ٿF�%�I��@�`^)�4@�����!?�����W�@���ٿF�%�I��@�`^)�4@�����!?�����W�@�6$FG�ٿ_�{	�@!��J	4@|�	���!?��i�+-�@�6$FG�ٿ_�{	�@!��J	4@|�	���!?��i�+-�@~�`s�ٿ!O�wUd�@�d���4@�R|Ȑ!?�]��'�@���__zٿ��*�k�@�&��4@��-���!?*U36��@���__zٿ��*�k�@�&��4@��-���!?*U36��@���__zٿ��*�k�@�&��4@��-���!?*U36��@���__zٿ��*�k�@�&��4@��-���!?*U36��@���__zٿ��*�k�@�&��4@��-���!?*U36��@���__zٿ��*�k�@�&��4@��-���!?*U36��@O����~ٿN���m@�@��җq4@"�1�!?�}N��%�@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@�+��ٿP�sq�Y�@�kk4@�ޠF�!?��n��@��ٿ�	�>��@-�oc4@�ۯ���!?�)���@���ڏٿUqM(%B�@��F4@��`ɳ�!?v����@���ڏٿUqM(%B�@��F4@��`ɳ�!?v����@��X�e�ٿ������@����"	4@�:�ʐ!?�]��8��@��X�e�ٿ������@����"	4@�:�ʐ!?�]��8��@��X�e�ٿ������@����"	4@�:�ʐ!?�]��8��@��?O��ٿc�+Kr��@�CCa4@+׹3��!?�T��
��@��?O��ٿc�+Kr��@�CCa4@+׹3��!?�T��
��@��?O��ٿc�+Kr��@�CCa4@+׹3��!?�T��
��@��?O��ٿc�+Kr��@�CCa4@+׹3��!?�T��
��@�Ts���ٿ��.��@�@�F��54@�͚�ِ!?�L1Sg��@F�H�̄ٿ������@ z��4@˦T�Ր!?LA��z��@F�H�̄ٿ������@ z��4@˦T�Ր!?LA��z��@F�H�̄ٿ������@ z��4@˦T�Ր!?LA��z��@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@Յ��Ćٿ�Й^�t�@�0n�4@b��~��!?9���h�@�A_��ٿ��k�֔�@ �	� 4@�����!?�j:߸��@�A_��ٿ��k�֔�@ �	� 4@�����!?�j:߸��@�A_��ٿ��k�֔�@ �	� 4@�����!?�j:߸��@�A_��ٿ��k�֔�@ �	� 4@�����!?�j:߸��@ZU��ٿ`L��1�@�M��Q4@�+���!?~��E�k�@ZU��ٿ`L��1�@�M��Q4@�+���!?~��E�k�@ZU��ٿ`L��1�@�M��Q4@�+���!?~��E�k�@�O�s��ٿ;�����@���4@b%���!?��2�3�@)G���ٿ01�N���@���f�4@!$&��!?� 7�@)G���ٿ01�N���@���f�4@!$&��!?� 7�@z��ڱ�ٿ�G,���@i�b�M4@�̀���!?�:�dB�@z��ڱ�ٿ�G,���@i�b�M4@�̀���!?�:�dB�@z��ڱ�ٿ�G,���@i�b�M4@�̀���!?�:�dB�@z��ڱ�ٿ�G,���@i�b�M4@�̀���!?�:�dB�@z��ڱ�ٿ�G,���@i�b�M4@�̀���!?�:�dB�@���كٿ�`��N��@Pl+�C4@es��!?ߘ��-Z�@���كٿ�`��N��@Pl+�C4@es��!?ߘ��-Z�@���كٿ�`��N��@Pl+�C4@es��!?ߘ��-Z�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@p^���ٿV�䉡�@�>j+4@ ԝ`~�!?��*h�@�W�Fr�ٿ�i���@��խw 4@X�\א!?'/�[��@�02n��ٿQ���\��@�r��54@X��=��!?��/d�@�02n��ٿQ���\��@�r��54@X��=��!?��/d�@�02n��ٿQ���\��@�r��54@X��=��!?��/d�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@�(�]�ٿ���s��@�?���4@O4��!?�<�G+�@et.��ٿj��j�	�@޺�R�4@������!?�n�bA��@et.��ٿj��j�	�@޺�R�4@������!?�n�bA��@1

�.ٿ��(��@>oc��4@�7�ݔ�!?�JP��@1

�.ٿ��(��@>oc��4@�7�ݔ�!?�JP��@1

�.ٿ��(��@>oc��4@�7�ݔ�!?�JP��@m�|��ٿ�[����@�Fp��4@�L䘐!?#CӤ��@w7�VU�ٿ�xF��@�E]Y� 4@;����!?pm��@w7�VU�ٿ�xF��@�E]Y� 4@;����!?pm��@w7�VU�ٿ�xF��@�E]Y� 4@;����!?pm��@w7�VU�ٿ�xF��@�E]Y� 4@;����!?pm��@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@�9�\�ٿ�Or����@�?C�� 4@<�AQ�!?f_Ni�@9�Ɔٿe���"��@v���4@IT���!?�@���@9�Ɔٿe���"��@v���4@IT���!?�@���@9�Ɔٿe���"��@v���4@IT���!?�@���@9�Ɔٿe���"��@v���4@IT���!?�@���@9�Ɔٿe���"��@v���4@IT���!?�@���@T�J��ٿ�`2���@>q��X4@]����!?E+����@O,Ĉ��ٿE��C|�@G�[U�4@Ӭo���!?h9���
�@O,Ĉ��ٿE��C|�@G�[U�4@Ӭo���!?h9���
�@O,Ĉ��ٿE��C|�@G�[U�4@Ӭo���!?h9���
�@O,Ĉ��ٿE��C|�@G�[U�4@Ӭo���!?h9���
�@O,Ĉ��ٿE��C|�@G�[U�4@Ӭo���!?h9���
�@���ٿ]�<9��@���4@�6��!?`k�"��@���ٿ]�<9��@���4@�6��!?`k�"��@���ٿ]�<9��@���4@�6��!?`k�"��@���6�ٿ'��_`��@����4@]��ʐ!?柲����@���6�ٿ'��_`��@����4@]��ʐ!?柲����@���6�ٿ'��_`��@����4@]��ʐ!?柲����@���6�ٿ'��_`��@����4@]��ʐ!?柲����@���6�ٿ'��_`��@����4@]��ʐ!?柲����@:���ٿ�F����@�Ȟ�i4@�_`���!?��jZ��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@e��u��ٿ�i��C�@k���4@Bw"�Ð!?*�&��@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@{3���ٿo� ���@��\�4@�!/&	�!?\�����@BX0�̇ٿ�;k(�F�@L{y_�4@�$�飐!?j��:[#�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@8�~i͇ٿ&>o�5�@2H%��4@�6���!?����ʤ�@9f�nO�ٿy���@A��4@�9��:�!?Gx�E*1�@9f�nO�ٿy���@A��4@�9��:�!?Gx�E*1�@9f�nO�ٿy���@A��4@�9��:�!?Gx�E*1�@Vώ��ٿ
�b��@�X��T4@�:�t��!?Պ9q8��@Vώ��ٿ
�b��@�X��T4@�:�t��!?Պ9q8��@Vώ��ٿ
�b��@�X��T4@�:�t��!?Պ9q8��@Vώ��ٿ
�b��@�X��T4@�:�t��!?Պ9q8��@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@��<�ٿ�L��@(�vT4@��E���!?�ݐROf�@���k�ٿ>���a�@_8A�K4@Xw�K��!?EK�o�@���k�ٿ>���a�@_8A�K4@Xw�K��!?EK�o�@���k�ٿ>���a�@_8A�K4@Xw�K��!?EK�o�@��|��ٿd���6��@�4��4@f��А!?}���S��@��|��ٿd���6��@�4��4@f��А!?}���S��@��|��ٿd���6��@�4��4@f��А!?}���S��@��|��ٿd���6��@�4��4@f��А!?}���S��@��|��ٿd���6��@�4��4@f��А!?}���S��@��|��ٿd���6��@�4��4@f��А!?}���S��@��:~�ٿ���/g��@�ɲt� 4@��S�̐!?�.}����@H����ٿ(g^����@�|�14@�h��!?= ��q�@H����ٿ(g^����@�|�14@�h��!?= ��q�@H����ٿ(g^����@�|�14@�h��!?= ��q�@H����ٿ(g^����@�|�14@�h��!?= ��q�@H����ٿ(g^����@�|�14@�h��!?= ��q�@�5m��ٿޟ�ۑO�@Q�A84@HP�:ѐ!?�{9�l��@�5m��ٿޟ�ۑO�@Q�A84@HP�:ѐ!?�{9�l��@�5m��ٿޟ�ۑO�@Q�A84@HP�:ѐ!?�{9�l��@�5m��ٿޟ�ۑO�@Q�A84@HP�:ѐ!?�{9�l��@֎���ٿ�����@A���3@s��y��!?�{;�X�@֎���ٿ�����@A���3@s��y��!?�{;�X�@o�p.�ٿ�͸���@͒⑊4@��c2Z�!?"���0�@o�p.�ٿ�͸���@͒⑊4@��c2Z�!?"���0�@o�p.�ٿ�͸���@͒⑊4@��c2Z�!?"���0�@�|@�ٿ��Ӆ:�@X�N|4@6��K��!?"·���@�|@�ٿ��Ӆ:�@X�N|4@6��K��!?"·���@�|@�ٿ��Ӆ:�@X�N|4@6��K��!?"·���@�|@�ٿ��Ӆ:�@X�N|4@6��K��!?"·���@$E�G�ٿ�(���@m�Ŀ#4@������!?t�4&R%�@$E�G�ٿ�(���@m�Ŀ#4@������!?t�4&R%�@��D���ٿ� ��@Ad��3@.ߐ!?g�6u��@��D���ٿ� ��@Ad��3@.ߐ!?g�6u��@��D���ٿ� ��@Ad��3@.ߐ!?g�6u��@��D���ٿ� ��@Ad��3@.ߐ!?g�6u��@��'�ٿJJH��[�@P�34@����!?oԀ���@�%&��ٿ�X��y�@y^hۖ4@Y�!?F��RI��@r����ٿB�gM�P�@���4@�� ~�!?E&n��@r����ٿB�gM�P�@���4@�� ~�!?E&n��@r����ٿB�gM�P�@���4@�� ~�!?E&n��@�,�_U�ٿ�e����@n�bk4@���g�!?~/��k �@�,�_U�ٿ�e����@n�bk4@���g�!?~/��k �@zSq�ٿ��ɱ���@�R �	4@���!?���^���@zSq�ٿ��ɱ���@�R �	4@���!?���^���@zSq�ٿ��ɱ���@�R �	4@���!?���^���@zSq�ٿ��ɱ���@�R �	4@���!?���^���@�M ��ٿ�L����@��*�
4@�tqTf�!?�h=��@�M ��ٿ�L����@��*�
4@�tqTf�!?�h=��@�M ��ٿ�L����@��*�
4@�tqTf�!?�h=��@�L ���ٿ1���¡�@�4��B4@WGi6��!?F�"�L�@�L ���ٿ1���¡�@�4��B4@WGi6��!?F�"�L�@�L ���ٿ1���¡�@�4��B4@WGi6��!?F�"�L�@�L ���ٿ1���¡�@�4��B4@WGi6��!?F�"�L�@F���ٿ@?�4sw�@��D6�4@8� ��!?s�^Ӎ��@F���ٿ@?�4sw�@��D6�4@8� ��!?s�^Ӎ��@F���ٿ@?�4sw�@��D6�4@8� ��!?s�^Ӎ��@F���ٿ@?�4sw�@��D6�4@8� ��!?s�^Ӎ��@F���ٿ@?�4sw�@��D6�4@8� ��!?s�^Ӎ��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@	i��ʍٿ�Hd��@r����4@	L��
�!?ߑ�1-��@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@���Fǉٿ2,���@� ��4@�@���!?����@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@=�΋�ٿȖ��@w�<Qr4@%��Ő!?ҢT��@_��2��ٿ��	��3�@'�I
�4@ioK���!?�}QG#l�@�p�d��ٿ>P��f2�@l�_��4@N�3y[�!?�Аi���@�p�d��ٿ>P��f2�@l�_��4@N�3y[�!?�Аi���@�p�d��ٿ>P��f2�@l�_��4@N�3y[�!?�Аi���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@A�%��ٿhe��-��@ma�<�4@�)i�[�!?�_�P���@�*��|�ٿ�#��N��@�Uk�4@y��:А!?�$����@�*��|�ٿ�#��N��@�Uk�4@y��:А!?�$����@�*��|�ٿ�#��N��@�Uk�4@y��:А!?�$����@�*��|�ٿ�#��N��@�Uk�4@y��:А!?�$����@�*��|�ٿ�#��N��@�Uk�4@y��:А!?�$����@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@Ny.�ٿn!�w)_�@�K���4@i�U�!?JӉ}q�@0kɣԆٿ(ĲX
��@Ά�4@�����!?���d��@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@{�C
�ٿJo4���@�w��A4@gЛ�!?�	_���@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�ʊٿ���DVS�@L���� 4@�^U\�!?�߉����@�10g*�ٿ��{���@G�m4@� �94�!?�\�Wo��@ߏc�B�ٿ�Y���@��e��4@-��5�!?\wt؏��@�t�/�ٿL��\8��@���c>4@�@ぐ!?�%}�@[�ɤ�ٿ���[��@�d_4@�� ��!?x��,, �@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@�!ퟠ�ٿƭ��x��@�˖>n4@Ma7��!?��V���@%�gҌٿ���e)<�@��(E4@�̥��!?>CE���@%�gҌٿ���e)<�@��(E4@�̥��!?>CE���@%�gҌٿ���e)<�@��(E4@�̥��!?>CE���@%�gҌٿ���e)<�@��(E4@�̥��!?>CE���@%�gҌٿ���e)<�@��(E4@�̥��!?>CE���@���S��ٿ<x,���@z��4@�PH��!?3ϙ	[6�@���S��ٿ<x,���@z��4@�PH��!?3ϙ	[6�@���S��ٿ<x,���@z��4@�PH��!?3ϙ	[6�@���S��ٿ<x,���@z��4@�PH��!?3ϙ	[6�@�>��ٿ��oy��@�V`��4@��'�!?P�η-��@�>��ٿ��oy��@�V`��4@��'�!?P�η-��@����bٿ����'b�@��^�,4@s�pҐ!?|��c6�@�X�ٿ�`�����@���&L4@0ap��!?T-�Q���@�X�ٿ�`�����@���&L4@0ap��!?T-�Q���@�X�ٿ�`�����@���&L4@0ap��!?T-�Q���@�X�ٿ�`�����@���&L4@0ap��!?T-�Q���@�X�ٿ�`�����@���&L4@0ap��!?T-�Q���@J˕��ٿ*F�k-��@�5�Y'4@����!?�$�����@J˕��ٿ*F�k-��@�5�Y'4@����!?�$�����@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@쎿��ٿ���j��@_Wn1	4@en���!?��RR�@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@.+z]��ٿK�M���@jv��/4@T�i�!?�+�v��@�$�ވٿ�ql(`��@:#A��4@܀��ݐ!?>���"�@�$�ވٿ�ql(`��@:#A��4@܀��ݐ!?>���"�@�$�ވٿ�ql(`��@:#A��4@܀��ݐ!?>���"�@bK4���ٿ�ekR���@����4@i��f��!?\ˎr,�@bK4���ٿ�ekR���@����4@i��f��!?\ˎr,�@bK4���ٿ�ekR���@����4@i��f��!?\ˎr,�@bK4���ٿ�ekR���@����4@i��f��!?\ˎr,�@bK4���ٿ�ekR���@����4@i��f��!?\ˎr,�@��5*��ٿ��B%G��@5���|4@:��b��!?|�a����@��5*��ٿ��B%G��@5���|4@:��b��!?|�a����@��5*��ٿ��B%G��@5���|4@:��b��!?|�a����@��5*��ٿ��B%G��@5���|4@:��b��!?|�a����@��5*��ٿ��B%G��@5���|4@:��b��!?|�a����@��Jk��ٿ.��H6�@O�s�H4@�v"Њ�!?����0>�@��Jk��ٿ.��H6�@O�s�H4@�v"Њ�!?����0>�@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@�
Ĭٿ��&�&�@bM��4@i��㳐!?�1GC��@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@E�s�ٿ�6�@	��?44@�_&��!?��m���@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@K�9ն�ٿ���HR�@(:ta%4@
TLO�!?�����@��� ��ٿ�ŏ���@�*}� 4@Sshɐ!?��!E,��@��� ��ٿ�ŏ���@�*}� 4@Sshɐ!?��!E,��@��� ��ٿ�ŏ���@�*}� 4@Sshɐ!?��!E,��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@���~��ٿ�(��z�@�#_�&4@qI�Ґ!?�*�\0��@��^��ٿi�6%i�@��z� 4@��=�6�!?�j��b/�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@�gWw��ٿMh� �S�@l��-t4@"��$�!?�k�\�[�@Cd�B�|ٿ-y`�V�@�C~��4@a��/�!?�E�D���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@��E{ٿg���@���4@�n��ؐ!?3�C���@�����xٿ�s�$M�@�aE��4@��k۾�!?�����@���B�yٿ�Z2��/�@A扗�4@�қ�!?"��@��@���B�yٿ�Z2��/�@A扗�4@�қ�!?"��@��@���B�yٿ�Z2��/�@A扗�4@�қ�!?"��@��@���B�yٿ�Z2��/�@A扗�4@�қ�!?"��@��@���B�yٿ�Z2��/�@A扗�4@�қ�!?"��@��@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@�x#�yٿ��p��4�@���4@;qȢ��!?�~4%�-�@ш�qq}ٿ���SB��@��w��4@4fȐ!?y�l���@ш�qq}ٿ���SB��@��w��4@4fȐ!?y�l���@ш�qq}ٿ���SB��@��w��4@4fȐ!?y�l���@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@��;�ٿ[�p	��@�U�Q�4@0!�ΐ!?~P�n��@1���уٿe\�U5��@���+4@d׌�ܐ!?`C��r�@1���уٿe\�U5��@���+4@d׌�ܐ!?`C��r�@1���уٿe\�U5��@���+4@d׌�ܐ!?`C��r�@1���уٿe\�U5��@���+4@d׌�ܐ!?`C��r�@1���уٿe\�U5��@���+4@d׌�ܐ!?`C��r�@yΣg��ٿFwBC:��@]��4@�]����!?�d���@yΣg��ٿFwBC:��@]��4@�]����!?�d���@yΣg��ٿFwBC:��@]��4@�]����!?�d���@yΣg��ٿFwBC:��@]��4@�]����!?�d���@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@Mr�w��ٿ�cS0/��@�x���4@ө.,А!?�Ϸ=Vw�@���aH�ٿm��y���@"҃��4@�6}��!?�?��<I�@���aH�ٿm��y���@"҃��4@�6}��!?�?��<I�@Қ��%�ٿ���	���@��4@;�c�֐!?;ˀ�9��@� *���ٿn9 �@���#�4@���UՐ!?����u��@� *���ٿn9 �@���#�4@���UՐ!?����u��@� *���ٿn9 �@���#�4@���UՐ!?����u��@� *���ٿn9 �@���#�4@���UՐ!?����u��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@Đ�c��ٿm��~���@�J��#	4@I��ו�!?d��6��@t����ٿȵ��U�@ƙ��4@��5�!?�?{����@t����ٿȵ��U�@ƙ��4@��5�!?�?{����@�lR�zٿ�#rL���@�9=14@6ր�̐!?��'ov
�@�lR�zٿ�#rL���@�9=14@6ր�̐!?��'ov
�@�lR�zٿ�#rL���@�9=14@6ր�̐!?��'ov
�@�lR�zٿ�#rL���@�9=14@6ր�̐!?��'ov
�@��K6�xٿ%)�Qţ�@9^ʡk4@Rnxi��!?����q�@��K6�xٿ%)�Qţ�@9^ʡk4@Rnxi��!?����q�@{�6*�ٿ�"x����@�bT
 4@-�#O��!?���.l�@{�6*�ٿ�"x����@�bT
 4@-�#O��!?���.l�@{�6*�ٿ�"x����@�bT
 4@-�#O��!?���.l�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@𐒘��ٿ0���5S�@+��4@n6y��!?H����]�@�pu��ٿY9�A��@Dᗚ4@>��!?:�|AD�@�pu��ٿY9�A��@Dᗚ4@>��!?:�|AD�@�pu��ٿY9�A��@Dᗚ4@>��!?:�|AD�@�pu��ٿY9�A��@Dᗚ4@>��!?:�|AD�@��F��}ٿy	����@��u�4@}�YIʐ!?�!>�{%�@��F��}ٿy	����@��u�4@}�YIʐ!?�!>�{%�@��F��}ٿy	����@��u�4@}�YIʐ!?�!>�{%�@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@��oٿ3���V��@N?bqi4@�w����!?.wZ$��@P�i̈́ٿ�n)N��@���&54@�4�ѐ!?+,����@P�i̈́ٿ�n)N��@���&54@�4�ѐ!?+,����@P�i̈́ٿ�n)N��@���&54@�4�ѐ!?+,����@P�i̈́ٿ�n)N��@���&54@�4�ѐ!?+,����@���|�ٿ�R�K�y�@k���t4@���g�!?h�/�J��@���|�ٿ�R�K�y�@k���t4@���g�!?h�/�J��@���|�ٿ�R�K�y�@k���t4@���g�!?h�/�J��@���|�ٿ�R�K�y�@k���t4@���g�!?h�/�J��@���|�ٿ�R�K�y�@k���t4@���g�!?h�/�J��@n_r�Јٿ��J�@TT�ؠ4@Y��2�!?'9�%_�@n_r�Јٿ��J�@TT�ؠ4@Y��2�!?'9�%_�@n_r�Јٿ��J�@TT�ؠ4@Y��2�!?'9�%_�@���u�ٿ�����@��T��4@ ���8�!?�}�Vx�@���u�ٿ�����@��T��4@ ���8�!?�}�Vx�@��q�x~ٿP�ʸ��@���ؗ4@�y`'�!?�(O��@���_~ٿw�.�@	"f�4@~k�{�!?�>[����@���_~ٿw�.�@	"f�4@~k�{�!?�>[����@���_~ٿw�.�@	"f�4@~k�{�!?�>[����@�b�Wn�ٿ�K�La$�@O`�<4@���@$�!?���AQ�@�b�Wn�ٿ�K�La$�@O`�<4@���@$�!?���AQ�@�G@;�ٿkEk
s��@���� 4@1�E��!?'l��yM�@�G@;�ٿkEk
s��@���� 4@1�E��!?'l��yM�@;�]��ٿđ�ȟ�@�Ѷ� 4@��_FҐ!?���ٚ�@;�]��ٿđ�ȟ�@�Ѷ� 4@��_FҐ!?���ٚ�@;�]��ٿđ�ȟ�@�Ѷ� 4@��_FҐ!?���ٚ�@;�]��ٿđ�ȟ�@�Ѷ� 4@��_FҐ!?���ٚ�@;�]��ٿđ�ȟ�@�Ѷ� 4@��_FҐ!?���ٚ�@����{ٿ���&��@���e�4@��ke�!?b�D�;O�@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@��Wىٿ=b����@��i�4@?o\�Ԑ!?������@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@B��ٿ��Z��@M+�4@�M���!?bg�����@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@��W�ٿ�w�q��@�/�k�4@�7�א!?U �3���@���T�ٿ���铘�@��/��4@<!&K��!?<�G���@Ww�L�ٿi�ך�@�5��	4@1�)��!?�v&���@>���]�ٿ=}�B$��@Gn�64@Z�]��!?r˫
��@>���]�ٿ=}�B$��@Gn�64@Z�]��!?r˫
��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@��U�čٿ���!�c�@4�9s�4@͞%��!?}�eG��@�y�uI�ٿ_T�q)�@?Q�"4@`��'�!?��D���@�y�uI�ٿ_T�q)�@?Q�"4@`��'�!?��D���@�y�uI�ٿ_T�q)�@?Q�"4@`��'�!?��D���@�y�uI�ٿ_T�q)�@?Q�"4@`��'�!?��D���@e�Pˆٿb�	ա��@0"}4@�ӕ/�!?c�C�|�@e�Pˆٿb�	ա��@0"}4@�ӕ/�!?c�C�|�@e�Pˆٿb�	ա��@0"}4@�ӕ/�!?c�C�|�@e�Pˆٿb�	ա��@0"}4@�ӕ/�!?c�C�|�@e�Pˆٿb�	ա��@0"}4@�ӕ/�!?c�C�|�@�u�T��ٿL��Ъ�@�e"F4@ZgZ�J�!?��ׅ(I�@�u�T��ٿL��Ъ�@�e"F4@ZgZ�J�!?��ׅ(I�@�u�T��ٿL��Ъ�@�e"F4@ZgZ�J�!?��ׅ(I�@�u�T��ٿL��Ъ�@�e"F4@ZgZ�J�!?��ׅ(I�@&Wn��ٿm_����@��O�{4@��>(�!?O	1V�
�@&Wn��ٿm_����@��O�{4@��>(�!?O	1V�
�@&Wn��ٿm_����@��O�{4@��>(�!?O	1V�
�@&Wn��ٿm_����@��O�{4@��>(�!?O	1V�
�@�gR�ٿ�r ��@�D@�k4@���F �!?>�����@�gR�ٿ�r ��@�D@�k4@���F �!?>�����@�gR�ٿ�r ��@�D@�k4@���F �!?>�����@�gR�ٿ�r ��@�D@�k4@���F �!?>�����@�42��ٿbX8'��@�d�4@J���!?!��_5\�@�42��ٿbX8'��@�d�4@J���!?!��_5\�@�42��ٿbX8'��@�d�4@J���!?!��_5\�@�42��ٿbX8'��@�d�4@J���!?!��_5\�@�42��ٿbX8'��@�d�4@J���!?!��_5\�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@���2��ٿ��y��@�}��2 4@�����!?�%&�@Q�{�f�ٿ��Mvw�@��	�4@��Ō�!?a謧�@Q�{�f�ٿ��Mvw�@��	�4@��Ō�!?a謧�@��-.�ٿ���˨l�@(w�HA4@E�=��!?o=Y5�@��-.�ٿ���˨l�@(w�HA4@E�=��!?o=Y5�@��-.�ٿ���˨l�@(w�HA4@E�=��!?o=Y5�@��-.�ٿ���˨l�@(w�HA4@E�=��!?o=Y5�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@��aĂ�ٿr�|���@�%Q�C4@v!��L�!?�JP��.�@t)Nٿ�)ӆ
�@3��4@}5��|�!?�㖬k��@t)Nٿ�)ӆ
�@3��4@}5��|�!?�㖬k��@t)Nٿ�)ӆ
�@3��4@}5��|�!?�㖬k��@t)Nٿ�)ӆ
�@3��4@}5��|�!?�㖬k��@�E�%�ٿc�TQb�@�6kb4@6�hĐ!?���#O��@�N�y�ٿw\�9�>�@`���4@{�wYߐ!?���d���@�N�y�ٿw\�9�>�@`���4@{�wYߐ!?���d���@�N�y�ٿw\�9�>�@`���4@{�wYߐ!?���d���@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@aL�櫂ٿ������@�w�J4@�%E�ΐ!?�d��K#�@S�3�B�ٿ*����@Ǜ��44@��`�!?���J6�@S�3�B�ٿ*����@Ǜ��44@��`�!?���J6�@S�3�B�ٿ*����@Ǜ��44@��`�!?���J6�@S�3�B�ٿ*����@Ǜ��44@��`�!?���J6�@�,��ٿU���{�@�By�4@P�e�ː!?Pp�Me�@�,��ٿU���{�@�By�4@P�e�ː!?Pp�Me�@(��?ɎٿH.;�:�@ވKp4@T�U�!?ǹ��F�@(��?ɎٿH.;�:�@ވKp4@T�U�!?ǹ��F�@(��?ɎٿH.;�:�@ވKp4@T�U�!?ǹ��F�@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@��[��ٿ5��_�f�@� ��=4@
Y ���!?��y)��@Թ�Άٿ:�>�S�@c]�#4@ZnMW�!?�گ�f�@��[��ٿ�M??���@�6�@4@��Omѐ!?��#ڶ�@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@����ٿ�'�<�p�@��s�4@o�
<А!?������@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@�Q^7��ٿ��3�wi�@i��af4@�c��!?ٓ5��@)Ż�ٿ��L���@8]xw4@0h��!?>��g�@)Ż�ٿ��L���@8]xw4@0h��!?>��g�@���ٿ��B�dj�@��[.�	4@ʥ�N��!?���:=�@���ٿ��B�dj�@��[.�	4@ʥ�N��!?���:=�@���ٿ��B�dj�@��[.�	4@ʥ�N��!?���:=�@���ٿ��B�dj�@��[.�	4@ʥ�N��!?���:=�@������ٿ{�B+��@v/Lq4@��{��!?l�X��'�@������ٿ{�B+��@v/Lq4@��{��!?l�X��'�@��=��ٿ�o��۱�@=�Y\�4@{����!?z��{��@��=��ٿ�o��۱�@=�Y\�4@{����!?z��{��@��=��ٿ�o��۱�@=�Y\�4@{����!?z��{��@���}#�ٿ�W�e�@P?��4@Lѐ!?�,R����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@�2����ٿ�v�#��@��L4@L/�驐!?}9����@kE��ٿ�k86�s�@컯�I4@(��!?�9\���@kE��ٿ�k86�s�@컯�I4@(��!?�9\���@���-~ٿ�T��~��@������3@��01�!??�We�Y�@!��ٿlԽ)L�@ێ��-�3@��쩐!?����! �@�t�Íٿ�tt�u�@25��$4@k`����!?,Rsd�C�@�t�Íٿ�tt�u�@25��$4@k`����!?,Rsd�C�@�L�ٿ9fڒ�;�@*[�l4@���Ա�!?���q�@�L�ٿ9fڒ�;�@*[�l4@���Ա�!?���q�@�L�ٿ9fڒ�;�@*[�l4@���Ա�!?���q�@��4G�ٿy�,��@3�p�u4@�g ���!?K�$���@��4G�ٿy�,��@3�p�u4@�g ���!?K�$���@��4G�ٿy�,��@3�p�u4@�g ���!?K�$���@��4G�ٿy�,��@3�p�u4@�g ���!?K�$���@J��Ԏ~ٿW��t���@̓���4@�bvn��!?���k?�@J��Ԏ~ٿW��t���@̓���4@�bvn��!?���k?�@�1L�!�ٿ�v��@�+b�4@a���{�!?a��@�;�@�1L�!�ٿ�v��@�+b�4@a���{�!?a��@�;�@�1L�!�ٿ�v��@�+b�4@a���{�!?a��@�;�@�1L�!�ٿ�v��@�+b�4@a���{�!?a��@�;�@[v,{�ٿX��?��@���ܤ4@^���!?�!�m�@[v,{�ٿX��?��@���ܤ4@^���!?�!�m�@[v,{�ٿX��?��@���ܤ4@^���!?�!�m�@[v,{�ٿX��?��@���ܤ4@^���!?�!�m�@v�Ņ�ٿ	q�4V��@g�4W\4@��zl��!?K�g�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@��e;\�ٿ'�d���@���H4@^ab�!?�G*�AG�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@���MR�ٿ��2SE��@�$�!C4@~�؞�!?�\�-�}�@�HQyO�ٿ�/5��@6��4@ ȴ��!?�v�e��@�HQyO�ٿ�/5��@6��4@ ȴ��!?�v�e��@�HQyO�ٿ�/5��@6��4@ ȴ��!?�v�e��@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�P)b�ٿ@����@�&�>#4@�W���!?i�y3�-�@�RlG�ٿl�,��@G��(4@�jƍ�!?Z�J�iu�@�RlG�ٿl�,��@G��(4@�jƍ�!?Z�J�iu�@�RlG�ٿl�,��@G��(4@�jƍ�!?Z�J�iu�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@C ��܂ٿw��ߕ
�@�̰S4@O����!?OKr=�@.�Vĩ�ٿ�z7���@�e�\4@�9���!?�Y&���@�{g��ٿ,���$�@U��e4@��淎�!?�~1��@}}�^�ٿ���|���@K�Qȶ4@̙��!?*��|���@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@���ׂٿ�6#����@�9%74@\MZ˚�!?n�'P�@XB%�M{ٿ���@M�?�4@SBy"��!?�\�?5�@XB%�M{ٿ���@M�?�4@SBy"��!?�\�?5�@XB%�M{ٿ���@M�?�4@SBy"��!?�\�?5�@XB%�M{ٿ���@M�?�4@SBy"��!?�\�?5�@`���ׂٿy�m5y��@�o�24@_���v�!?�q%����@`���ׂٿy�m5y��@�o�24@_���v�!?�q%����@`���ׂٿy�m5y��@�o�24@_���v�!?�q%����@r���ٿL��� X�@~�����3@.�,!?�eŸ���@2X>%�ٿ Qt�(`�@���A�3@ �&�!?^#�"�@2X>%�ٿ Qt�(`�@���A�3@ �&�!?^#�"�@2X>%�ٿ Qt�(`�@���A�3@ �&�!?^#�"�@2X>%�ٿ Qt�(`�@���A�3@ �&�!?^#�"�@2X>%�ٿ Qt�(`�@���A�3@ �&�!?^#�"�@����ٿݡT����@��S 4@&��V��!?��Ն;��@��ծ��ٿ�_�@���" 4@h�ҁΐ!?:B�,��@��ծ��ٿ�_�@���" 4@h�ҁΐ!?:B�,��@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�;��ٿ�	��Y��@����4@r�y���!?���M���@�z��*�ٿ�XlO^��@˗��l4@�"N��!?Q���4��@�z��*�ٿ�XlO^��@˗��l4@�"N��!?Q���4��@�z��*�ٿ�XlO^��@˗��l4@�"N��!?Q���4��@�IF
��ٿ�.�h̨�@bb��v4@)U�} �!?Q����@]H�~ٿ�׀���@uL5j4@�E�	�!?�tN�!�@]H�~ٿ�׀���@uL5j4@�E�	�!?�tN�!�@]H�~ٿ�׀���@uL5j4@�E�	�!?�tN�!�@]H�~ٿ�׀���@uL5j4@�E�	�!?�tN�!�@�yZ,s�ٿz�̮��@s���4@=-��!?��t�Y�@�yZ,s�ٿz�̮��@s���4@=-��!?��t�Y�@g(�@ٿ
����@3�5�4@^h�x��!?��l+N�@7�Jah}ٿ�y�&>�@�1��H4@��v�Ȑ!?�;�(?��@�&�i�zٿ��h��@k�y�4@W���!?x����@?ZFeٿ�ٿ����@�����	4@�ڐ!?$�?r"u�@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@��J�~ٿ�;m��
�@��e�4@y�͊��!?K.�Y��@c�j\}ٿ�;�U��@��_��4@��a�ِ!?�f"����@c�j\}ٿ�;�U��@��_��4@��a�ِ!?�f"����@��nC&}ٿ�J՞�@\���*4@V���̐!?X������@��nC&}ٿ�J՞�@\���*4@V���̐!?X������@��nC&}ٿ�J՞�@\���*4@V���̐!?X������@_��P�ٿ�!`�I�@��5$4@���Ð!?j�w�h��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@;�&�ٿd	�Ɠ�@��qd�4@���e�!?��L��@�Y��ٿ�X{�l��@�Q�#4@ܞ����!?{��ʒ�@��5�ٿ�_�1�F�@��Ea4@�-��!?df~ �@��snU�ٿ{��F���@��&4@W�{�d�!?��V7�@o R�D�ٿںD5��@`��4@W��!?|�W�@o R�D�ٿںD5��@`��4@W��!?|�W�@��g�ٿ)��=(��@1�|�4@� Sﳐ!?%��`��@���
Ȇٿ֘���@�� 4@C��Ð!?���'d�@���
Ȇٿ֘���@�� 4@C��Ð!?���'d�@ڮ��ōٿ�>� R��@���0��3@�nOo��!?����(��@ڮ��ōٿ�>� R��@���0��3@�nOo��!?����(��@ڮ��ōٿ�>� R��@���0��3@�nOo��!?����(��@Z�S�X�ٿf�f!f��@��D�'4@z�}w��!?ە���
�@<N\U��ٿ�[P>�@j��c;4@�G�!��!?"�2�U�@<N\U��ٿ�[P>�@j��c;4@�G�!��!?"�2�U�@<N\U��ٿ�[P>�@j��c;4@�G�!��!?"�2�U�@&W���ٿؕ5�^��@u��|=4@��;ِ!?ɞ���o�@&W���ٿؕ5�^��@u��|=4@��;ِ!?ɞ���o�@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�'��ٿu�H��3�@���Y4@�C]���!?K��8��@�4�ٿ��#��@�����4@R��|��!?�R���@�4�ٿ��#��@�����4@R��|��!?�R���@�4�ٿ��#��@�����4@R��|��!?�R���@�4�ٿ��#��@�����4@R��|��!?�R���@�4�ٿ��#��@�����4@R��|��!?�R���@�4�ٿ��#��@�����4@R��|��!?�R���@�b$�~ٿ5�G�{�@�Yʏ� 4@��g֐!?��>�%�@��˪R�ٿ�J.����@�N�44@��g|"�!?��ܰ�s�@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@���ٿ��h#�@�\�(l4@MnFh�!?Hn��]��@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@6�ٿ?�&��@��.��4@�
����!?H	�jz1�@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@�:��}ٿ=C�$��@��)��4@�eH���!?�j;��@LbÒ��ٿplH�s��@yl��L4@$�ݻ��!?��V5��@LbÒ��ٿplH�s��@yl��L4@$�ݻ��!?��V5��@LbÒ��ٿplH�s��@yl��L4@$�ݻ��!?��V5��@���+�ٿ�g����@R O5V4@Fv�ꤐ!?�]���@�9��ٿ3��9�@*�@ 4@rc����!?�����@�>�}p�ٿ�d�-��@��
J4@/��g��!?B
W�[�@�>�}p�ٿ�d�-��@��
J4@/��g��!?B
W�[�@�>�}p�ٿ�d�-��@��
J4@/��g��!?B
W�[�@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�=��"�ٿ*��w���@�%���4@:~���!?E�X�z��@�b��]�ٿ�����@����4@�7S���!?��y���@�?���ٿ�XI��@� 64@��*~�!?��f�)�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@��ڙ�ٿ6��4��@��wB4@9�Y��!?�q�(�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@j~�U�ٿ������@/�#j&4@�|k��!?�\Hz�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@Y�ނٿױY)��@'�tX44@fi�r��!?:(�@�@�����ٿ�e�U ��@Ռx4@tq��t�!?�:5>.�@�����ٿ�e�U ��@Ռx4@tq��t�!?�:5>.�@�����ٿ�e�U ��@Ռx4@tq��t�!?�:5>.�@�����ٿ�e�U ��@Ռx4@tq��t�!?�:5>.�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@s�J:�}ٿeί��@9�X~�4@���>��!?U�B;y�@��xٿT9�"��@��zzs4@e�ߐ!?�����C�@��xٿT9�"��@��zzs4@e�ߐ!?�����C�@��xٿT9�"��@��zzs4@e�ߐ!?�����C�@��xٿT9�"��@��zzs4@e�ߐ!?�����C�@�x�ٿ'��@���@����4@�Qmq��!?�����@�b�0�ٿ�MT�@��#:4@8K�\�!?�����@�b�0�ٿ�MT�@��#:4@8K�\�!?�����@�b�0�ٿ�MT�@��#:4@8K�\�!?�����@�b�0�ٿ�MT�@��#:4@8K�\�!?�����@�DNٿ� ����@
\�24@��	n�!?V(��@�DNٿ� ����@
\�24@��	n�!?V(��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@���Ã�ٿ�AEEX��@�L���4@�P娐!?8Wٕy��@�Ew��ٿ���M��@����<4@�<���!?J��A�@��^tD�ٿ>�����@�Q� 4@�Ž
�!?��x[�M�@��^tD�ٿ>�����@�Q� 4@�Ž
�!?��x[�M�@��^tD�ٿ>�����@�Q� 4@�Ž
�!?��x[�M�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@�HA~ٿﺙ�s=�@��JC��3@��h���!?�f�2�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@1�Y��ٿ��K���@i���4@,��f�!?ΚA�ra�@2��g��ٿ��P��@���C;4@�4���!?d垥���@2��g��ٿ��P��@���C;4@�4���!?d垥���@�#�쳇ٿ�>~q��@ӎBQx 4@�A� ��!?C`�{[��@�#�쳇ٿ�>~q��@ӎBQx 4@�A� ��!?C`�{[��@�#�쳇ٿ�>~q��@ӎBQx 4@�A� ��!?C`�{[��@�#�쳇ٿ�>~q��@ӎBQx 4@�A� ��!?C`�{[��@���Vٿ��w	&�@�ȷ?4@ǋ��ΐ!?��i����@���Vٿ��w	&�@�ȷ?4@ǋ��ΐ!?��i����@���Vٿ��w	&�@�ȷ?4@ǋ��ΐ!?��i����@��t�|ٿ5k�N�@����4@�/�ڝ�!?����T�@�iV�}�ٿ(g�p���@hZ5�L4@i@�F�!?�s~����@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�{[Dn�ٿ� ��@�;vT�4@kPQ�!?��V�\v�@�̰G]�ٿ�ڤT�@�p�L4@M+y�l�!?�=#�w��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@��+�ٿ�P�&g�@"��54@��w��!?�abd��@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@jU��ٿA�����@��f��4@�0���!?m��so�@z�)0|ٿ�#�s���@��\m;4@B�ni �!?}%g��_�@�ʐ��ٿH"� -�@� ��4@A'���!?�&��~�@�ʐ��ٿH"� -�@� ��4@A'���!?�&��~�@�ʐ��ٿH"� -�@� ��4@A'���!?�&��~�@�ʐ��ٿH"� -�@� ��4@A'���!?�&��~�@������ٿ�Ks?�@���S�4@b��O��!?����6�@������ٿ�Ks?�@���S�4@b��O��!?����6�@wU��i�ٿ���xQ�@������3@�ݥ:��!?FbU����@wU��i�ٿ���xQ�@������3@�ݥ:��!?FbU����@wU��i�ٿ���xQ�@������3@�ݥ:��!?FbU����@wU��i�ٿ���xQ�@������3@�ݥ:��!?FbU����@wU��i�ٿ���xQ�@������3@�ݥ:��!?FbU����@q�VgM�ٿ�d�w"x�@,\q�l4@p6 �L�!?��a���@q�VgM�ٿ�d�w"x�@,\q�l4@p6 �L�!?��a���@q�VgM�ٿ�d�w"x�@,\q�l4@p6 �L�!?��a���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@����K�ٿ����f�@w�q���3@}snO��!?���:���@�4Cu"�ٿ$�ح-��@�5∼�3@ �i.�!?�t���@�4Cu"�ٿ$�ح-��@�5∼�3@ �i.�!?�t���@�4Cu"�ٿ$�ح-��@�5∼�3@ �i.�!?�t���@����4�ٿ����@��4@QY��!�!?#�#�a�@E��ٿU=��)��@�S�F9 4@'ϧ��!? �����@E��ٿU=��)��@�S�F9 4@'ϧ��!? �����@E��ٿU=��)��@�S�F9 4@'ϧ��!? �����@E��ٿU=��)��@�S�F9 4@'ϧ��!? �����@E��ٿU=��)��@�S�F9 4@'ϧ��!? �����@ȷ�b@�ٿ_(~K~�@m?o�4@�Y ���!?�?�P��@�B��΋ٿ���8�}�@�J�]�4@^����!?��x,��@�B��΋ٿ���8�}�@�J�]�4@^����!?��x,��@|���K�ٿ��Φ��@�|4@'+#z�!?WA�4��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@��=i��ٿ3���d�@��:4@�%�8��!?��~��@R�$X�ٿM@!���@��_�4@�R�~�!?�$�[���@R�$X�ٿM@!���@��_�4@�R�~�!?�$�[���@V�|��ٿ��6H��@"��74@!�m�`�!?j^�W��@��:a��ٿ3���@��C4@Ï(��!?�����7�@���h�ٿ�p*퓋�@�Y�E�4@2����!?sW�7��@���h�ٿ�p*퓋�@�Y�E�4@2����!?sW�7��@���h�ٿ�p*퓋�@�Y�E�4@2����!?sW�7��@���h�ٿ�p*퓋�@�Y�E�4@2����!?sW�7��@���h�ٿ�p*퓋�@�Y�E�4@2����!?sW�7��@����ٿ�j���@5�RΆ4@���!?�,8�v��@ju?���ٿ�E��U��@�H�s4@����!?�a��9:�@ju?���ٿ�E��U��@�H�s4@����!?�a��9:�@ju?���ٿ�E��U��@�H�s4@����!?�a��9:�@ju?���ٿ�E��U��@�H�s4@����!?�a��9:�@6oe":ٿ�wR���@e�n4@N�����!?�N�}�@��kB�ٿ�7k���@��)4@�^@子!?;��j���@��kB�ٿ�7k���@��)4@�^@子!?;��j���@��kB�ٿ�7k���@��)4@�^@子!?;��j���@�l[x�ٿ��(!+��@i.}	4@)BTՐ!?���Lo0�@�	�ׄٿ��%	��@��24@ܗ%/C�!?k�Rq5��@�	�ׄٿ��%	��@��24@ܗ%/C�!?k�Rq5��@�	�ׄٿ��%	��@��24@ܗ%/C�!?k�Rq5��@�	�ׄٿ��%	��@��24@ܗ%/C�!?k�Rq5��@�	�ׄٿ��%	��@��24@ܗ%/C�!?k�Rq5��@8<��ٿ�%�:���@[rV��4@����!?\{�8���@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@��	��ٿ�.W�U�@ЋD��4@/(=�>�!?�Z�x&��@K�q�d�ٿ.�E7@�@�tݢ4@�O��>�!?��1��@���� �ٿ������@�
4@�5����!?�X�S1��@��X��ٿ�蠌��@�o���
4@h��퐐!?w�[�@;?ԥ�ٿ�iC�ϯ�@.|�<4@�l0.��!?&	E��@;?ԥ�ٿ�iC�ϯ�@.|�<4@�l0.��!?&	E��@;?ԥ�ٿ�iC�ϯ�@.|�<4@�l0.��!?&	E��@��0�ʂٿY�j~��@Z 4@+$���!?g�h~�@��0�ʂٿY�j~��@Z 4@+$���!?g�h~�@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�F�4�ٿ��ת��@�A��54@}�"��!?��1N���@�!��S�ٿ:�fP��@i*��4@")!?�\��bB�@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@
Ba{v�ٿ~v�/e�@�h�@4@ p7�!?I+�m��@,�>A�ٿ��t��Z�@H�}.@4@zJ�(��!?���qi�@,�>A�ٿ��t��Z�@H�}.@4@zJ�(��!?���qi�@yo�h��ٿ+��r�R�@ȼ�G4@\~֍�!? 	�h��@yo�h��ٿ+��r�R�@ȼ�G4@\~֍�!? 	�h��@�.h}ٿ��yx��@��ۣ4@�5>��!?/Q����@�.h}ٿ��yx��@��ۣ4@�5>��!?/Q����@�.h}ٿ��yx��@��ۣ4@�5>��!?/Q����@�.h}ٿ��yx��@��ۣ4@�5>��!?/Q����@�.h}ٿ��yx��@��ۣ4@�5>��!?/Q����@-7��ٿd�}s���@��d� 4@ő!Ɛ!?���o�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ ��=#�ٿݝye���@#T�E4@�º�!?�2E3�@ӻ.�ٿAż��@��Y04@�S]0��!?k�=����@ӻ.�ٿAż��@��Y04@�S]0��!?k�=����@ӻ.�ٿAż��@��Y04@�S]0��!?k�=����@	>&�ٿh&)��^�@�@B}�4@w.�L�!?���q���@	>&�ٿh&)��^�@�@B}�4@w.�L�!?���q���@	>&�ٿh&)��^�@�@B}�4@w.�L�!?���q���@�8���ٿ���F�j�@���~4@P��仐!?�_v����@�8���ٿ���F�j�@���~4@P��仐!?�_v����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@�r�W�ٿ�Q��x��@��ט4@U�� ��!?Mմ����@f�)l4�ٿE��3���@dj��W4@z�ֆ��!?:���s�@ NH��ٿ������@���� 4@}1C�!?���.`u�@ NH��ٿ������@���� 4@}1C�!?���.`u�@�B�ٿ��ʽ�@:Bv�K4@���i�!?�V���@�B�ٿ��ʽ�@:Bv�K4@���i�!?�V���@�B�ٿ��ʽ�@:Bv�K4@���i�!?�V���@H����ٿ�E��"�@��=�~4@��޹8�!?D��>���@H����ٿ�E��"�@��=�~4@��޹8�!?D��>���@H����ٿ�E��"�@��=�~4@��޹8�!?D��>���@H����ٿ�E��"�@��=�~4@��޹8�!?D��>���@�t����ٿ�ؿ�١�@��414@�Gu��!?i�ܷE<�@�t����ٿ�ؿ�١�@��414@�Gu��!?i�ܷE<�@�t����ٿ�ؿ�١�@��414@�Gu��!?i�ܷE<�@�t����ٿ�ؿ�١�@��414@�Gu��!?i�ܷE<�@�����ٿ����X�@ۥ~G4@4V��ܐ!?؈aw�@�����ٿ����X�@ۥ~G4@4V��ܐ!?؈aw�@�����ٿ����X�@ۥ~G4@4V��ܐ!?؈aw�@�����ٿ����X�@ۥ~G4@4V��ܐ!?؈aw�@�����ٿ����X�@ۥ~G4@4V��ܐ!?؈aw�@�f;xɈٿЎ�e�m�@W��4@��Ɛ!?zI��@�f;xɈٿЎ�e�m�@W��4@��Ɛ!?zI��@����j�ٿq�F�{�@ȓ�a 4@z����!?̑�D�n�@����j�ٿq�F�{�@ȓ�a 4@z����!?̑�D�n�@����j�ٿq�F�{�@ȓ�a 4@z����!?̑�D�n�@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@�
��4�ٿ4��?A��@�N����3@3ˎ��!?��~����@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@8�#�ӆٿq���ќ�@�ݢ�64@J,D���!?4�?�7��@�p}��ٿ�\3����@�j��4@d��yҐ!?�D�J�|�@�p}��ٿ�\3����@�j��4@d��yҐ!?�D�J�|�@�p}��ٿ�\3����@�j��4@d��yҐ!?�D�J�|�@�p}��ٿ�\3����@�j��4@d��yҐ!?�D�J�|�@%+��Áٿ�3~5���@�"�S�	4@QUy�!?�����@�<C�ٿ�����H�@���G�4@�a�;��!?�s��:�@�<C�ٿ�����H�@���G�4@�a�;��!?�s��:�@�8ٿ\�Nk�M�@�8�w�4@�īt�!?�i�_�	�@�8ٿ\�Nk�M�@�8�w�4@�īt�!?�i�_�	�@�8ٿ\�Nk�M�@�8�w�4@�īt�!?�i�_�	�@�8ٿ\�Nk�M�@�8�w�4@�īt�!?�i�_�	�@�8ٿ\�Nk�M�@�8�w�4@�īt�!?�i�_�	�@i�gϋٿ�Gd��@���NQ4@*DG�S�!?1)H�t�@i�gϋٿ�Gd��@���NQ4@*DG�S�!?1)H�t�@i�gϋٿ�Gd��@���NQ4@*DG�S�!?1)H�t�@i�gϋٿ�Gd��@���NQ4@*DG�S�!?1)H�t�@i�gϋٿ�Gd��@���NQ4@*DG�S�!?1)H�t�@�5lC�ٿ�襟C��@ٙ���4@��,m�!?�׾!���@�5lC�ٿ�襟C��@ٙ���4@��,m�!?�׾!���@�5lC�ٿ�襟C��@ٙ���4@��,m�!?�׾!���@v��O��ٿ �|K_g�@�@[��4@}R����!?���qs�@v��O��ٿ �|K_g�@�@[��4@}R����!?���qs�@�4�)�ٿ%I��9��@+�s?4@����!?Hn�t�@M;�I�ٿ1�{ˣ��@�X�;~�3@�\j���!?�b�e&�@M;�I�ٿ1�{ˣ��@�X�;~�3@�\j���!?�b�e&�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@2/���ٿ�D^)
�@�~Υ��3@�����!?�jQ�NW�@���	�ٿl�6��@����94@P$j�+�!?�_C6B�@�I��ٿ[�(��@F��3%4@6{T���!?M_4�4��@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@݃����ٿ�&f��|�@,X[��4@�ѐ�!?��D�4%�@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@���j��ٿ4�b``�@���o�4@P�鶹�!?CJf+'��@�_��ٿ	��*���@K�!U4@��D�А!?���T��@��5���ٿ$��A��@��c��4@�}�+�!?S��s=0�@��5���ٿ$��A��@��c��4@�}�+�!?S��s=0�@��5���ٿ$��A��@��c��4@�}�+�!?S��s=0�@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�[ ��ٿ�͚�h�@4���4@zw�Hא!?+T�2��@�
ė]�ٿ3L@�[��@�Hg^�4@�{�Wɐ!?D���>}�@Ѭ��ٿ�������@��m��4@o4�u�!?��|���@Ѭ��ٿ�������@��m��4@o4�u�!?��|���@Ѭ��ٿ�������@��m��4@o4�u�!?��|���@Ѭ��ٿ�������@��m��4@o4�u�!?��|���@Ѭ��ٿ�������@��m��4@o4�u�!?��|���@[��u͏ٿ����6��@�Z�4@�"�ޥ�!?IbQ���@s8�~��ٿ@Y�g-�@�<���4@���uؐ!?B�g�/�@s8�~��ٿ@Y�g-�@�<���4@���uؐ!?B�g�/�@s8�~��ٿ@Y�g-�@�<���4@���uؐ!?B�g�/�@s8�~��ٿ@Y�g-�@�<���4@���uؐ!?B�g�/�@s8�~��ٿ@Y�g-�@�<���4@���uؐ!?B�g�/�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�,Y��ٿ�-݄��@����44@�ɉ/��!?i�B� X�@�UY�K�ٿ[�b��@5;S�4@ljZ��!?2>�����@a�Ӻ�ٿ�a�����@.?)��3@�DXc�!?I�����@a�Ӻ�ٿ�a�����@.?)��3@�DXc�!?I�����@a�Ӻ�ٿ�a�����@.?)��3@�DXc�!?I�����@a�Ӻ�ٿ�a�����@.?)��3@�DXc�!?I�����@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@���R��ٿR���y��@WG��y4@^&����!?�9_fQ�@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@��\8Յٿ���0�@�]���4@�@z��!?
*�h��@�jcL�ٿ��B"�@��8�4@EnkÚ�!?S׬����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����ˆٿ_G�w���@h���4@����!?�����@����K�ٿ��u���@����q4@�-����!?������@����K�ٿ��u���@����q4@�-����!?������@����K�ٿ��u���@����q4@�-����!?������@����K�ٿ��u���@����q4@�-����!?������@AX�&�~ٿξc*&�@ ��4@���֐!?*�Y�a'�@� ͮ�ٿK��R��@ ��_�3@sg��Ր!?^"�����@� ͮ�ٿK��R��@ ��_�3@sg��Ր!?^"�����@++,��ٿT�;|�!�@�kb-��3@�e�F�!?�/.F���@++,��ٿT�;|�!�@�kb-��3@�e�F�!?�/.F���@qe�ٿ�C|힧�@��V4@^��(�!?�N�(D�@qe�ٿ�C|힧�@��V4@^��(�!?�N�(D�@7�`H�ٿ�r�y0�@�j��4@�Ça�!??s&����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@#���r�ٿC�:7~x�@�Qo~4@������!?DS����@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@C8�+b�ٿ�r|��@.&pA|4@�m;�!?xԼ8v�@1v(��}ٿv݉`�@�9V~� 4@!����!?P�����@����ٿ��Jv��@=xY44@jE�(ǐ!?���tj�@����ٿ��Jv��@=xY44@jE�(ǐ!?���tj�@����ٿ��Jv��@=xY44@jE�(ǐ!?���tj�@����ٿ��Jv��@=xY44@jE�(ǐ!?���tj�@$��0,�ٿ�1�O^�@�34@P��!?+�si���@$��0,�ٿ�1�O^�@�34@P��!?+�si���@$��0,�ٿ�1�O^�@�34@P��!?+�si���@$��0,�ٿ�1�O^�@�34@P��!?+�si���@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@���!�ٿE�5*�@`�=�4@W�V�!?b兺i��@����ٿx��4�3�@=T>���3@w�_*�!?�ab �@����P�ٿ��k��c�@�c Z4@�Z��!?��Z�3�@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@O
;�ٿ�ݟ\m�@A�f=4@͠�C�!?�����@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@�.�s'�ٿTf��p��@y�8m84@q8���!?q�N	 ��@~��n��ٿ,B�TD[�@u �Kt4@�{�ː!?;�c�O��@~��n��ٿ,B�TD[�@u �Kt4@�{�ː!?;�c�O��@~��n��ٿ,B�TD[�@u �Kt4@�{�ː!?;�c�O��@�OM��ٿ���/��@Ii�R�4@�$���!?`�8��@����u�ٿ�8�i��@�f��4@sPO�}�!?���C6Y�@����u�ٿ�8�i��@�f��4@sPO�}�!?���C6Y�@K�&ݿ�ٿT��o��@����r4@���F��!?�����@K�&ݿ�ٿT��o��@����r4@���F��!?�����@K�&ݿ�ٿT��o��@����r4@���F��!?�����@K�&ݿ�ٿT��o��@����r4@���F��!?�����@7I$ҽ�ٿ���:�@���4@u�y���!?�p�t��@7I$ҽ�ٿ���:�@���4@u�y���!?�p�t��@7I$ҽ�ٿ���:�@���4@u�y���!?�p�t��@7I$ҽ�ٿ���:�@���4@u�y���!?�p�t��@�r	�߈ٿo�ԓD�@�P�!�4@�j�0��!?�V-�@�r	�߈ٿo�ԓD�@�P�!�4@�j�0��!?�V-�@�r	�߈ٿo�ԓD�@�P�!�4@�j�0��!?�V-�@3M���ٿ������@�ss�~4@�;�ؐ!?�+����@3M���ٿ������@�ss�~4@�;�ؐ!?�+����@3M���ٿ������@�ss�~4@�;�ؐ!?�+����@��f�]�ٿ��<t$��@^ZL4@��wh|�!?���I�@��f�]�ٿ��<t$��@^ZL4@��wh|�!?���I�@��f�]�ٿ��<t$��@^ZL4@��wh|�!?���I�@��f�]�ٿ��<t$��@^ZL4@��wh|�!?���I�@
�\�؂ٿ�A��=��@0�(G4@^�2��!?���|�@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�8�ٿ�_y�%��@�DhW�4@�A�d��!?�s�?��@�;�k�ٿs(�٣��@\�pE4@r�ڐ!?F[�ı�@�;�k�ٿs(�٣��@\�pE4@r�ڐ!?F[�ı�@d딢�ٿSV��P��@ ���4@�ӸS�!?SZ5D�E�@d딢�ٿSV��P��@ ���4@�ӸS�!?SZ5D�E�@d딢�ٿSV��P��@ ���4@�ӸS�!?SZ5D�E�@d딢�ٿSV��P��@ ���4@�ӸS�!?SZ5D�E�@d딢�ٿSV��P��@ ���4@�ӸS�!?SZ5D�E�@���H
�ٿն�'��@��?B�4@��	w��!?fLF�O��@���H
�ٿն�'��@��?B�4@��	w��!?fLF�O��@���H
�ٿն�'��@��?B�4@��	w��!?fLF�O��@���H
�ٿն�'��@��?B�4@��	w��!?fLF�O��@�%�	�ٿ[�����@�p`�T4@�����!?t����@�%�	�ٿ[�����@�p`�T4@�����!?t����@�%�	�ٿ[�����@�p`�T4@�����!?t����@�%�	�ٿ[�����@�p`�T4@�����!?t����@�yeՀ�ٿ݅�g���@8��gr4@���"��!?�J�@�yeՀ�ٿ݅�g���@8��gr4@���"��!?�J�@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@8dn�c�ٿv�wM��@��y��4@��˩e�!?`�U`B��@��3�ٿ�e��ߙ�@*]�N�4@Mh��d�!?C�V�u�@�V؂�ٿ���)�@�3���4@�=�"��!?a3���@�V؂�ٿ���)�@�3���4@�=�"��!?a3���@�V؂�ٿ���)�@�3���4@�=�"��!?a3���@�V؂�ٿ���)�@�3���4@�=�"��!?a3���@�V؂�ٿ���)�@�3���4@�=�"��!?a3���@3"�H�ٿ.����@�Mv��4@���0��!?���Cd��@3"�H�ٿ.����@�Mv��4@���0��!?���Cd��@��c�ٿa ���@��'�4@�1���!?&<�ӆ�@��c�ٿa ���@��'�4@�1���!?&<�ӆ�@�����ٿ�1�B��@}���4@K�/��!?\���1�@�����ٿ�1�B��@}���4@K�/��!?\���1�@�����ٿ�1�B��@}���4@K�/��!?\���1�@�����ٿ�1�B��@}���4@K�/��!?\���1�@�^r��ٿ�m�C��@��	�\ 4@}�*�ڐ!?)�x��@�^r��ٿ�m�C��@��	�\ 4@}�*�ڐ!?)�x��@*��#E�ٿ��h��)�@����4@>��u��!?�@%���@*��#E�ٿ��h��)�@����4@>��u��!?�@%���@*��#E�ٿ��h��)�@����4@>��u��!?�@%���@�ֽ�ٿ�E�r�@0�K4@T惝��!?21md��@ݾ>���ٿ?�����@{�։�4@L�q�!?蔆���@	{���ٿ-}8B��@���� 4@�+E}�!?����i��@	{���ٿ-}8B��@���� 4@�+E}�!?����i��@	{���ٿ-}8B��@���� 4@�+E}�!?����i��@=4S���ٿH"�A��@s3@^4@���!?��/��@=4S���ٿH"�A��@s3@^4@���!?��/��@f|�d��ٿ�N�����@9�l�4@|�_��!?w��Q���@0�~d�ٿ�������@�+O84@�*�V��!?(\s��@0�~d�ٿ�������@�+O84@�*�V��!?(\s��@0�~d�ٿ�������@�+O84@�*�V��!?(\s��@���?ǅٿ��G?0��@
�٭4@s�����!?�W%��r�@���?ǅٿ��G?0��@
�٭4@s�����!?�W%��r�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@������ٿ\��ѣ�@��d/4@�
��!?[�ce?�@y��`{ٿYSG5��@����g4@�鬙�!?�ؖ���@y��`{ٿYSG5��@����g4@�鬙�!?�ؖ���@y��`{ٿYSG5��@����g4@�鬙�!?�ؖ���@y��`{ٿYSG5��@����g4@�鬙�!?�ؖ���@y��`{ٿYSG5��@����g4@�鬙�!?�ؖ���@q���-}ٿ1�t���@��h�E 4@DK����!?�8�f��@5w0�*{ٿ�鴲�2�@�u���3@q��!?������@5w0�*{ٿ�鴲�2�@�u���3@q��!?������@5w0�*{ٿ�鴲�2�@�u���3@q��!?������@�ي�_�ٿu��~�{�@�6>�4@9w�K\�!?R��E��@�ي�_�ٿu��~�{�@�6>�4@9w�K\�!?R��E��@d5�}}ٿ�и�9�@�,��4@��PՁ�!?#qy�@}��v�ٿu����@TQ�]4@��-��!?1�0hl��@}��v�ٿu����@TQ�]4@��-��!?1�0hl��@l�y)�ٿ6t-��@$^�=4@,�X��!?���x�e�@{�̃ӇٿH�6w0�@8��h4@���^��!?�\\�S�@{�̃ӇٿH�6w0�@8��h4@���^��!?�\\�S�@{�̃ӇٿH�6w0�@8��h4@���^��!?�\\�S�@���K�ٿT�����@\���r4@WC-���!?..�����@���K�ٿT�����@\���r4@WC-���!?..�����@���K�ٿT�����@\���r4@WC-���!?..�����@���K�ٿT�����@\���r4@WC-���!?..�����@���K�ٿT�����@\���r4@WC-���!?..�����@���K�ٿT�����@\���r4@WC-���!?..�����@��J�;�ٿ��e���@E���4@k����!?�I��B�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@|���ٿ��-����@�86�E4@@?㚐!?�6��@�@��>�g�ٿܾ{���@'��5�4@]��!?�'�X�-�@�8��+�ٿQ�L���@�98hP4@�Z�А!?2h�t��@�8��+�ٿQ�L���@�98hP4@�Z�А!?2h�t��@�8��+�ٿQ�L���@�98hP4@�Z�А!?2h�t��@�4�@b�ٿ�%���#�@"��4@������!?[��95u�@�4�@b�ٿ�%���#�@"��4@������!?[��95u�@�4�@b�ٿ�%���#�@"��4@������!?[��95u�@�4�@b�ٿ�%���#�@"��4@������!?[��95u�@�4�@b�ٿ�%���#�@"��4@������!?[��95u�@wE|��ٿ�����l�@��\�4@w��~�!?���q1�@wE|��ٿ�����l�@��\�4@w��~�!?���q1�@zS����ٿ5��(�
�@
A74@:����!?�#�x���@zS����ٿ5��(�
�@
A74@:����!?�#�x���@��0ѷ�ٿ����m�@˅���4@}Q���!?@�kE��@��0ѷ�ٿ����m�@˅���4@}Q���!?@�kE��@��0ѷ�ٿ����m�@˅���4@}Q���!?@�kE��@e����ٿz�qe�@@"ʱ4@�$2�!?ܖ
TZ�@e����ٿz�qe�@@"ʱ4@�$2�!?ܖ
TZ�@e����ٿz�qe�@@"ʱ4@�$2�!?ܖ
TZ�@e����ٿz�qe�@@"ʱ4@�$2�!?ܖ
TZ�@e����ٿz�qe�@@"ʱ4@�$2�!?ܖ
TZ�@k$�<P�ٿ��^!��@a"�i�4@z����!?*�<џe�@k$�<P�ٿ��^!��@a"�i�4@z����!?*�<џe�@C�9�L�ٿ����2\�@�m��
4@�d�v�!?�~��N�@C�9�L�ٿ����2\�@�m��
4@�d�v�!?�~��N�@��I�l�ٿ��U�|�@�Yn4@ ��=��!?Zr��@r�����ٿ���K��@��e�4@�4B�!?5�}RM�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@ˋ��	�ٿ��<̝-�@c�m�4@k��!?R�]�գ�@f��³�ٿ���a��@�Ce4@i����!?dx��/�@E���'�ٿb9�Û�@&	:w4@$��{��!?�6���|�@E���'�ٿb9�Û�@&	:w4@$��{��!?�6���|�@E���'�ٿb9�Û�@&	:w4@$��{��!?�6���|�@E���'�ٿb9�Û�@&	:w4@$��{��!?�6���|�@���-�ٿ*��Z��@܇���4@����!?������@���-�ٿ*��Z��@܇���4@����!?������@Ac�tG�ٿ^�����@�	��4@�>�ݐ!?�Wl����@Ac�tG�ٿ^�����@�	��4@�>�ݐ!?�Wl����@ �_J$�ٿ~�>D���@/�w4@@=ڐ!?[^�j��@.��%�ٿ}���.�@�H�p 4@�/5�!?�P��`q�@.��%�ٿ}���.�@�H�p 4@�/5�!?�P��`q�@�+7�ٿ�i,�@���4@`�Yj��!?S�Oط��@�+7�ٿ�i,�@���4@`�Yj��!?S�Oط��@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��!H�ٿ����@��P��3@8�U�Ԑ!?	���M�@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@��Z��ٿ	vgp~N�@��F�q�3@R��aԐ!?_�����@�bc��ٿ����S��@D�۶W 4@:���ѐ!?�4�c	��@SB�5k�ٿ��k���@��3�4@!��Tؐ!?5�IZe`�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@tWԌ|�ٿ�Hy#��@��X�4@D��+��!?}�h uI�@E  ��ٿ�� �@s�@���4@����!?Esj�<��@E  ��ٿ�� �@s�@���4@����!?Esj�<��@E  ��ٿ�� �@s�@���4@����!?Esj�<��@E  ��ٿ�� �@s�@���4@����!?Esj�<��@E  ��ٿ�� �@s�@���4@����!?Esj�<��@���ˍٿ*k��rp�@�s��4@����!?�*�G�o�@A�!��ٿ�{:y��@돁�"4@���!?�
Zn�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@q���ٿ@Q"��@W�1�4@�#��!?�����M�@���Zߌٿ��;��@�m�&4@�/5帐!?@5�� ��@���Zߌٿ��;��@�m�&4@�/5帐!?@5�� ��@v��긅ٿyV{X�C�@Gi�m�4@��@��!?nCb�@v��긅ٿyV{X�C�@Gi�m�4@��@��!?nCb�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@7q�-�ٿq��LW�@u4�e�4@��7#��!?;#�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ձ��C�ٿ������@Tj�ֵ4@ʨ?j��!?���Uv�@ H��ٿsB��@i�� 4@}����!?��[]W�@ H��ٿsB��@i�� 4@}����!?��[]W�@ H��ٿsB��@i�� 4@}����!?��[]W�@ H��ٿsB��@i�� 4@}����!?��[]W�@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@�S��ٿ�h��6 �@Z���v4@��p���!?����@��9Ɩ�ٿھR��@2�sz�4@�$��А!?a�4�"�@��9Ɩ�ٿھR��@2�sz�4@�$��А!?a�4�"�@��9Ɩ�ٿھR��@2�sz�4@�$��А!?a�4�"�@��9Ɩ�ٿھR��@2�sz�4@�$��А!?a�4�"�@��9Ɩ�ٿھR��@2�sz�4@�$��А!?a�4�"�@���T��ٿ��v����@7x*K�4@X��!?��f&U��@�u۟��ٿ��` ��@{ @Μ4@-�>ڐ�!?�+�@�u۟��ٿ��` ��@{ @Μ4@-�>ڐ�!?�+�@ߴ����ٿ���;&�@&���� 4@	�"��!?���'��@ߴ����ٿ���;&�@&���� 4@	�"��!?���'��@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@.BkcE�ٿ���1l��@,�B]\ 4@��@ƀ�!?5
uN���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@x��!:vٿYú�?��@�ԱM4@��/��!?�%P#���@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@볊ȅٿ�Q����@�ݘ�Z4@�~| Ȑ!?�F��XG�@a�q�ٿ�]�N"��@��244@{�`Ő!?>�G���@a�q�ٿ�]�N"��@��244@{�`Ő!?>�G���@a�q�ٿ�]�N"��@��244@{�`Ő!?>�G���@����ٿ�K����@�nM��4@0�����!?Q�2F��@����ٿ�K����@�nM��4@0�����!?Q�2F��@����ٿ�K����@�nM��4@0�����!?Q�2F��@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@>�l���ٿ��F��#�@3�7�4@�GH��!?����@�Ͱ�ٿ?�W����@����4@sm�T�!?�?�-�Y�@�A@��ٿK�V��h�@	sJ�4@[{�$��!?�
�2�[�@�A@��ٿK�V��h�@	sJ�4@[{�$��!?�
�2�[�@�A@��ٿK�V��h�@	sJ�4@[{�$��!?�
�2�[�@�A@��ٿK�V��h�@	sJ�4@[{�$��!?�
�2�[�@�A@��ٿK�V��h�@	sJ�4@[{�$��!?�
�2�[�@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@�䅽��ٿ�!�E�E�@��41T 4@Afr�!?R��4��@+4��Q�ٿ��!��@:�AYP 4@�����!?	o����@+4��Q�ٿ��!��@:�AYP 4@�����!?	o����@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�N�R�ٿ�<g��@.Qq}� 4@�剐!?�؂ϋ��@�!���ٿt�H�3|�@nFv��4@���Ő!?_���;�@�!���ٿt�H�3|�@nFv��4@���Ő!?_���;�@�!���ٿt�H�3|�@nFv��4@���Ő!?_���;�@}�'/�ٿ6�z�	�@�� 4@Z�����!?m���6h�@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@/;-��ٿ6a�q�@�"�<Y4@�G�Ȑ!?C�� ���@p����ٿ>T\Ƕ�@��j4@dm`7��!?و�����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@�C�*�ٿDY�8���@mM�4@��%̐!?��}����@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@����:�ٿo�J��@��k��4@��^�ِ!?d �t���@��B��ٿV����u�@d*�4@5��ߐ!?�u�I��@��B��ٿV����u�@d*�4@5��ߐ!?�u�I��@��B��ٿV����u�@d*�4@5��ߐ!?�u�I��@��Iݨ�ٿ�5�����@�}V�4@����!?1�v$��@�����ٿ�����1�@�k��4@4 ����!?����z�@�����ٿ�����1�@�k��4@4 ����!?����z�@�����ٿ�����1�@�k��4@4 ����!?����z�@�lU��ٿ:n!wZ�@��q��4@qH�5��!?{2�e��@�lU��ٿ:n!wZ�@��q��4@qH�5��!?{2�e��@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@a��W��ٿޑ��9�@�~F�	4@$��)�!?kƚI3O�@I۔Äٿܑ�����@�|g�	4@)K��!?�����@I۔Äٿܑ�����@�|g�	4@)K��!?�����@I۔Äٿܑ�����@�|g�	4@)K��!?�����@� ���ٿ��YC��@j��_�	4@ٙ}ߐ!?@�c�S�@��?s�ٿ������@���.�4@�m�ߐ!?�AB�e��@��?s�ٿ������@���.�4@�m�ߐ!?�AB�e��@��?s�ٿ������@���.�4@�m�ߐ!?�AB�e��@��?s�ٿ������@���.�4@�m�ߐ!?�AB�e��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@SN (�ٿǔm|�
�@ܴ�"�4@AQ�+��!?�żߔ��@�S�P��ٿ0��[���@�ʃS4@���	�!?�pJ �@�S�P��ٿ0��[���@�ʃS4@���	�!?�pJ �@�S�P��ٿ0��[���@�ʃS4@���	�!?�pJ �@�S�P��ٿ0��[���@�ʃS4@���	�!?�pJ �@@ΐ��}ٿ7Ԋ���@����4@��$�!?L ,>I�@@ΐ��}ٿ7Ԋ���@����4@��$�!?L ,>I�@ 4��/}ٿ^�{&�B�@���4@+� �$�!?�𽼴��@&H��O|ٿ�e>��@�t*4�4@�����!?פ���@&H��O|ٿ�e>��@�t*4�4@�����!?פ���@&H��O|ٿ�e>��@�t*4�4@�����!?פ���@&H��O|ٿ�e>��@�t*4�4@�����!?פ���@&K0q�ٿ�4k���@Z�cĢ4@}@RY�!?+uJF�_�@&K0q�ٿ�4k���@Z�cĢ4@}@RY�!?+uJF�_�@&K0q�ٿ�4k���@Z�cĢ4@}@RY�!?+uJF�_�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@Z���K�ٿ�)��@,ڄ�04@&X�E��!?(+�]�!�@|�1߹�ٿ8��w��@ZT1��4@��;㪐!?R��y?��@|�1߹�ٿ8��w��@ZT1��4@��;㪐!?R��y?��@|�1߹�ٿ8��w��@ZT1��4@��;㪐!?R��y?��@|�1߹�ٿ8��w��@ZT1��4@��;㪐!?R��y?��@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@�ؖ�Ɂٿ�A�L���@1+5g4@��f��!?p�$��u�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@w&A]��ٿ������@�{4@��|�̐!?��!`�'�@��P���ٿ���4���@r�C���3@w��L��!?|��?�P�@��P���ٿ���4���@r�C���3@w��L��!?|��?�P�@/Sf7{ٿ�˒{�s�@���V 4@FE[א!?3T%F�I�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@C�rˀٿQ c��@�,v*4@����!?��7 um�@����
�ٿ���|ص�@V��o4@D�`���!?���,��@u���`�ٿ9�w���@�Wuw4@v7�ɐ!?��JҊ8�@u���`�ٿ9�w���@�Wuw4@v7�ɐ!?��JҊ8�@u���`�ٿ9�w���@�Wuw4@v7�ɐ!?��JҊ8�@u���`�ٿ9�w���@�Wuw4@v7�ɐ!?��JҊ8�@�2���ٿ�N� :�@i*�ln4@�G����!?0�LM�@�2���ٿ�N� :�@i*�ln4@�G����!?0�LM�@�2���ٿ�N� :�@i*�ln4@�G����!?0�LM�@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@��$���ٿ�l��(X�@u��84@xn��!?�*�%
��@F_��E�ٿ�kE5~��@���Z4@	�fqސ!?�ܲċH�@F_��E�ٿ�kE5~��@���Z4@	�fqސ!?�ܲċH�@F_��E�ٿ�kE5~��@���Z4@	�fqސ!?�ܲċH�@F_��E�ٿ�kE5~��@���Z4@	�fqސ!?�ܲċH�@F_��E�ٿ�kE5~��@���Z4@	�fqސ!?�ܲċH�@p6����ٿ�A�iY�@J'��4@B��4��!?���8�7�@�i�[��ٿ{Dh���@J�b��4@����!?:�gj�4�@�i�[��ٿ{Dh���@J�b��4@����!?:�gj�4�@�i�[��ٿ{Dh���@J�b��4@����!?:�gj�4�@�w;�~ٿI$=����@��7�z4@���	�!?H$��@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@kҜ�ٿ���
��@*��^4@&���!?vj[�4]�@a��ZL�ٿ;���j��@+����4@�W����!?@1�KHp�@a��ZL�ٿ;���j��@+����4@�W����!?@1�KHp�@a��ZL�ٿ;���j��@+����4@�W����!?@1�KHp�@a��ZL�ٿ;���j��@+����4@�W����!?@1�KHp�@a��ZL�ٿ;���j��@+����4@�W����!?@1�KHp�@Ï�n�ٿ�����@B�~4@ȁ!\e�!?��ݬ�@Ï�n�ٿ�����@B�~4@ȁ!\e�!?��ݬ�@�Z:��ٿ�(Z���@`�/e�4@�»�T�!?�v�YM�@�Z:��ٿ�(Z���@`�/e�4@�»�T�!?�v�YM�@�Z:��ٿ�(Z���@`�/e�4@�»�T�!?�v�YM�@�%�g�ٿ@�b��@#�@	4@�D�hy�!?Ð����@�%�g�ٿ@�b��@#�@	4@�D�hy�!?Ð����@d{�|ٿ���B��@�keP4@���5ې!?@�JH�@!�i�P�ٿ�3/���@�^e�4@���8�!?����Z�@!�i�P�ٿ�3/���@�^e�4@���8�!?����Z�@!�i�P�ٿ�3/���@�^e�4@���8�!?����Z�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@�z����ٿ�f���@9���+�3@0��u,�!?���P�p�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@9u� �ٿ���@��r4@3��!?;���w.�@��i�h�ٿ0w#���@�.k>~4@�)T�!?�:�,V�@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@_�,�ˇٿef��^�@v|�4@#�l�0�!?#�z��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@3'ҳ�ٿ���BO�@� U�4@����Ȑ!?�20��@�>7~ٿ��?�
�@���<$4@�BA��!?�}�
�-�@>O�z�ٿ!�R���@��l�4@�iL�D�!?'�ON��@#����ٿ2�C���@efM$4@��n��!?�*�"��@Sd�+�~ٿ�)1�m��@��w4@�.��ސ!?!z=1���@Sd�+�~ٿ�)1�m��@��w4@�.��ސ!?!z=1���@Sd�+�~ٿ�)1�m��@��w4@�.��ސ!?!z=1���@T�V b�ٿ��z���@eh�^T4@9r��!?HY��K��@T�V b�ٿ��z���@eh�^T4@9r��!?HY��K��@T�V b�ٿ��z���@eh�^T4@9r��!?HY��K��@ey_(C�ٿ�r7x� �@���(�4@Cf����!?1=ʔ/�@+�y=W�ٿ�iY���@��Df*4@�6/�!?�y#��@+�y=W�ٿ�iY���@��Df*4@�6/�!?�y#��@c��v^�ٿ6�s�i�@<o�\4@�T���!? X�k�@%����|ٿ^���y�@�o��c	4@)vo�Ɛ!?`��WǸ�@%����|ٿ^���y�@�o��c	4@)vo�Ɛ!?`��WǸ�@�b�8E�ٿ������@oE��4@U����!?K-�4d�@�b�8E�ٿ������@oE��4@U����!?K-�4d�@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�P 2�ٿ���;��@1��v4@U#M�!?e��P	��@�����ٿ��ϸm�@�R���4@���D�!?@����@�����ٿ��ϸm�@�R���4@���D�!?@����@��t�
zٿ���m�@���4@��2��!?������@��t�
zٿ���m�@���4@��2��!?������@��t�
zٿ���m�@���4@��2��!?������@��t�
zٿ���m�@���4@��2��!?������@��t�
zٿ���m�@���4@��2��!?������@�>힎yٿ�H����@�c<4@-�=}�!?�$�3��@�>힎yٿ�H����@�c<4@-�=}�!?�$�3��@�>힎yٿ�H����@�c<4@-�=}�!?�$�3��@Ʈ�Mzٿ��pS�(�@zq*4@�T5_�!?;�0���@Ʈ�Mzٿ��pS�(�@zq*4@�T5_�!?;�0���@Ʈ�Mzٿ��pS�(�@zq*4@�T5_�!?;�0���@��v�zٿ���J�[�@�Y"F4@M�Q(��!?͙J���@��v�zٿ���J�[�@�Y"F4@M�Q(��!?͙J���@��v�zٿ���J�[�@�Y"F4@M�Q(��!?͙J���@��v�zٿ���J�[�@�Y"F4@M�Q(��!?͙J���@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@��53Ƈٿ�_H�]�@��/���3@Ɂ鷍�!?R��W�@�7����ٿ�j�����@��	��3@kE�rl�!?��
�9�@R�z�~ٿ�Cށ��@J$�4@�ʰ%ǐ!?�k����@R�z�~ٿ�Cށ��@J$�4@�ʰ%ǐ!?�k����@R�z�~ٿ�Cށ��@J$�4@�ʰ%ǐ!?�k����@R�z�~ٿ�Cށ��@J$�4@�ʰ%ǐ!?�k����@R�z�~ٿ�Cށ��@J$�4@�ʰ%ǐ!?�k����@�h����ٿ�H�4���@�~�$ 4@_JRo�!?�����@�Ëi�ٿ�@K'6g�@�����4@�c-^�!?o�'�ދ�@�Ëi�ٿ�@K'6g�@�����4@�c-^�!?o�'�ދ�@�Ëi�ٿ�@K'6g�@�����4@�c-^�!?o�'�ދ�@�Ëi�ٿ�@K'6g�@�����4@�c-^�!?o�'�ދ�@�Ëi�ٿ�@K'6g�@�����4@�c-^�!?o�'�ދ�@,��ٿ��4Q
�@��H 4@��9k�!?�#ԗ�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@$Y����ٿ"�����@����84@�c¡��!?���9�@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@IF�ɺ�ٿ�w�U�l�@~��74@��vh�!?s������@<��?�ٿ< :}��@r����4@���ל�!?*��8�@��]���ٿ|x�"(��@N�Ik�	4@Vj���!?������@e0�ٿ�,=�@/���54@T��|�!?5����@V0��ٿw"h���@^���n4@B����!?�Y�.$6�@V0��ٿw"h���@^���n4@B����!?�Y�.$6�@V0��ٿw"h���@^���n4@B����!?�Y�.$6�@V0��ٿw"h���@^���n4@B����!?�Y�.$6�@� @2�ٿ����z�@
zKz�4@MUm�!?j�b�^��@� @2�ٿ����z�@
zKz�4@MUm�!?j�b�^��@��hZ�ٿ����A�@�z;;�4@c�FPH�!?�[�t,&�@��hZ�ٿ����A�@�z;;�4@c�FPH�!?�[�t,&�@��hZ�ٿ����A�@�z;;�4@c�FPH�!?�[�t,&�@��hZ�ٿ����A�@�z;;�4@c�FPH�!?�[�t,&�@��hZ�ٿ����A�@�z;;�4@c�FPH�!?�[�t,&�@Cz���ٿ���B�'�@���!~	4@�{��!?���G�@Cz���ٿ���B�'�@���!~	4@�{��!?���G�@Cz���ٿ���B�'�@���!~	4@�{��!?���G�@Cz���ٿ���B�'�@���!~	4@�{��!?���G�@����ٿ�7��{K�@�<C4@�!$ڐ!?&90$`�@����ٿ�7��{K�@�<C4@�!$ڐ!?&90$`�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@�GmZ��ٿ��TOS�@���|4@CJ��А!?�9�h%/�@@Aؒٿ6v�,���@}�ף�4@�����!?h�89�@@Aؒٿ6v�,���@}�ף�4@�����!?h�89�@@Aؒٿ6v�,���@}�ף�4@�����!?h�89�@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@�`Q)�ٿ�{>Y��@�yUt4@�#�9!?5���]��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@���.�ٿX��R ��@�1���4@"�Nn�!?���K��@"%��ٿG�����@6%4��4@q��͐!?�9島�@"%��ٿG�����@6%4��4@q��͐!?�9島�@"%��ٿG�����@6%4��4@q��͐!?�9島�@"%��ٿG�����@6%4��4@q��͐!?�9島�@"%��ٿG�����@6%4��4@q��͐!?�9島�@^�"��ٿ�ts��@�H�i4@�꙾��!?=�O����@^�"��ٿ�ts��@�H�i4@�꙾��!?=�O����@^�"��ٿ�ts��@�H�i4@�꙾��!?=�O����@^�"��ٿ�ts��@�H�i4@�꙾��!?=�O����@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@齻���ٿ�np���@J�G>/4@�u����!?���y�A�@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@
����ٿ�H^[���@�M)<4@3rِ֧!? E����@U*���ٿ�q����@��[�4@W�犐!? �}W�@l���ٿk�n��@i�аu4@#鍕�!?a�A;{~�@l���ٿk�n��@i�аu4@#鍕�!?a�A;{~�@l���ٿk�n��@i�аu4@#鍕�!?a�A;{~�@��+���ٿh�*I�v�@|m_�4@�Yjw��!?�~�"��@��+���ٿh�*I�v�@|m_�4@�Yjw��!?�~�"��@��+���ٿh�*I�v�@|m_�4@�Yjw��!?�~�"��@�Zh���ٿZ�tP+��@���4@����א!?�P�>�@�@�Zh���ٿZ�tP+��@���4@����א!?�P�>�@�@�Zh���ٿZ�tP+��@���4@����א!?�P�>�@�@�Zh���ٿZ�tP+��@���4@����א!?�P�>�@�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@�	4�E{ٿ�.�e���@�B�4@ܗ5-��!?�U�@O33�ٿ�F�Cs�@����14@'Z-���!?��h���@O33�ٿ�F�Cs�@����14@'Z-���!?��h���@O33�ٿ�F�Cs�@����14@'Z-���!?��h���@O33�ٿ�F�Cs�@����14@'Z-���!?��h���@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�x��ٿ� ����@e�\�4@�z�2�!?xn�i��@�3�I�ٿҩӠ��@����4@]8��A�!?�fc��@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@�W]�q�ٿ�hd~[��@�0�{4@���K�!?U^6���@1U-��ٿ�9֙���@��;���3@s�9l��!?$7,�!N�@1U-��ٿ�9֙���@��;���3@s�9l��!?$7,�!N�@�r�ǋٿ o����@]i��4@�\E�!?���x���@�r�ǋٿ o����@]i��4@�\E�!?���x���@�r�ǋٿ o����@]i��4@�\E�!?���x���@�r�ǋٿ o����@]i��4@�\E�!?���x���@ڗRNk�ٿ*N}�Y�@dǡ!4@Y�q��!?j$=l26�@��8�ٿ�n'e���@��^U=4@θ���!?E0��@��8�ٿ�n'e���@��^U=4@θ���!?E0��@h��=Տٿu�oca��@e��4@A[�Bb�!?8��e��@h��=Տٿu�oca��@e��4@A[�Bb�!?8��e��@�.0���ٿ��~7ƭ�@7�}� 4@0/p��!?>ʉ~�F�@�.0���ٿ��~7ƭ�@7�}� 4@0/p��!?>ʉ~�F�@�.0���ٿ��~7ƭ�@7�}� 4@0/p��!?>ʉ~�F�@�.0���ٿ��~7ƭ�@7�}� 4@0/p��!?>ʉ~�F�@�.0���ٿ��~7ƭ�@7�}� 4@0/p��!?>ʉ~�F�@�8"�>�ٿ������@�*�Ɣ4@�V∟�!?G�u�?�@�8"�>�ٿ������@�*�Ɣ4@�V∟�!?G�u�?�@�8"�>�ٿ������@�*�Ɣ4@�V∟�!?G�u�?�@X��a�ٿ����@�{��4@<���!?x�͎��@X��a�ٿ����@�{��4@<���!?x�͎��@C�*E�ٿ�}-�s?�@���ڂ4@m��;�!?��'����@C�*E�ٿ�}-�s?�@���ڂ4@m��;�!?��'����@C�*E�ٿ�}-�s?�@���ڂ4@m��;�!?��'����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@C����ٿZA��O��@��ȗK4@��,��!?;^����@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@7=`~�ٿ��Y;��@�"�+4@<;����!?����_�@ LJ�1�ٿ��h_�'�@&��4@�+��y�!?����@ LJ�1�ٿ��h_�'�@&��4@�+��y�!?����@ LJ�1�ٿ��h_�'�@&��4@�+��y�!?����@�[˄�ٿ��x4�@�^F�4@1�%�s�!?�0��@�[˄�ٿ��x4�@�^F�4@1�%�s�!?�0��@�[˄�ٿ��x4�@�^F�4@1�%�s�!?�0��@�[˄�ٿ��x4�@�^F�4@1�%�s�!?�0��@�����ٿ��\����@��ǀ�4@\�{i�!?)�f���@�����ٿ��\����@��ǀ�4@\�{i�!?)�f���@	s�lS�ٿR�̓u��@�^>8b4@�qא!?�rv3*��@	s�lS�ٿR�̓u��@�^>8b4@�qא!?�rv3*��@�\�lw�ٿa�셄�@�����4@cp%��!?䰑����@�\�lw�ٿa�셄�@�����4@cp%��!?䰑����@�`'#ٿ6;��X��@��cK�4@�'>�!?� |if��@�`'#ٿ6;��X��@��cK�4@�'>�!?� |if��@�`'#ٿ6;��X��@��cK�4@�'>�!?� |if��@�`'#ٿ6;��X��@��cK�4@�'>�!?� |if��@�ܟ-�ٿ�M�����@8��x�4@&��k�!?n� ٺ�@�ܟ-�ٿ�M�����@8��x�4@&��k�!?n� ٺ�@�Q�?s�ٿMH��L��@� d�4@"3�Wf�!?qW���@�Q�?s�ٿMH��L��@� d�4@"3�Wf�!?qW���@�Q�?s�ٿMH��L��@� d�4@"3�Wf�!?qW���@��D�ٿ7��嬘�@�1��;4@`ҵ;d�!?4�Q����@��D�ٿ7��嬘�@�1��;4@`ҵ;d�!?4�Q����@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@8g�]�ٿ���q<��@�vD�4@S1;�~�!?���;i]�@��a�K�ٿ�2�ߥi�@�6�^4@.���!?Kwr�&��@I��څٿk(�mJ}�@\]?�4@��Գ�!?�6**��@I��څٿk(�mJ}�@\]?�4@��Գ�!?�6**��@I��څٿk(�mJ}�@\]?�4@��Գ�!?�6**��@I��څٿk(�mJ}�@\]?�4@��Գ�!?�6**��@I��څٿk(�mJ}�@\]?�4@��Գ�!?�6**��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@�>�~s�ٿh�8/�=�@qM�74@����!?�GQ�2��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@w�c7��ٿ��Z�\�@�+<] 4@���=��!?�4�B@��@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@[>����ٿȤi���@i6&�! 4@I�Qn�!?�5�(�{�@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@]><���ٿ�8����@�� 7�4@�k��!?B�\jF��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@j�8�ٿ ���P�@�}C�	4@��N2��!?��G��@����ٿ���`ӊ�@�����4@�����!?Ц�����@����ٿ���`ӊ�@�����4@�����!?Ц�����@����ٿ���`ӊ�@�����4@�����!?Ц�����@����ٿ���`ӊ�@�����4@�����!?Ц�����@����ٿ���`ӊ�@�����4@�����!?Ц�����@����ٿiɉ� �@Ѻz�4@�r8�5�!?���l�@1�n:�ٿN:�	���@R�r>�4@���a4�!?����Xg�@1�n:�ٿN:�	���@R�r>�4@���a4�!?����Xg�@�PB&rٿ#�-�0��@���}4@'%d9�!?�J�����@b���ٿ��O��\�@���4@�H<�!?���A��@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@��O|�ٿ�`Y}���@�����4@*�@�ǐ!?��_�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@_
eS��ٿ�*E�Z��@����4@0�<沐!?@6̰�u�@�'�裋ٿv���=�@G�ԝ?4@��FI��!?4�f9�c�@�'�裋ٿv���=�@G�ԝ?4@��FI��!?4�f9�c�@�'�裋ٿv���=�@G�ԝ?4@��FI��!?4�f9�c�@�'�裋ٿv���=�@G�ԝ?4@��FI��!?4�f9�c�@˭Mb��ٿo��'���@؍�4@���p|�!?r/���t�@����B�ٿ�o�O�P�@���4@af��ɐ!?��ڋp�@"���ٿ�	O�@�.FzZ4@�����!?������@"���ٿ�	O�@�.FzZ4@�����!?������@"���ٿ�	O�@�.FzZ4@�����!?������@"���ٿ�	O�@�.FzZ4@�����!?������@"���ٿ�	O�@�.FzZ4@�����!?������@"���ٿ�	O�@�.FzZ4@�����!?������@4ڸeS�ٿ�y3�TW�@���� 4@{�Gg5�!?�@�%��@4ڸeS�ٿ�y3�TW�@���� 4@{�Gg5�!?�@�%��@6��"�zٿv�]����@��<4@}�>���!?��b�I�@����~ٿcR��+��@��d3�4@5���!?/�3P��@����~ٿcR��+��@��d3�4@5���!?/�3P��@7�l;�ٿ�q�/���@f
 �=4@�\u��!?y'�wE��@7�l;�ٿ�q�/���@f
 �=4@�\u��!?y'�wE��@u�m'�ٿJ�'un�@_g�z24@� ����!?s?0�u�@u�m'�ٿJ�'un�@_g�z24@� ����!?s?0�u�@u�m'�ٿJ�'un�@_g�z24@� ����!?s?0�u�@u�m'�ٿJ�'un�@_g�z24@� ����!?s?0�u�@abF�{ٿ=�L!z�@4D4@��DHV�!?�V� �$�@abF�{ٿ=�L!z�@4D4@��DHV�!?�V� �$�@abF�{ٿ=�L!z�@4D4@��DHV�!?�V� �$�@abF�{ٿ=�L!z�@4D4@��DHV�!?�V� �$�@abF�{ٿ=�L!z�@4D4@��DHV�!?�V� �$�@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@���Ѡ{ٿ�=oT���@o`�4@���א!?��N��@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@j�&��ٿ�pPK���@i%o�4@�2d���!?�V�X2s�@B�fL�ٿ��9�ح�@f?���4@DLH�א!?��@���@B�fL�ٿ��9�ح�@f?���4@DLH�א!?��@���@B�fL�ٿ��9�ح�@f?���4@DLH�א!?��@���@B�fL�ٿ��9�ح�@f?���4@DLH�א!?��@���@B�fL�ٿ��9�ح�@f?���4@DLH�א!?��@���@-:،ٿ��;��S�@k��X4@/��Q��!?�-!�߼�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@��J`�ٿ�D���@���`4@�-���!?�lP�V�@�d&\�ٿ�>��^�@���ކ4@�2��!?8�O`�@�d&\�ٿ�>��^�@���ކ4@�2��!?8�O`�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@(�*�Y�ٿ%��m�@�P}��4@��k6��!?*�W��(�@����ٿ��F��:�@#�ԕ<4@a$fא!?�7]J@'�@����ٿ��F��:�@#�ԕ<4@a$fא!?�7]J@'�@����ٿ��F��:�@#�ԕ<4@a$fא!?�7]J@'�@����ٿ��F��:�@#�ԕ<4@a$fא!?�7]J@'�@����ٿ��F��:�@#�ԕ<4@a$fא!?�7]J@'�@���~�ٿ� �x�@��~�4@�4��!?`����Q�@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@[ ��ٿ
�Z6���@є=b�4@�[�;ϐ!?�R1���@F�̶f�ٿn��<1b�@�{��4@
���!?��=����@F�̶f�ٿn��<1b�@�{��4@
���!?��=����@F�̶f�ٿn��<1b�@�{��4@
���!?��=����@F�̶f�ٿn��<1b�@�{��4@
���!?��=����@B��ٿp�J%`�@��s�4@jT0䔐!?ST475��@B��ٿp�J%`�@��s�4@jT0䔐!?ST475��@B��ٿp�J%`�@��s�4@jT0䔐!?ST475��@2��~ٿ���:���@�E$�4@�9aP�!?�� �-�@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@V���ٿy��M0��@�n�4@�;�]g�!?���-?��@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@��I`�ٿH��3��@5��2�4@�YEې!?��/�/|�@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@v���F�ٿ����r�@MX4@������!? �g����@��7��~ٿ�>q����@�N"�/4@�gE��!?A���V��@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@���Ńٿ��X�Y��@<Nb]4@ ��Dd�!?��E>�v�@
.���ٿs�)(��@=�܂�4@�f�.��!??	�f��@
.���ٿs�)(��@=�܂�4@�f�.��!??	�f��@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@�L�x��ٿ/٨8-��@�%� 4@�u �!?T% �1�@��@�l�ٿ�n�����@�p�\�4@'�z�!?�����@��@�l�ٿ�n�����@�p�\�4@'�z�!?�����@��@�l�ٿ�n�����@�p�\�4@'�z�!?�����@�ַ���ٿC	�d+��@�H���4@ ��3ߐ!?�,H|��@5�M^�ٿ�G�4[�@��4@�|�I͐!?W8_�wR�@5�M^�ٿ�G�4[�@��4@�|�I͐!?W8_�wR�@8�˨?�ٿxk�����@��\A�4@��-�!?�3y����@�Zڂٿ��e�	��@pYI��4@C��,N�!?%TR��@�Zڂٿ��e�	��@pYI��4@C��,N�!?%TR��@�Zڂٿ��e�	��@pYI��4@C��,N�!?%TR��@�Zڂٿ��e�	��@pYI��4@C��,N�!?%TR��@k����ٿ�: D��@��4@�_��)�!?��E~��@6,9,�ٿL����Z�@U�ݏ�4@,��!?I�pL�@6,9,�ٿL����Z�@U�ݏ�4@,��!?I�pL�@ �S��ٿD�����@��14@�(�!?$��x�X�@ �S��ٿD�����@��14@�(�!?$��x�X�@ �S��ٿD�����@��14@�(�!?$��x�X�@,H�ﶈٿb�d���@����,4@����!?$�4��@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@��� ��ٿ�p����@a��4@+c����!?�I�Q�@�(�[�ٿÏ���@t��|(4@/�O��!?2t����@�(�[�ٿÏ���@t��|(4@/�O��!?2t����@�(�[�ٿÏ���@t��|(4@/�O��!?2t����@�(�[�ٿÏ���@t��|(4@/�O��!?2t����@�(�[�ٿÏ���@t��|(4@/�O��!?2t����@�7%���ٿ����,�@z��֩4@�1ڐ!?��� ��@�7%���ٿ����,�@z��֩4@�1ڐ!?��� ��@�7%���ٿ����,�@z��֩4@�1ڐ!?��� ��@�7%���ٿ����,�@z��֩4@�1ڐ!?��� ��@^�j���ٿ) 	�.��@�Xf��4@��	��!? ��Tp�@^�j���ٿ) 	�.��@�Xf��4@��	��!? ��Tp�@^�j���ٿ) 	�.��@�Xf��4@��	��!? ��Tp�@^�j���ٿ) 	�.��@�Xf��4@��	��!? ��Tp�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@  ]�.�ٿ&.�/���@�]�"%4@vz�2ݐ!?�VB�&�@���ٿ��>����@"�gz�4@���ڐ!?�q(��@���ٿ��>����@"�gz�4@���ڐ!?�q(��@���ٿ��>����@"�gz�4@���ڐ!?�q(��@���ٿ��>����@"�gz�4@���ڐ!?�q(��@G,4�ٿE1��[��@!\+��4@�����!?d�;Uib�@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@om��4�ٿz�=״��@�%�N�4@�{��i�!?L�����@��*�#�ٿ6�S���@�Js��4@5�u��!?�4��
��@��*�#�ٿ6�S���@�Js��4@5�u��!?�4��
��@��*�#�ٿ6�S���@�Js��4@5�u��!?�4��
��@��*�#�ٿ6�S���@�Js��4@5�u��!?�4��
��@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@b��ٿ[��	߃�@@�Ta4@)G+^��!?��uk�@Y�.Φ�ٿ�	�Lx��@��!L4@��N���!?�h����@�T��ώٿƇ���@k�Ua�4@�O�Sk�!?�TBec��@�T��ώٿƇ���@k�Ua�4@�O�Sk�!?�TBec��@�T��ώٿƇ���@k�Ua�4@�O�Sk�!?�TBec��@r��_y�ٿ�5|Ȃ��@��B�j	4@��o�Ő!?eA��!�@r��_y�ٿ�5|Ȃ��@��B�j	4@��o�Ő!?eA��!�@r��_y�ٿ�5|Ȃ��@��B�j	4@��o�Ő!?eA��!�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@�n�ٿ��a����@Ԇa�� 4@����!?p�穫�@|N�)}ٿ��NJ.'�@��v��3@ut$��!?Bc��<�@@�
�G�ٿj*�HK��@$�T!��3@��57�!?�(��`�@@�
�G�ٿj*�HK��@$�T!��3@��57�!?�(��`�@@�
�G�ٿj*�HK��@$�T!��3@��57�!?�(��`�@@�
�G�ٿj*�HK��@$�T!��3@��57�!?�(��`�@���Ӂٿ���D��@����Z�3@�܂�ߐ!?�y�h��@���Ӂٿ���D��@����Z�3@�܂�ߐ!?�y�h��@���|'�ٿ��4����@2Ӯ��3@��Ȓ��!?8��G���@���|'�ٿ��4����@2Ӯ��3@��Ȓ��!?8��G���@���|'�ٿ��4����@2Ӯ��3@��Ȓ��!?8��G���@���|'�ٿ��4����@2Ӯ��3@��Ȓ��!?8��G���@���|'�ٿ��4����@2Ӯ��3@��Ȓ��!?8��G���@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�ď���ٿ�n�d��@ŧ��W 4@�#��!?��[�+�@�S_�ٿ���;��@�iR+4@\٣嘐!?���E �@���rٿ����\��@�^���4@϶���!?������@���rٿ����\��@�^���4@϶���!?������@��cn��ٿ��(�A�@ō&Q�4@z7��Ӑ!?��~h�@��cn��ٿ��(�A�@ō&Q�4@z7��Ӑ!?��~h�@��ٿ�z�{i��@��lIP4@V|�*ѐ!?��[��@��ٿ�z�{i��@��lIP4@V|�*ѐ!?��[��@��ٿ�z�{i��@��lIP4@V|�*ѐ!?��[��@��ٿ�z�{i��@��lIP4@V|�*ѐ!?��[��@� �߁ٿ���rQ�@K`74@���\��!?�g|�U�@� �߁ٿ���rQ�@K`74@���\��!?�g|�U�@� �߁ٿ���rQ�@K`74@���\��!?�g|�U�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@�-�*փٿ2L?�@.�%M�4@��&��!?���T�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@Dm'Y�ٿ�b_o��@�I�4@����K�!?e�N��X�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@֛<�2�ٿLk�1��@;`��4@G���!?�j8R-M�@��O�ٿhK�$�f�@�u�4@��,	�!?��jIO�@��O�ٿhK�$�f�@�u�4@��,	�!?��jIO�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@�?W���ٿ���:c�@���ۿ4@�C��͐!?g<_l�@��8�ٿ��ò��@�>	��4@�)"�̐!?�e�A���@�s�҄ٿ�J�Q��@(���Q4@��{�!?���-�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@�B��(�ٿ�ْkVj�@�(� �4@�����!?���%�H�@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@^�#G��ٿ�K�d���@�R_KG4@Ю�'ݐ!?��iP���@�����ٿ��ә�@_��T4@b,�Fʐ!?�Ճ	V��@�����ٿ��ә�@_��T4@b,�Fʐ!?�Ճ	V��@�����ٿ��ә�@_��T4@b,�Fʐ!?�Ճ	V��@�����ٿ��ә�@_��T4@b,�Fʐ!?�Ճ	V��@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@V��V�ٿ h��nc�@R��4@p"	��!?�B�8�@�la	��ٿ�o�K�v�@#:� 4@T��!?�D���@�la	��ٿ�o�K�v�@#:� 4@T��!?�D���@�la	��ٿ�o�K�v�@#:� 4@T��!?�D���@�la	��ٿ�o�K�v�@#:� 4@T��!?�D���@�la	��ٿ�o�K�v�@#:� 4@T��!?�D���@Ifn�N�ٿݎ,�Z+�@G�0�#4@�8|%��!?�������@Ifn�N�ٿݎ,�Z+�@G�0�#4@�8|%��!?�������@Ifn�N�ٿݎ,�Z+�@G�0�#4@�8|%��!?�������@j���ٿ�Xߚ�Q�@w4�Z4@��%���!?��S(e�@j���ٿ�Xߚ�Q�@w4�Z4@��%���!?��S(e�@j���ٿ�Xߚ�Q�@w4�Z4@��%���!?��S(e�@j���ٿ�Xߚ�Q�@w4�Z4@��%���!?��S(e�@j���ٿ�Xߚ�Q�@w4�Z4@��%���!?��S(e�@�����ٿ���@d\�b 4@Xx�۟�!?� ���@�����ٿ���@d\�b 4@Xx�۟�!?� ���@�����ٿ���@d\�b 4@Xx�۟�!?� ���@�����ٿ���@d\�b 4@Xx�۟�!?� ���@�6ύy�ٿ�?���@��]b 4@9�=A��!?�ϡ��q�@�6ύy�ٿ�?���@��]b 4@9�=A��!?�ϡ��q�@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@l�8���ٿ����\��@��R{4@�)���!?��S���@+|=G�ٿ,��vO��@�,�by4@��4�!?Ƌ�L�@+|=G�ٿ,��vO��@�,�by4@��4�!?Ƌ�L�@+|=G�ٿ,��vO��@�,�by4@��4�!?Ƌ�L�@+|=G�ٿ,��vO��@�,�by4@��4�!?Ƌ�L�@+|=G�ٿ,��vO��@�,�by4@��4�!?Ƌ�L�@qf�@��ٿ����@|�	�D4@���!?d�b���@qf�@��ٿ����@|�	�D4@���!?d�b���@qf�@��ٿ����@|�	�D4@���!?d�b���@qf�@��ٿ����@|�	�D4@���!?d�b���@qf�@��ٿ����@|�	�D4@���!?d�b���@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@d�jn�ٿ���v��@�</W4@׺�ː!?�jd�8�@I6��ٿx4��K�@�9	��4@���+ݐ!?���EV��@Q3��ٿ�ksm�%�@�>Ma�4@��.�!?�9}$e��@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@)$��n�ٿ;��!UL�@��S��4@'��� �!?f����@���ٿ�B��v��@��i�e4@�£i�!?��#�m��@���ٿ�B��v��@��i�e4@�£i�!?��#�m��@���ٿ�B��v��@��i�e4@�£i�!?��#�m��@���ٿ�B��v��@��i�e4@�£i�!?��#�m��@�|���ٿp����@xw�M4@��m���!?�h�i�T�@�|���ٿp����@xw�M4@��m���!?�h�i�T�@�|���ٿp����@xw�M4@��m���!?�h�i�T�@�|���ٿp����@xw�M4@��m���!?�h�i�T�@�|���ٿp����@xw�M4@��m���!?�h�i�T�@�Fw6��ٿmC�و�@7�f�04@)>�9��!?�tC��8�@�Fw6��ٿmC�و�@7�f�04@)>�9��!?�tC��8�@�Fw6��ٿmC�و�@7�f�04@)>�9��!?�tC��8�@�Fw6��ٿmC�و�@7�f�04@)>�9��!?�tC��8�@�ð��ٿ���F��@�>�%�4@��W�q�!?��9����@�ð��ٿ���F��@�>�%�4@��W�q�!?��9����@�ð��ٿ���F��@�>�%�4@��W�q�!?��9����@�ð��ٿ���F��@�>�%�4@��W�q�!?��9����@�����ٿ��k>Bq�@j���4@@;r�w�!?��e��@�����ٿ��k>Bq�@j���4@@;r�w�!?��e��@N�,W�ٿ�njx���@C�j*O4@��w�!?����?�@�*����ٿ�%�J��@I[0�z4@�)3m�!?���f��@�*����ٿ�%�J��@I[0�z4@�)3m�!?���f��@�*����ٿ�%�J��@I[0�z4@�)3m�!?���f��@�*����ٿ�%�J��@I[0�z4@�)3m�!?���f��@�*����ٿ�%�J��@I[0�z4@�)3m�!?���f��@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@8ౡ��ٿ�:{�n��@�Vi�d4@�$���!?�J@�b�@�T���ٿġ����@�ǥ�4@�#���!?6�-�R�@�T���ٿġ����@�ǥ�4@�#���!?6�-�R�@�T���ٿġ����@�ǥ�4@�#���!?6�-�R�@�T���ٿġ����@�ǥ�4@�#���!?6�-�R�@�!�֮�ٿ_���W��@�*y4@��3."�!?R���s�@�!�֮�ٿ_���W��@�*y4@��3."�!?R���s�@�g�p��ٿ�	6�!Q�@�WS6�4@��XW�!?���6q��@�g�p��ٿ�	6�!Q�@�WS6�4@��XW�!?���6q��@m�����ٿ�g���@g���m4@�h�?��!?�����@m�����ٿ�g���@g���m4@�h�?��!?�����@m�����ٿ�g���@g���m4@�h�?��!?�����@m�����ٿ�g���@g���m4@�h�?��!?�����@m�����ٿ�g���@g���m4@�h�?��!?�����@m�����ٿ�g���@g���m4@�h�?��!?�����@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@	���ٿQu�OO��@���{�4@�ө��!?:m�Sȴ�@�� ���ٿ�ʪ��$�@)EXv4@H�y���!?`�G Dk�@��:��ٿ���9�@.rC</4@�E��!?Z�'S̵�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@aq�;�ٿ�	+����@��DBq4@���!?�=�r^[�@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@����ٿ�X����@�	�4@9,+c��!?#�}X��@��<�ٿ��N���@���4@�qu��!?�p�Y�@��<�ٿ��N���@���4@�qu��!?�p�Y�@4GN��ٿ�Y�=6��@Ko鵟4@)�ݫy�!?����w@�@4GN��ٿ�Y�=6��@Ko鵟4@)�ݫy�!?����w@�@4GN��ٿ�Y�=6��@Ko鵟4@)�ݫy�!?����w@�@4GN��ٿ�Y�=6��@Ko鵟4@)�ݫy�!?����w@�@�\,M�ٿWPI�,��@�]m�	4@��`��!?�����G�@�\,M�ٿWPI�,��@�]m�	4@��`��!?�����G�@�\,M�ٿWPI�,��@�]m�	4@��`��!?�����G�@�\,M�ٿWPI�,��@�]m�	4@��`��!?�����G�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@�H�Qߊٿ<�o5�@�lF��4@-n����!?���._�@جN�|�ٿ��^�}��@㬩_�4@�T���!?���[�s�@جN�|�ٿ��^�}��@㬩_�4@�T���!?���[�s�@�ͯ�s�ٿc?8z/�@[����4@����ǐ!? ��N�@�ͯ�s�ٿc?8z/�@[����4@����ǐ!? ��N�@�ͯ�s�ٿc?8z/�@[����4@����ǐ!? ��N�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@���閄ٿ���I<9�@X���4@2�7�Ő!?�G��/�@,j"�ٿTizZ�@�*�G74@}����!?^���*��@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@e�?��~ٿ�)Vs��@=Ƽ�>4@�� �Ɛ!?גn�zG�@�Z����ٿ�#ϗ�\�@��BhY4@�Y�Ő!?+�i�Fa�@�Z����ٿ�#ϗ�\�@��BhY4@�Y�Ő!?+�i�Fa�@�Z����ٿ�#ϗ�\�@��BhY4@�Y�Ő!?+�i�Fa�@7$++߇ٿ�8෢p�@�0�l4@m�0���!?F~p�@��@7$++߇ٿ�8෢p�@�0�l4@m�0���!?F~p�@��@7$++߇ٿ�8෢p�@�0�l4@m�0���!?F~p�@��@�&�Qt�ٿ�7<�3�@�}�4@�/	߯�!?f��'�o�@�&�Qt�ٿ�7<�3�@�}�4@�/	߯�!?f��'�o�@�&�Qt�ٿ�7<�3�@�}�4@�/	߯�!?f��'�o�@�&�Qt�ٿ�7<�3�@�}�4@�/	߯�!?f��'�o�@�&�Qt�ٿ�7<�3�@�}�4@�/	߯�!?f��'�o�@�d�H�ٿd���:�@��ގ4@�+�9��!?1�D�4�@���#�ٿl
�CuP�@M�I��4@a��b�!?�f�sxv�@��R�|ٿ vU�h9�@�E�4@��vU��!?Q��a�@��R�|ٿ vU�h9�@�E�4@��vU��!?Q��a�@��R�|ٿ vU�h9�@�E�4@��vU��!?Q��a�@�_�8X}ٿS�nfo�@c�M9	4@E L�А!?++��Á�@�_�8X}ٿS�nfo�@c�M9	4@E L�А!?++��Á�@�_�8X}ٿS�nfo�@c�M9	4@E L�А!?++��Á�@aGe-{ٿ%���	�@���WO4@~c͐!?���f�@t[�D��ٿ:�W��@�@�JeA�4@���g�!?;u��\Q�@t[�D��ٿ:�W��@�@�JeA�4@���g�!?;u��\Q�@t[�D��ٿ:�W��@�@�JeA�4@���g�!?;u��\Q�@t[�D��ٿ:�W��@�@�JeA�4@���g�!?;u��\Q�@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@mR�ٿ2��"�@��4@����\�!?�ى���@�����ٿ�m�gV��@F�`�"4@�an\��!?�O��}d�@�����ٿ�m�gV��@F�`�"4@�an\��!?�O��}d�@�����ٿ�m�gV��@F�`�"4@�an\��!?�O��}d�@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�+W��ٿ�N�O��@�89��4@2�G�!?$�~���@�k�ٿZ.����@I���Y4@��gC�!?��մ��@4�7O͈ٿ����'�@Z`���4@�p����!?|�$��@��u�ٿ����T��@O`0��4@�S2:��!?�}��,�@��u�ٿ����T��@O`0��4@�S2:��!?�}��,�@��u�ٿ����T��@O`0��4@�S2:��!?�}��,�@��u�ٿ����T��@O`0��4@�S2:��!?�}��,�@� x)�ٿ���*�@�/�4@�w.���!?l?~�n�@m�I`�ٿ���+��@���*�4@o^ǝ��!?�u�F�(�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@}�%�ٿ+��g�@:��K�4@�#�^��!?�p�f%�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@�:3���ٿ�"��P�@���4@%}
���!?1�xƯ�@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@���ІٿE�@��@=wZ�4@.<����!?=�����@.��뎂ٿ�k���@{���4@8���!?���G��@.��뎂ٿ�k���@{���4@8���!?���G��@d��b�ٿ业���@���?4@�^`�Ԑ!?�s�X(�@d��b�ٿ业���@���?4@�^`�Ԑ!?�s�X(�@�
ժ�ٿ�h\s�@���׆4@Lm�Y�!?���L��@�
ժ�ٿ�h\s�@���׆4@Lm�Y�!?���L��@�
ժ�ٿ�h\s�@���׆4@Lm�Y�!?���L��@�
ժ�ٿ�h\s�@���׆4@Lm�Y�!?���L��@�
ժ�ٿ�h\s�@���׆4@Lm�Y�!?���L��@g�eȻ�ٿ]��J�@�Ԩ4@k3ҩ��!?92��Y��@g�eȻ�ٿ]��J�@�Ԩ4@k3ҩ��!?92��Y��@ ��~ٿ����z��@�����4@
�~��!?ewx����@ ��~ٿ����z��@�����4@
�~��!?ewx����@ ��~ٿ����z��@�����4@
�~��!?ewx����@ ��~ٿ����z��@�����4@
�~��!?ewx����@ ��~ٿ����z��@�����4@
�~��!?ewx����@ ��~ٿ����z��@�����4@
�~��!?ewx����@����ٿ��9���@{BW[
4@�O͐!?G�����@����ٿ��9���@{BW[
4@�O͐!?G�����@����ٿ��9���@{BW[
4@�O͐!?G�����@��?�5�ٿ	2�r\b�@O�B0�4@iw!t�!?�����n�@��?�5�ٿ	2�r\b�@O�B0�4@iw!t�!?�����n�@��?�5�ٿ	2�r\b�@O�B0�4@iw!t�!?�����n�@��?�5�ٿ	2�r\b�@O�B0�4@iw!t�!?�����n�@��?�5�ٿ	2�r\b�@O�B0�4@iw!t�!?�����n�@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@�����ٿ�)H>��@���� 4@�?5�4�!?��[
I��@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@S����ٿ@gs����@4��|4@{}�Tʐ!?eg���@,$�{ٿ.m�7c��@�'�4@$��Uې!?��ЗG�@,$�{ٿ.m�7c��@�'�4@$��Uې!?��ЗG�@��7WzٿY�'|,��@f�^��4@����Ȑ!?�t�Z�H�@��7WzٿY�'|,��@f�^��4@����Ȑ!?�t�Z�H�@��7WzٿY�'|,��@f�^��4@����Ȑ!?�t�Z�H�@��p�"ٿ��u
��@Kk��4@B�&:�!?��e�Ѿ�@��p�"ٿ��u
��@Kk��4@B�&:�!?��e�Ѿ�@��p�"ٿ��u
��@Kk��4@B�&:�!?��e�Ѿ�@���F�ٿ�{(����@��j�Q4@����͐!?1��h�	�@���F�ٿ�{(����@��j�Q4@����͐!?1��h�	�@��rMٿ�:)�,@�@��w|�4@�"a��!?�Z����@��rMٿ�:)�,@�@��w|�4@�"a��!?�Z����@��rMٿ�:)�,@�@��w|�4@�"a��!?�Z����@��rMٿ�:)�,@�@��w|�4@�"a��!?�Z����@��rMٿ�:)�,@�@��w|�4@�"a��!?�Z����@"�$��ٿ�Ub�T�@{�G�� 4@��,��!?���r�!�@"�$��ٿ�Ub�T�@{�G�� 4@��,��!?���r�!�@��u*Àٿ�7̷���@A�q"g�3@iW�ཐ!?��6� �@��u*Àٿ�7̷���@A�q"g�3@iW�ཐ!?��6� �@��u*Àٿ�7̷���@A�q"g�3@iW�ཐ!?��6� �@��u*Àٿ�7̷���@A�q"g�3@iW�ཐ!?��6� �@���ٿ�zƉC_�@�0�� 4@M�	��!?B��>l5�@�^2~ٿR��^�@����4@Đ�@�!?-Q��	�@�^2~ٿR��^�@����4@Đ�@�!?-Q��	�@�^2~ٿR��^�@����4@Đ�@�!?-Q��	�@�}w��ٿ`e>N�@�a�4[4@e�z��!?�OD��8�@�}w��ٿ`e>N�@�a�4[4@e�z��!?�OD��8�@�}w��ٿ`e>N�@�a�4[4@e�z��!?�OD��8�@�}w��ٿ`e>N�@�a�4[4@e�z��!?�OD��8�@"�9Նٿ��n����@�Lz4@�`�߆�!?��L����@"�9Նٿ��n����@�Lz4@�`�߆�!?��L����@"�9Նٿ��n����@�Lz4@�`�߆�!?��L����@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@�[WLʂٿ��'�@'sY)4@�?���!?�h7���@v�y}ٿ)��Q���@�u|4@�HgQ��!?xL���@pYɘՀٿ>��Dy�@&Vi\�4@
3Wp�!?vg8q@��@k�v�ٿ}'��s�@�j4@��C��!?��	��@k�v�ٿ}'��s�@�j4@��C��!?��	��@k�v�ٿ}'��s�@�j4@��C��!?��	��@k�v�ٿ}'��s�@�j4@��C��!?��	��@p��"�{ٿM���\�@"T���4@�*����!?��4��@p��"�{ٿM���\�@"T���4@�*����!?��4��@p��"�{ٿM���\�@"T���4@�*����!?��4��@dw�`wٿ�{R����@y���3@b(��!?�VT� �@dw�`wٿ�{R����@y���3@b(��!?�VT� �@ �1�wٿ;>����@e�-�4@�em��!?�<���@ �1�wٿ;>����@e�-�4@�em��!?�<���@ �1�wٿ;>����@e�-�4@�em��!?�<���@y:M��ٿb�ɖ�@���FB4@�����!?Qx����@y:M��ٿb�ɖ�@���FB4@�����!?Qx����@�ׄ<�ٿK��+�@I'>��4@a1�!?(�\����@ƨ���ٿ�%~z��@�}0�74@W�s�!?k�����@�:��ևٿLo��I��@@�P�i4@St�.�!?��l%��@�:��ևٿLo��I��@@�P�i4@St�.�!?��l%��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@8�>'5�ٿ���Q"��@�G�4@J���!?�i=GP��@{q�h̏ٿ/�����@�I%�4@�#��!?��1���@{q�h̏ٿ/�����@�I%�4@�#��!?��1���@*ɝ�6�ٿ���@�cq�4@��!���!?8��%�@*ɝ�6�ٿ���@�cq�4@��!���!?8��%�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@g�sO�ٿ���:�@g�^.q4@;l7�!?�i�E�@.��
�ٿX�e�ow�@6�V4@�	�!?�7�d(��@.��
�ٿX�e�ow�@6�V4@�	�!?�7�d(��@.��
�ٿX�e�ow�@6�V4@�	�!?�7�d(��@(/�?ňٿ�r�����@����N4@�mِ!?�U��@(/�?ňٿ�r�����@����N4@�mِ!?�U��@(/�?ňٿ�r�����@����N4@�mِ!?�U��@��0���ٿ��]~��@Y)F-4@Sh�!�!?�3�5+��@iy�"�ٿV��;��@�r���4@� �c��!?�VM�S�@iy�"�ٿV��;��@�r���4@� �c��!?�VM�S�@iy�"�ٿV��;��@�r���4@� �c��!?�VM�S�@�;"�$�ٿ�M]��h�@w�ґ4@�5��!?��3����@�;"�$�ٿ�M]��h�@w�ґ4@�5��!?��3����@�;"�$�ٿ�M]��h�@w�ґ4@�5��!?��3����@�;"�$�ٿ�M]��h�@w�ґ4@�5��!?��3����@��9�ԃٿ�G����@7'�E�3@�,����!?a�Qi���@��9�ԃٿ�G����@7'�E�3@�,����!?a�Qi���@��9�ԃٿ�G����@7'�E�3@�,����!?a�Qi���@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@2;4�U�ٿ{4(8��@�磊+4@���Ӑ!?�7,����@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@>1�ÃٿU�ܢW��@G��a�4@I��!?^�^�A�@�5���ٿ"�����@�k:���3@�!?��L���@�5���ٿ"�����@�k:���3@�!?��L���@�5���ٿ"�����@�k:���3@�!?��L���@�5���ٿ"�����@�k:���3@�!?��L���@�˄jȍٿ0�s7��@V#@�W4@��ѐ!?<�7���@�˄jȍٿ0�s7��@V#@�W4@��ѐ!?<�7���@�˄jȍٿ0�s7��@V#@�W4@��ѐ!?<�7���@�˄jȍٿ0�s7��@V#@�W4@��ѐ!?<�7���@�|�%��ٿ��'9���@<�Zc�4@�5�!?=��6~|�@�|�%��ٿ��'9���@<�Zc�4@�5�!?=��6~|�@�|�%��ٿ��'9���@<�Zc�4@�5�!?=��6~|�@�|�%��ٿ��'9���@<�Zc�4@�5�!?=��6~|�@�_�Ȏ�ٿ4���y��@M�h�4@��/*�!?��8�&L�@�_�Ȏ�ٿ4���y��@M�h�4@��/*�!?��8�&L�@�&@L�ٿ����0�@��Y��4@C~?�!? 7��fZ�@�&@L�ٿ����0�@��Y��4@C~?�!? 7��fZ�@^��Q�ٿʝ�߳;�@�q���4@p�矫�!?�P){�@^��Q�ٿʝ�߳;�@�q���4@p�矫�!?�P){�@��h#�ٿE�'���@�� U4@�����!?]z�L�&�@��h#�ٿE�'���@�� U4@�����!?]z�L�&�@��h#�ٿE�'���@�� U4@�����!?]z�L�&�@�:�OQ�ٿ�k\��@ ��M�4@�͞mҐ!?�H����@�:�OQ�ٿ�k\��@ ��M�4@�͞mҐ!?�H����@�:�OQ�ٿ�k\��@ ��M�4@�͞mҐ!?�H����@���{�ٿ�]sK��@4�㩉4@uVv
q�!?�Z��Rv�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@cLM���ٿ��1b,��@g�C(�4@�敭�!?v9�ʡ�@�~a6�ٿ�9��{�@ɝ���4@�B��Ő!?��ab��@�~a6�ٿ�9��{�@ɝ���4@�B��Ő!?��ab��@�~a6�ٿ�9��{�@ɝ���4@�B��Ő!?��ab��@�~a6�ٿ�9��{�@ɝ���4@�B��Ő!?��ab��@�~a6�ٿ�9��{�@ɝ���4@�B��Ő!?��ab��@0����ٿ�l���@A��Ti4@db�1��!?�ғ(A��@0����ٿ�l���@A��Ti4@db�1��!?�ғ(A��@0����ٿ�l���@A��Ti4@db�1��!?�ғ(A��@�z�
�ٿ{nj��;�@����m4@{���~�!?��8��M�@�z�
�ٿ{nj��;�@����m4@{���~�!?��8��M�@�2�Ѝ�ٿ-�����@�Hǩ4@m|
���!?4J�" k�@����ٿD*W���@�Ϣ��4@��慒�!?�%�3�@����ٿD*W���@�Ϣ��4@��慒�!?�%�3�@����ٿD*W���@�Ϣ��4@��慒�!?�%�3�@F�,�ٿ��)��@TM�c(4@MSﺐ!?�"j9��@F�,�ٿ��)��@TM�c(4@MSﺐ!?�"j9��@F�,�ٿ��)��@TM�c(4@MSﺐ!?�"j9��@F�,�ٿ��)��@TM�c(4@MSﺐ!?�"j9��@F�,�ٿ��)��@TM�c(4@MSﺐ!?�"j9��@�>.�ٿ�v�~�!�@_���4@>F��!?'�����@�����ٿ-��F���@;S�64@��Đ!?�A���@�����ٿ-��F���@;S�64@��Đ!?�A���@�(�`�ٿ�t���@	�S
4@��6���!?����/�@�(�`�ٿ�t���@	�S
4@��6���!?����/�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@��M��ٿ��_m�B�@T���4@�����!?���t <�@�9�͈ٿ�tQ'��@^��Z;4@�;A���!?���H��@�9�͈ٿ�tQ'��@^��Z;4@�;A���!?���H��@��g�ٿC�R�p�@� J��4@�᥯�!?�܂��Y�@��g�ٿC�R�p�@� J��4@�᥯�!?�܂��Y�@��g�ٿC�R�p�@� J��4@�᥯�!?�܂��Y�@��g�ٿC�R�p�@� J��4@�᥯�!?�܂��Y�@��g�ٿC�R�p�@� J��4@�᥯�!?�܂��Y�@ ��7��ٿ�5v����@o7O�4@3r�;��!?1�����@ ��7��ٿ�5v����@o7O�4@3r�;��!?1�����@�w� ٿ���VZ�@Zc2�4@UP��!?Rx���@�w� ٿ���VZ�@Zc2�4@UP��!?Rx���@�H�ٿI�ȡ*z�@E*Y�4@� �@�!?��{_��@�H�ٿI�ȡ*z�@E*Y�4@� �@�!?��{_��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�};m��ٿ�Q����@�5�M�4@IL���!?ڛ羗��@�妳V�ٿ�6ߡ�<�@� 
-4@|Ԓ���!?�'��.2�@�妳V�ٿ�6ߡ�<�@� 
-4@|Ԓ���!?�'��.2�@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@ޛ��{�ٿ�i�,�@5n���4@��mǐ!?������@W�?=׆ٿ\'�H�l�@5t�Q4@ˮw�!?�e���I�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@)�4i�ٿ�}{+���@�	�C�4@����!?�)f1�D�@	��v�ٿʸ�ގ�@� �-4@y�̘�!?mC�*Y�@���&�ٿ�׺�)2�@oW��4@u5��!?#���x/�@���&�ٿ�׺�)2�@oW��4@u5��!?#���x/�@���&�ٿ�׺�)2�@oW��4@u5��!?#���x/�@���&�ٿ�׺�)2�@oW��4@u5��!?#���x/�@w��鬋ٿ�3R�_��@���I4@<�y�Ґ!?������@��8�_�ٿ-��c��@D��� 4@�,r��!?' y�/�@��8�_�ٿ-��c��@D��� 4@�,r��!?' y�/�@��8�_�ٿ-��c��@D��� 4@�,r��!?' y�/�@��8�_�ٿ-��c��@D��� 4@�,r��!?' y�/�@��8�_�ٿ-��c��@D��� 4@�,r��!?' y�/�@�����ٿ�;3���@@{-<;4@ke�!?�Jıta�@�����ٿ�;3���@@{-<;4@ke�!?�Jıta�@^�UI�ٿAW��KK�@!�Y�H4@��շ�!?K����@��t1̄ٿgT҂���@����4@'����!? )���m�@��t1̄ٿgT҂���@����4@'����!? )���m�@��t1̄ٿgT҂���@����4@'����!? )���m�@��t1̄ٿgT҂���@����4@'����!? )���m�@,�D惆ٿ���y�=�@���S�4@Is��h�!?cݟ#B�@Q����ٿ�'��Z�@l��4@��J�j�!?��#܁�@%q)sz�ٿG�?!���@b��$4@���I�!?+�R���@��];��ٿ�Rz��u�@[�u&��3@�l2cK�!?��m�n��@}{�Ĝ�ٿ:��b{P�@����3@9NbR��!?�lpu�@��?.�ٿ� �.?�@)�;MA4@���!?Pȁ&���@��?.�ٿ� �.?�@)�;MA4@���!?Pȁ&���@��?.�ٿ� �.?�@)�;MA4@���!?Pȁ&���@3�Z�ٿ�S���@��Y94@K#���!?�d�����@3�Z�ٿ�S���@��Y94@K#���!?�d�����@3�Z�ٿ�S���@��Y94@K#���!?�d�����@3�Z�ٿ�S���@��Y94@K#���!?�d�����@�;�J�ٿ��?�x��@P]�B� 4@�!�Uΐ!?br.��c�@�;�J�ٿ��?�x��@P]�B� 4@�!�Uΐ!?br.��c�@�;�J�ٿ��?�x��@P]�B� 4@�!�Uΐ!?br.��c�@�;�J�ٿ��?�x��@P]�B� 4@�!�Uΐ!?br.��c�@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@����ٿ��FR��@�lV&4@�4��!?�o�����@<_>N�ٿ����@:U��	4@�o��Ɛ!?�,�77�@<_>N�ٿ����@:U��	4@�o��Ɛ!?�,�77�@�Y���ٿN�l���@(f>�N	4@)o�� �!?%�L��@�Y���ٿN�l���@(f>�N	4@)o�� �!?%�L��@�Y���ٿN�l���@(f>�N	4@)o�� �!?%�L��@a����ٿ��e57��@iFM�A	4@IZ	Q�!?�#�,��@a����ٿ��e57��@iFM�A	4@IZ	Q�!?�#�,��@a����ٿ��e57��@iFM�A	4@IZ	Q�!?�#�,��@l�$��ٿ�k`��@��[4@Ր{X�!?D�P�Rv�@l�$��ٿ�k`��@��[4@Ր{X�!?D�P�Rv�@l�$��ٿ�k`��@��[4@Ր{X�!?D�P�Rv�@l�$��ٿ�k`��@��[4@Ր{X�!?D�P�Rv�@w�����ٿT��<�@W�_P�4@���[�!?���o ��@�m޽��ٿy\���J�@b\���4@�	���!?�P+����@si���ٿz��@�K� 4@~�H^��!?_4�^��@�B�D�ٿ(���@ ��4@�l�w�!?o�1�w�@lhF)�ٿB�כ��@x):P4@�D��!?v%�����@`y��ٿ������@a���44@�եX�!?^W���@`y��ٿ������@a���44@�եX�!?^W���@`y��ٿ������@a���44@�եX�!?^W���@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@M�۪��ٿ?�G_(�@����4@���̐!?"��N��@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@V�g?A�ٿ;Fk���@H��:84@@mĐ!?�&7���@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@�e��ٿ�f��3�@�4N4@4�;΅�!?%B�s��@��"u�ٿ�o���@��:��4@y�!?P1���@��"u�ٿ�o���@��:��4@y�!?P1���@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@N�yPP�ٿ_l{8��@�?>�4@ଋ:k�!?md�a�@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Lh}Çٿ����@����4@��~ʐ!?�ަ���@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@Ζ?Ɖٿyб���@O�	;4@�ƙ���!?ϵ �x�@pMY�ٿI�6���@��-�4@�&�*��!?�Z�ƨF�@��m��ٿ��2_{�@]64d�4@_Q�?��!?[dAr�@��m��ٿ��2_{�@]64d�4@_Q�?��!?[dAr�@�lcS�ٿ���0���@��!2�4@�"8uܐ!?�*wP�@�lcS�ٿ���0���@��!2�4@�"8uܐ!?�*wP�@t�[�f�ٿ�f=����@�-1g4@N �4��!?3���ch�@t�[�f�ٿ�f=����@�-1g4@N �4��!?3���ch�@t�[�f�ٿ�f=����@�-1g4@N �4��!?3���ch�@t�[�f�ٿ�f=����@�-1g4@N �4��!?3���ch�@t�[�f�ٿ�f=����@�-1g4@N �4��!?3���ch�@7�Z�ٿn���n�@p�W,4@����!?�p�hR�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@"0U��ٿׅ�g��@�2\°4@���%�!?�w�IF�@:�;菀ٿBj |N��@U���44@��x8�!?s%X�A��@:�;菀ٿBj |N��@U���44@��x8�!?s%X�A��@��@ٿ�a�[��@�@X&<4@O[Ĥ��!?J�P=%_�@��@ٿ�a�[��@�@X&<4@O[Ĥ��!?J�P=%_�@��@ٿ�a�[��@�@X&<4@O[Ĥ��!?J�P=%_�@��@ٿ�a�[��@�@X&<4@O[Ĥ��!?J�P=%_�@��@ٿ�a�[��@�@X&<4@O[Ĥ��!?J�P=%_�@{�ͮ�{ٿ���r���@SD���4@��W;��!?����8��@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@��r�|ٿ���6�@�`͚H4@ng�!?��<9���@KcU~a�ٿo�T/��@t�JwK4@l�R_P�!?��1�`H�@U7A��ٿ%ɖ���@�!��4@����!?�E�^��@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@���e�ٿ�x��w�@����4@�M#��!?<�����@�2~�C�ٿk|�j�u�@;$��4@�ϐ!?��c���@eet�ٿ�l|�Dk�@C�	�o4@R�����!?���6��@ ̠���ٿ��'�-�@ޯ�E�4@���Y�!?���QV��@ ̠���ٿ��'�-�@ޯ�E�4@���Y�!?���QV��@ ̠���ٿ��'�-�@ޯ�E�4@���Y�!?���QV��@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@�Ԛ�ǃٿ@���1��@���&�4@�   G�!?H��+�@����o�ٿ�U6,(��@�C,4@��%�s�!?6��w��@����o�ٿ�U6,(��@�C,4@��%�s�!?6��w��@�E����ٿ41P���@r4@���j�!?Ϋ�L���@�E����ٿ41P���@r4@���j�!?Ϋ�L���@�E����ٿ41P���@r4@���j�!?Ϋ�L���@����ٿ6\�����@d�	4@N[TU�!?�,J ���@����ٿ6\�����@d�	4@N[TU�!?�,J ���@����ٿ6\�����@d�	4@N[TU�!?�,J ���@�_�ٿ(�4" ��@`mK#4@����ϐ!?�/	��@�_�ٿ(�4" ��@`mK#4@����ϐ!?�/	��@�_�ٿ(�4" ��@`mK#4@����ϐ!?�/	��@Ga�_�ٿ������@\�~P4@X�����!?ڒ�K�@Ga�_�ٿ������@\�~P4@X�����!?ڒ�K�@'�MM�ٿz����@�+��4@K��'�!?
hj���@'�MM�ٿz����@�+��4@K��'�!?
hj���@'�MM�ٿz����@�+��4@K��'�!?
hj���@D&��o�ٿQؓ�>�@��n4@(�<��!?����9��@D&��o�ٿQؓ�>�@��n4@(�<��!?����9��@D&��o�ٿQؓ�>�@��n4@(�<��!?����9��@D&��o�ٿQؓ�>�@��n4@(�<��!?����9��@�2�|ٿ������@0�E��4@Ψ-o�!?��\��P�@�2�|ٿ������@0�E��4@Ψ-o�!?��\��P�@�2�|ٿ������@0�E��4@Ψ-o�!?��\��P�@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@F���|ٿ��>+���@���b4@Y����!?\�>҆��@�p�s �ٿ���l�@3☀M4@��E��!?9��	��@�p�s �ٿ���l�@3☀M4@��E��!?9��	��@�p�s �ٿ���l�@3☀M4@��E��!?9��	��@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@��!t�ٿ�r� &�@��f��4@Z����!?Gm�����@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@"0Ԛ�ٿ3�b��@��*#�4@�_jѐ!?���_�@`�,�ٿ�@�S�@/~��4@�<Q��!?6PH�@`�,�ٿ�@�S�@/~��4@�<Q��!?6PH�@`�,�ٿ�@�S�@/~��4@�<Q��!?6PH�@��w�c�ٿ��d�	�@���e4@�ɐ!?��9h��@��w�c�ٿ��d�	�@���e4@�ɐ!?��9h��@��w�c�ٿ��d�	�@���e4@�ɐ!?��9h��@��w�c�ٿ��d�	�@���e4@�ɐ!?��9h��@��Ӽ�ٿtWnh��@��(4@�Ф��!?�0&u��@��Ӽ�ٿtWnh��@��(4@�Ф��!?�0&u��@��-<��ٿ�\��`�@<��ն4@�3Y���!?�N�?�@��-<��ٿ�\��`�@<��ն4@�3Y���!?�N�?�@��-<��ٿ�\��`�@<��ն4@�3Y���!?�N�?�@��-<��ٿ�\��`�@<��ն4@�3Y���!?�N�?�@���嬎ٿh�N��H�@�ڦ]�4@����!?��11w�@�����ٿ�gfL�*�@��8@4@p���p�!?Q)����@(0)�ٿgn���H�@S�`�`4@��kBn�!?���,�@(0)�ٿgn���H�@S�`�`4@��kBn�!?���,�@(0)�ٿgn���H�@S�`�`4@��kBn�!?���,�@�Va�ӊٿ���eT�@Qz[��3@\�ܲ��!?�<R��<�@�Va�ӊٿ���eT�@Qz[��3@\�ܲ��!?�<R��<�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@��U�Ԁٿ�.V���@h�@^ 4@��[�!?Vj�Ӌ�@�:�,�ٿ��B�S�@��6>�4@��6���!?�Z�N��@�:�,�ٿ��B�S�@��6>�4@��6���!?�Z�N��@� i�ٿ��^��@��*�4@�Qݚ�!?���g��@� i�ٿ��^��@��*�4@�Qݚ�!?���g��@� i�ٿ��^��@��*�4@�Qݚ�!?���g��@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�q���ٿ��?��o�@��4@ns��Ր!?�1����@�4"��ٿ�vX��@���4@b�,ǐ!?���w���@�4"��ٿ�vX��@���4@b�,ǐ!?���w���@�4"��ٿ�vX��@���4@b�,ǐ!?���w���@{H��N�ٿs�_���@�;�4@��ѐ!?��S���@{H��N�ٿs�_���@�;�4@��ѐ!?��S���@{H��N�ٿs�_���@�;�4@��ѐ!?��S���@{H��N�ٿs�_���@�;�4@��ѐ!?��S���@{H��N�ٿs�_���@�;�4@��ѐ!?��S���@t���ٿ����BE�@���2�4@Q�1#��!?'3�9��@t���ٿ����BE�@���2�4@Q�1#��!?'3�9��@t���ٿ����BE�@���2�4@Q�1#��!?'3�9��@�-��f�ٿ<�L��@7��f4@n/!?OH?��C�@!��Ϗٿ�����s�@�F4�4@��@��!?���!>��@K���ٿ�K5�s�@W=g�4@8����!?Md����@K���ٿ�K5�s�@W=g�4@8����!?Md����@K���ٿ�K5�s�@W=g�4@8����!?Md����@\��?m�ٿ���R�@&j0��4@�2���!?����A�@4	e��ٿ������@(��4@y<��!?��ï�@4	e��ٿ������@(��4@y<��!?��ï�@4	e��ٿ������@(��4@y<��!?��ï�@4	e��ٿ������@(��4@y<��!?��ï�@4	e��ٿ������@(��4@y<��!?��ï�@4	e��ٿ������@(��4@y<��!?��ï�@�5��ߐٿq�q��@�O0R24@F5t���!?���u;��@�5��ߐٿq�q��@�O0R24@F5t���!?���u;��@c��p�ٿU�.im�@N�eS�4@}����!?+�^ce�@c��p�ٿU�.im�@N�eS�4@}����!?+�^ce�@c��p�ٿU�.im�@N�eS�4@}����!?+�^ce�@c��p�ٿU�.im�@N�eS�4@}����!?+�^ce�@c��p�ٿU�.im�@N�eS�4@}����!?+�^ce�@N�̎�ٿ)�/�~�@�=�4�4@��>�!?��
���@N�̎�ٿ)�/�~�@�=�4�4@��>�!?��
���@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@;w���ٿa���L�@z�ACW4@@��͐!?���yi]�@�`���ٿ�j�*y[�@�a�Ժ4@%�I���!?'��G�`�@�`���ٿ�j�*y[�@�a�Ժ4@%�I���!?'��G�`�@ǭA�ٿ���E�@�R]
�4@�=a��!?:^��-�@ǭA�ٿ���E�@�R]
�4@�=a��!?:^��-�@ǭA�ٿ���E�@�R]
�4@�=a��!?:^��-�@h)^��ٿ��4Xu��@R� "�4@�L|��!?����r��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@�ii���ٿ^V��&�@�d	J�4@-��#��!??k�H8��@hUi�2�ٿ�]�0G3�@ �# ^4@�Gy�j�!?H�!M"�@8n&+�ٿf�V2M0�@�v�4@���k�!?��Š��@8n&+�ٿf�V2M0�@�v�4@���k�!?��Š��@8n&+�ٿf�V2M0�@�v�4@���k�!?��Š��@�m�}ٿ�>+�_��@�+��4@ڝHf��!?px�U�@�m�}ٿ�>+�_��@�+��4@ڝHf��!?px�U�@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@�`<�ٿ�f�D��@��4@Ԫ��z�!?Tl�*U��@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@E]1]�ٿ�b4���@��fU�4@z�r��!?(���T�@�&�"ٿ��7]�@wo7�4@Ѳ4���!?X#x�ʥ�@�&�"ٿ��7]�@wo7�4@Ѳ4���!?X#x�ʥ�@���Le�ٿڛ��d��@{�[l"4@�m�f�!?�x8���@��{&��ٿ��F% ��@o�L�84@q�"��!?Ȇ{�C��@��{&��ٿ��F% ��@o�L�84@q�"��!?Ȇ{�C��@��{&��ٿ��F% ��@o�L�84@q�"��!?Ȇ{�C��@��{&��ٿ��F% ��@o�L�84@q�"��!?Ȇ{�C��@��{&��ٿ��F% ��@o�L�84@q�"��!?Ȇ{�C��@�V���ٿ+��I��@F/
,�4@/�"��!?u��k��@S㨅�ٿ �M��@�b��,4@r�=
�!?�ͭ~��@S㨅�ٿ �M��@�b��,4@r�=
�!?�ͭ~��@S㨅�ٿ �M��@�b��,4@r�=
�!?�ͭ~��@S㨅�ٿ �M��@�b��,4@r�=
�!?�ͭ~��@S㨅�ٿ �M��@�b��,4@r�=
�!?�ͭ~��@��I܉ٿ�{�7�@�Ĭ�a4@�����!?�q�IK\�@Xwצ$�ٿ�kbU=��@�CM�4@
�U��!?���1�X�@Xwצ$�ٿ�kbU=��@�CM�4@
�U��!?���1�X�@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@V�nr��ٿk�鄬�@�E��+4@aj)N��!?��|���@7�.�ٿL�r��@0 �4@��B0��!?B�����@|6SH�ٿ�����@Q9���4@t!5ې!?2�����@|6SH�ٿ�����@Q9���4@t!5ې!?2�����@|6SH�ٿ�����@Q9���4@t!5ې!?2�����@d�vCy�ٿ�F��j��@��`I4@����!?�1��k��@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���ٿa�����@),c%G4@��y	��!?M��T#Q�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@���|΅ٿ}O��O��@�C�&4@7�.{��!?�&�%�@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@�׽�s�ٿb�]"Ū�@�3��:4@�$��Đ!?t0����@���S|�ٿ�rUY�@O��� 4@Xp����!?n�;���@���S|�ٿ�rUY�@O��� 4@Xp����!?n�;���@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@#W��Ձٿ�fA�4�@� �94@��GZ��!?�#�`�@�)(]�zٿ9ج�?��@�ra�4@6Z�(ސ!?f�/�r�@�>�Ayٿ�o�E���@���#4@�����!?|ߔ��@�>�Ayٿ�o�E���@���#4@�����!?|ߔ��@XDs{ٿP�OX%=�@bq���4@sit�!?�YF��A�@XDs{ٿP�OX%=�@bq���4@sit�!?�YF��A�@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@�s��/vٿPv��a#�@G%�
�4@�~��!?��)]��@����zٿ��7R�@����4@ϊ���!?�b�W?�@����zٿ��7R�@����4@ϊ���!?�b�W?�@0�2IG�ٿ-��~�@$�h� 4@R셩А!?Ԑ���i�@h�n+�ٿe�
�:�@�lkћ4@�N�J�!?C����~�@��#�ٿWS���@� ��-4@��؄ݐ!?����z��@��#�ٿWS���@� ��-4@��؄ݐ!?����z��@��#�ٿWS���@� ��-4@��؄ݐ!?����z��@��#�ٿWS���@� ��-4@��؄ݐ!?����z��@��#�ٿWS���@� ��-4@��؄ݐ!?����z��@Ln9��ٿQ��UM��@�+�~4@H��1ؐ!?�,va��@Ln9��ٿQ��UM��@�+�~4@H��1ؐ!?�,va��@Ln9��ٿQ��UM��@�+�~4@H��1ؐ!?�,va��@Ln9��ٿQ��UM��@�+�~4@H��1ؐ!?�,va��@����~ٿ���v��@F�5 4@
,�X�!?uh�k]�@����~ٿ���v��@F�5 4@
,�X�!?uh�k]�@Gv%�d�ٿ?G]$���@�����3@i����!?� ]���@qJ��%{ٿ�*����@���U4@Z���!?�ß0���@5d�)�ٿ8�*;���@��)�4@ff#��!?�\C���@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@.2@�ٿd��t��@H	�4@�W�~�!?S�	��V�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@��%h�ٿ��cʆ�@aK�pF4@g5>��!?�1� �<�@L����ٿ섛�jl�@pyS�4@e�#�!?�o���@�&<��ٿ�q�]�#�@�T0�|4@�.N��!?$9����@�&<��ٿ�q�]�#�@�T0�|4@�.N��!?$9����@�	r���ٿ�*��2�@�N�p4@@�ǥ/�!?S�
N��@�	r���ٿ�*��2�@�N�p4@@�ǥ/�!?S�
N��@rҦ8�ٿ��<�s�@�����4@���ِ!? $��ct�@�A�ٿ��6-5�@[#�À4@e�:H�!?&W�K��@6y"���ٿ���#Qg�@�>��4@�e�-̐!?���Ai�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@q�7J؃ٿ������@3�al4@������!?S/G�t�@���ٿ ֓+��@��ⲍ4@��>[�!?n�W�@���ٿ ֓+��@��ⲍ4@��>[�!?n�W�@���ٿ ֓+��@��ⲍ4@��>[�!?n�W�@�B%:[�ٿ�{E^��@���g�4@��bN�!?�k8����@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@(Ǩ��ٿ�ҭ]�@3�G�P4@�O���!?��U���@��fz�ٿs��x�Q�@v���w4@���3�!?�� ��@��fz�ٿs��x�Q�@v���w4@���3�!?�� ��@��fz�ٿs��x�Q�@v���w4@���3�!?�� ��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@�V����ٿ�H?p���@�&N7f4@N^Z�!?��T��@X-.�w�ٿ*�M���@�T"�4@x� =�!?00��B�@X-.�w�ٿ*�M���@�T"�4@x� =�!?00��B�@�'���ٿ��o16�@p�!4@C}�=%�!?S��"�J�@�'���ٿ��o16�@p�!4@C}�=%�!?S��"�J�@��#R��ٿ��V���@��$΂4@?�׎O�!?�\w�{+�@�Տ#�ٿ�/��@\���4@����l�!?���cW��@cyA�ٿ��B�6?�@�_{�I4@̞�!?�*��>��@cyA�ٿ��B�6?�@�_{�I4@̞�!?�*��>��@cyA�ٿ��B�6?�@�_{�I4@̞�!?�*��>��@cyA�ٿ��B�6?�@�_{�I4@̞�!?�*��>��@cyA�ٿ��B�6?�@�_{�I4@̞�!?�*��>��@�Ƅ�~ٿ�Eu!�@�+�4@V���!?IN����@�Ƅ�~ٿ�Eu!�@�+�4@V���!?IN����@�Ƅ�~ٿ�Eu!�@�+�4@V���!?IN����@�,3�ٿ�Qϟ���@�-/�4@ ����!?W}�t�@�,3�ٿ�Qϟ���@�-/�4@ ����!?W}�t�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@Ҹ��Ņٿ����y�@j|��4@uNo�!?�z�.,�@�3��ٿn����@>�4@�!�ſ�!?��p��@���v+�ٿ�Y�1��@���z_4@�����!?�-�z���@���v+�ٿ�Y�1��@���z_4@�����!?�-�z���@���v+�ٿ�Y�1��@���z_4@�����!?�-�z���@���v+�ٿ�Y�1��@���z_4@�����!?�-�z���@2�6ىٿ�ۯ���@eq�O4@�<��!?2p'%7��@2�6ىٿ�ۯ���@eq�O4@�<��!?2p'%7��@��	]�ٿ���<��@Z�u��
4@!]���!?��1&j�@��	]�ٿ���<��@Z�u��
4@!]���!?��1&j�@��	]�ٿ���<��@Z�u��
4@!]���!?��1&j�@��	]�ٿ���<��@Z�u��
4@!]���!?��1&j�@��	]�ٿ���<��@Z�u��
4@!]���!?��1&j�@P��/%�ٿ�/ ����@P����4@x��ai�!?�zS!��@P��/%�ٿ�/ ����@P����4@x��ai�!?�zS!��@P��/%�ٿ�/ ����@P����4@x��ai�!?�zS!��@���y�ٿ���q���@�Bg�4@~(K�!?:f)v���@���y�ٿ���q���@�Bg�4@~(K�!?:f)v���@���y�ٿ���q���@�Bg�4@~(K�!?:f)v���@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@��d�;�ٿ_k�oe}�@�q�� 4@D��l�!?
��@��@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@�,����ٿ����D�@�b.�f�3@9C��!?�o��jo�@唼��ٿko�6�D�@�;�]�3@A��f̐!?C����/�@�
ͪ��ٿd���[n�@��7��3@d�,!?��Y��@�b��ٿ9Z/�%�@���� 4@�F���!?�8�9��@�b��ٿ9Z/�%�@���� 4@�F���!?�8�9��@�b��ٿ9Z/�%�@���� 4@�F���!?�8�9��@�b��ٿ9Z/�%�@���� 4@�F���!?�8�9��@>��5�ٿ��,�g��@؀��7 4@���!?�Rh�$�@>��5�ٿ��,�g��@؀��7 4@���!?�Rh�$�@>��5�ٿ��,�g��@؀��7 4@���!?�Rh�$�@k�o#�ٿW���;�@3%N�^4@�ä��!?ah��5��@k�o#�ٿW���;�@3%N�^4@�ä��!?ah��5��@�,W5}ٿ�������@ j,3�4@����!?T��S��@�,W5}ٿ�������@ j,3�4@����!?T��S��@�,W5}ٿ�������@ j,3�4@����!?T��S��@�,W5}ٿ�������@ j,3�4@����!?T��S��@*V�*{ٿh����@�3I� 4@I4$]��!?��>��@*V�*{ٿh����@�3I� 4@I4$]��!?��>��@�?zٿ#�H���@"!q�4@�hC)�!?��u�i�@�?zٿ#�H���@"!q�4@�hC)�!?��u�i�@�?zٿ#�H���@"!q�4@�hC)�!?��u�i�@�?zٿ#�H���@"!q�4@�hC)�!?��u�i�@�?zٿ#�H���@"!q�4@�hC)�!?��u�i�@��,�
{ٿ�<�C��@\��/�4@�q�n��!?��q��]�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@�]��ٿ�y�g���@7\M�s4@x�m뷐!?�s�Q�@LD6���ٿ(�R�@G���4@	�K��!?�N�s[^�@LD6���ٿ(�R�@G���4@	�K��!?�N�s[^�@LD6���ٿ(�R�@G���4@	�K��!?�N�s[^�@q`��ٿ�x,+m��@	�#4@[g@�ؐ!?����[�@q`��ٿ�x,+m��@	�#4@[g@�ؐ!?����[�@q`��ٿ�x,+m��@	�#4@[g@�ؐ!?����[�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@���=݅ٿ���}�@]1��	4@L��z�!?9W ��D�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@� :�ٿ����e)�@^O�n4@c) 8��!?V��mV�@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@sT�c�ٿ-�P.�5�@����4@v�	�ː!?�����@��ɬn�ٿ�TA��X�@���1W4@k��(��!?n�ԃK��@��ɬn�ٿ�TA��X�@���1W4@k��(��!?n�ԃK��@B �9�ٿW��22�@�`�R�4@;���!?��V�M��@B �9�ٿW��22�@�`�R�4@;���!?��V�M��@B �9�ٿW��22�@�`�R�4@;���!?��V�M��@$@��ɇٿ�A��Jv�@��i"�4@��񏲐!?�S���@i�=�ٿ
�}���@�|"Na4@|f��Ɛ!?R���N'�@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@;"��"�ٿ��k�b��@Cz�o�4@A�^��!?<�g�L��@����ٿr������@��W� 4@e��Ő!?�.��6�@����ٿr������@��W� 4@e��Ő!?�.��6�@����ٿr������@��W� 4@e��Ő!?�.��6�@����ٿr������@��W� 4@e��Ő!?�.��6�@x��6�ٿ5$��3�@�/W�4@��p�!?M?���@x��6�ٿ5$��3�@�/W�4@��p�!?M?���@x��6�ٿ5$��3�@�/W�4@��p�!?M?���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��u�؅ٿ!>O(��@a���4@��y��!?�T�k���@��V�C�ٿq<7���@n�l-4@���nU�!?G0��6��@��V�C�ٿq<7���@n�l-4@���nU�!?G0��6��@��V�C�ٿq<7���@n�l-4@���nU�!?G0��6��@��V�C�ٿq<7���@n�l-4@���nU�!?G0��6��@��V�C�ٿq<7���@n�l-4@���nU�!?G0��6��@u�R�`�ٿ8�����@��gu4@�R�a�!?�I7۔�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@|.���ٿ�AC7K��@�`K�4@qDeAސ!?�9u	_�@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@Xpn�4�ٿ����-�@�<�m4@��>d�!?�)-���@�ߙ��ٿU1�h4I�@��04@fm7Ð!?{VX��`�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��d."�ٿ�i5Ki]�@�h/4@���ߐ!?z��40�@��y2��ٿt��*��@6��c44@z2(���!?�C���K�@��y2��ٿt��*��@6��c44@z2(���!?�C���K�@��y2��ٿt��*��@6��c44@z2(���!?�C���K�@��y2��ٿt��*��@6��c44@z2(���!?�C���K�@��%X��ٿ�w����@�����4@��AҐ!?��z&�\�@��%X��ٿ�w����@�����4@��AҐ!?��z&�\�@��%X��ٿ�w����@�����4@��AҐ!?��z&�\�@��%X��ٿ�w����@�����4@��AҐ!?��z&�\�@��%X��ٿ�w����@�����4@��AҐ!?��z&�\�@E��A}ٿ�ͪ���@W�ϸ� 4@��TTɐ!?
��@�@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@|ʮ���ٿܠj��@�;��*4@e ��H�!?a�����@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@�,�{M�ٿ�7O��@8&V-�4@�9w�Q�!?�O�gw��@N��#�ٿ��b%�@۪E�4@�b&��!?Ꮌ@���@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@2�Oˊٿ�=�\@�@�H��u4@�K����!?"Ym4��@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@E�2U>�ٿ����5��@(�7)�4@{Ǥ0s�!?���&�@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@Ȯ؃c�ٿ�W�{��@k(Gb�4@�|����!?���a��@,���ʉٿ���n��@�1�4@������!?�}��@,���ʉٿ���n��@�1�4@������!?�}��@,���ʉٿ���n��@�1�4@������!?�}��@,���ʉٿ���n��@�1�4@������!?�}��@����ٿ�cg���@|���4@#�}ƪ�!?\����@����ٿ�cg���@|���4@#�}ƪ�!?\����@����ٿ�cg���@|���4@#�}ƪ�!?\����@����ٿ�cg���@|���4@#�}ƪ�!?\����@����ٿ�cg���@|���4@#�}ƪ�!?\����@k��jq�ٿ�7���@�q��4@?�hT��!?���J�@k��jq�ٿ�7���@�q��4@?�hT��!?���J�@k��jq�ٿ�7���@�q��4@?�hT��!?���J�@k��jq�ٿ�7���@�q��4@?�hT��!?���J�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@/�^�a�ٿ�|k����@@�S�4@��s�!?h>�,+_�@ƀ��ٿ������@���L4@� l蝐!?@�2�l��@ƀ��ٿ������@���L4@� l蝐!?@�2�l��@ƀ��ٿ������@���L4@� l蝐!?@�2�l��@ƀ��ٿ������@���L4@� l蝐!?@�2�l��@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@������ٿ}��y2�@�#	�B4@�dv��!?���@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@�ۖ��ٿ7�	a��@�l�j� 4@
�^��!?�������@3_Z�ٿ�6QK
�@���� 4@3��0�!?������@3_Z�ٿ�6QK
�@���� 4@3��0�!?������@�ٛ�-|ٿ�՗���@\$���4@b��&��!?�f���@�ٛ�-|ٿ�՗���@\$���4@b��&��!?�f���@�ٛ�-|ٿ�՗���@\$���4@b��&��!?�f���@��!��|ٿ� nJs��@�+�04@p{F�~�!?�>@����@��!��|ٿ� nJs��@�+�04@p{F�~�!?�>@����@��!��|ٿ� nJs��@�+�04@p{F�~�!?�>@����@��o=��ٿݛ8?�;�@N��4@��;Iѐ!?h���>u�@��o=��ٿݛ8?�;�@N��4@��;Iѐ!?h���>u�@��o=��ٿݛ8?�;�@N��4@��;Iѐ!?h���>u�@��o=��ٿݛ8?�;�@N��4@��;Iѐ!?h���>u�@��o=��ٿݛ8?�;�@N��4@��;Iѐ!?h���>u�@����܊ٿ�,>5F�@��M]4@�YkIT�!?����2�@����܊ٿ�,>5F�@��M]4@�YkIT�!?����2�@����܊ٿ�,>5F�@��M]4@�YkIT�!?����2�@�<�F؋ٿ�Џ��;�@��#��4@���h�!?��`�
�@�<�F؋ٿ�Џ��;�@��#��4@���h�!?��`�
�@�<�F؋ٿ�Џ��;�@��#��4@���h�!?��`�
�@�<�F؋ٿ�Џ��;�@��#��4@���h�!?��`�
�@�<�F؋ٿ�Џ��;�@��#��4@���h�!?��`�
�@��ٿ�FҜ�2�@oP�4@v���!?VR����@��ٿ�FҜ�2�@oP�4@v���!?VR����@��ٿ�FҜ�2�@oP�4@v���!?VR����@��ٿ�FҜ�2�@oP�4@v���!?VR����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�촷��ٿE{��w�@}�V��4@ՙ�!?P����@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@�Bҙ��ٿ�w��H^�@Ϛꥴ4@����!?S�C_���@����}ٿjí�z�@�I�u4@�V�1�!?@����w�@�S�ktyٿ%�j;l��@�_�U>4@���]D�!?|��M8<�@�S�ktyٿ%�j;l��@�_�U>4@���]D�!?|��M8<�@�S�ktyٿ%�j;l��@�_�U>4@���]D�!?|��M8<�@^8��R�ٿ�H6 .Z�@b�_�F4@>`D�Ɛ!?�u-	ɓ�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��cXǀٿja��6�@D�+b4@g_O���!?*��jr
�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@��D��~ٿ5�MI���@���Ի4@Vx�Ő!?��ج6]�@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@.;fٿMɼ+���@�Rbc4@/�w�!?�������@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@�h:'��ٿV�`ՠY�@Eɻ�	4@H����!?%��x���@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@={R�ٿ8x��>��@t�o��4@*X$vߐ!?&��w�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�C��ٿK�`���@{�4@�[��ڐ!?��G��h�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�{��Ąٿ~Ʉ���@���334@&9[e��!?�5�ǁ�@�v�  �ٿ���H��@�ȘT4@��xĳ�!?�V�I�(�@�v�  �ٿ���H��@�ȘT4@��xĳ�!?�V�I�(�@�X��{�ٿ�v��L�@��a4@рGW��!?X������@�����ٿ�y����@���B4@i��jv�!?���u�@N���N�ٿe���B��@�#�w4@�m��!?��v+��@N���N�ٿe���B��@�#�w4@�m��!?��v+��@N���N�ٿe���B��@�#�w4@�m��!?��v+��@N���N�ٿe���B��@�#�w4@�m��!?��v+��@N���N�ٿe���B��@�#�w4@�m��!?��v+��@���dV�ٿ|؞��E�@�m�( 4@��c�!?Vf�9�,�@\J���ٿ5�,�z��@ ��G4@@��!?��d\�@\J���ٿ5�,�z��@ ��G4@@��!?��d\�@\J���ٿ5�,�z��@ ��G4@@��!?��d\�@\J���ٿ5�,�z��@ ��G4@@��!?��d\�@\J���ٿ5�,�z��@ ��G4@@��!?��d\�@
���ٿ!�ķCY�@���4@��f�!?�O���,�@�8�]�ٿJ1�8���@30X4@uE��!?A2^�e��@�'� +�ٿ�Ȧ���@�)��4@Ʀ�fE�!?8��u���@�'� +�ٿ�Ȧ���@�)��4@Ʀ�fE�!?8��u���@�'� +�ٿ�Ȧ���@�)��4@Ʀ�fE�!?8��u���@�L-C�}ٿ�U����@ͨ*%4@��!?��Q����@lu ��~ٿGV�{�e�@1��4@$5�}Đ!?2��p��@lu ��~ٿGV�{�e�@1��4@$5�}Đ!?2��p��@lu ��~ٿGV�{�e�@1��4@$5�}Đ!?2��p��@P�=�ٿ�����@��?�4@R���ǐ!?%�m�r�@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���s�ٿ���!��@�Mߓ4@Rίn��!?�)Ю��@���F~ٿ��8���@�,�@�	4@Ȓ���!?8x�U��@���F~ٿ��8���@�,�@�	4@Ȓ���!?8x�U��@�E�KٿY��4���@�\�B�4@
��9g�!?��R-\��@�E�KٿY��4���@�\�B�4@
��9g�!?��R-\��@�E�KٿY��4���@�\�B�4@
��9g�!?��R-\��@�E�KٿY��4���@�\�B�4@
��9g�!?��R-\��@�H��ٿJ�!_Ee�@d�u�4@���!?K��I<��@�H��ٿJ�!_Ee�@d�u�4@���!?K��I<��@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@Rɝ3F�ٿ��J�@�2�U4@e�謐!?X}_��C�@�*��s�ٿ◙:Gw�@�,2ed4@�D
��!?�vv�^�@�*��s�ٿ◙:Gw�@�,2ed4@�D
��!?�vv�^�@�*��s�ٿ◙:Gw�@�,2ed4@�D
��!?�vv�^�@6[�xU�ٿ��RI���@�b�d4@��y�Ӑ!?#K�^9�@6[�xU�ٿ��RI���@�b�d4@��y�Ӑ!?#K�^9�@6[�xU�ٿ��RI���@�b�d4@��y�Ӑ!?#K�^9�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@$1�r�ٿ}$����@�\��4@�}t�Ԑ!?hWa[�@�6�y�ٿl&9���@����4@���k��!?�8�|�@�6�y�ٿl&9���@����4@���k��!?�8�|�@�6�y�ٿl&9���@����4@���k��!?�8�|�@�6�y�ٿl&9���@����4@���k��!?�8�|�@�6�y�ٿl&9���@����4@���k��!?�8�|�@�6�y�ٿl&9���@����4@���k��!?�8�|�@ �A��ٿ�Z)-�U�@��N���3@#Z�S��!?������@ �A��ٿ�Z)-�U�@��N���3@#Z�S��!?������@Y�����ٿ9)���@py����3@�#�q��!?�դ� �@Y�����ٿ9)���@py����3@�#�q��!?�դ� �@Y�����ٿ9)���@py����3@�#�q��!?�դ� �@��$׈ٿ�!���)�@`�����3@ �q��!?$&���@��$׈ٿ�!���)�@`�����3@ �q��!?$&���@��$׈ٿ�!���)�@`�����3@ �q��!?$&���@��$׈ٿ�!���)�@`�����3@ �q��!?$&���@��$׈ٿ�!���)�@`�����3@ �q��!?$&���@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@�^�ٿK�}Y�@���d�4@��GR[�!?}$�3�r�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��X�܆ٿP��7���@�e��4@"n����!?�R��n�@��i���ٿ�!���@��J4@yL���!?�خ�o�@3@��ٿ��#���@l��;]4@"5m� �!?=X��"�@3@��ٿ��#���@l��;]4@"5m� �!?=X��"�@3@��ٿ��#���@l��;]4@"5m� �!?=X��"�@��|���ٿ�}ÉV��@�q�S04@�l����!?6i�(s��@��|���ٿ�}ÉV��@�q�S04@�l����!?6i�(s��@��|���ٿ�}ÉV��@�q�S04@�l����!?6i�(s��@�tQ�l�ٿ�F���	�@nC��i4@��	��!?dk�{H�@�tQ�l�ٿ�F���	�@nC��i4@��	��!?dk�{H�@��_�ٿ��TL�@���~�4@�R�[Ґ!?]�}\-�@��_�ٿ��TL�@���~�4@�R�[Ґ!?]�}\-�@��_�ٿ��TL�@���~�4@�R�[Ґ!?]�}\-�@Ԭu�~ٿ�n4�j��@(���4@�"@��!?TV�|�.�@Ԭu�~ٿ�n4�j��@(���4@�"@��!?TV�|�.�@Ԭu�~ٿ�n4�j��@(���4@�"@��!?TV�|�.�@�dk�S�ٿo N.���@���/c4@��+ΐ!?�*m*��@�dk�S�ٿo N.���@���/c4@��+ΐ!?�*m*��@T�N�ٿ��?�F�@O�Ȅ4@×�\�!?rX糊��@T�N�ٿ��?�F�@O�Ȅ4@×�\�!?rX糊��@T�N�ٿ��?�F�@O�Ȅ4@×�\�!?rX糊��@T�N�ٿ��?�F�@O�Ȅ4@×�\�!?rX糊��@T�N�ٿ��?�F�@O�Ȅ4@×�\�!?rX糊��@�R6�T�ٿ��"L�@�	8��4@X��?�!?y��=��@����ٿ��ʴF��@�r�4z4@��e��!?4= ����@��هٿ��[EvA�@���+�4@�S|<��!?��I����@��هٿ��[EvA�@���+�4@�S|<��!?��I����@��هٿ��[EvA�@���+�4@�S|<��!?��I����@��هٿ��[EvA�@���+�4@�S|<��!?��I����@l���ٿ?@�b�@���eg4@�L�:��!?�8�dg�@l���ٿ?@�b�@���eg4@�L�:��!?�8�dg�@l���ٿ?@�b�@���eg4@�L�:��!?�8�dg�@�s��ٿ�
0Mc�@��6,�4@M
�ϐ!?�a���@�s��ٿ�
0Mc�@��6,�4@M
�ϐ!?�a���@T���O�ٿ�`���@�x�ӈ 4@��rt�!?��*-b�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@��+��ٿ�)i�L9�@?�}� 4@#q4��!?�҄9'9�@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@KfF�ʆٿ� ݚ<G�@����4@j
���!?+�|8W��@/�CCQ�ٿ�L}����@��t(q4@�+[���!?U2���@/�CCQ�ٿ�L}����@��t(q4@�+[���!?U2���@/�CCQ�ٿ�L}����@��t(q4@�+[���!?U2���@IƢ�{ٿAS��TS�@Άԯ4@����ǐ!?P�����@IƢ�{ٿAS��TS�@Άԯ4@����ǐ!?P�����@�9qh�ٿ=ۃSc��@yL<qi4@έ����!?ߵ0��\�@�9qh�ٿ=ۃSc��@yL<qi4@έ����!?ߵ0��\�@�9qh�ٿ=ۃSc��@yL<qi4@έ����!?ߵ0��\�@�9qh�ٿ=ۃSc��@yL<qi4@έ����!?ߵ0��\�@�9qh�ٿ=ۃSc��@yL<qi4@έ����!?ߵ0��\�@�\k�ފٿ\Ku�5�@��T:4@�Iet�!?�C/��@�J��n�ٿ�1���C�@9v�4@sKm��!?�k�X0�@�5��ؔٿ���9���@�F�z4@�/���!?�r�!7�@�5��ؔٿ���9���@�F�z4@�/���!?�r�!7�@�5��ؔٿ���9���@�F�z4@�/���!?�r�!7�@�,(�ٿF�ޣ+��@����
4@(�Xj��!?+�t�]��@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@I^��ٿ�|����@}��u94@� �sא!?�j2��I�@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@y�w��ٿ�'�\��@L���4@A�8ʔ�!?��#(���@A��ײ�ٿ���"��@��24@|��!?"p��N��@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�m䧉ٿ��v8��@���4@�Ţ�!�!?Q��~�@�LF��ٿ���v��@]����4@�^\9��!?H�wH��@�LF��ٿ���v��@]����4@�^\9��!?H�wH��@�LF��ٿ���v��@]����4@�^\9��!?H�wH��@�LF��ٿ���v��@]����4@�^\9��!?H�wH��@ӫ���ٿ�M,)h�@��F"m4@$��/��!?���L���@�u�Ԏٿn��sU�@�>��4@୩ʐ!?�\\����@���"�ٿ��\�t��@g�7�4@���i�!?;����8�@���"�ٿ��\�t��@g�7�4@���i�!?;����8�@8����ٿy���$��@���"�4@�3|pŐ!?�t����@���Ќٿ@1\=�@s�=b4@��8���!?��2�U�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�2�F��ٿ?!y����@5U�~a4@��݃��!?Pù��t�@�!���ٿX93n��@E!?��4@���ǹ�!?����5�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�,@	�ٿ�;r*�@��Q 4@�W��!?�g��!�@�N���ٿ�ڽW��@S�F2�4@���2̐!?G	�H��@��xE<�ٿ�Ly��@�g��4@�@�q�!?�L\ ��@X:6�ٿֈø4 �@]���4@�8;_
�!?V�$,z��@X:6�ٿֈø4 �@]���4@�8;_
�!?V�$,z��@C/r��ٿ�6_t���@�(A4@#�`ΐ!?�b��@C/r��ٿ�6_t���@�(A4@#�`ΐ!?�b��@C/r��ٿ�6_t���@�(A4@#�`ΐ!?�b��@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@N ��f�ٿd���	I�@{��0K4@Rv�Ր!?��P���@��8�ٿ�"��`�@`��m4@�<G�!?[����R�@P �@�ٿGl̷��@�AX4@�ht���!?�|���@P �@�ٿGl̷��@�AX4@�ht���!?�|���@P �@�ٿGl̷��@�AX4@�ht���!?�|���@P �@�ٿGl̷��@�AX4@�ht���!?�|���@P �@�ٿGl̷��@�AX4@�ht���!?�|���@P �@�ٿGl̷��@�AX4@�ht���!?�|���@C���/�ٿ�{����@2�ؙ�4@Yhd���!? ���.1�@C���/�ٿ�{����@2�ؙ�4@Yhd���!? ���.1�@_�ľ9�ٿl�U�xs�@W�|�4@Tʹv�!?y@2����@_�ľ9�ٿl�U�xs�@W�|�4@Tʹv�!?y@2����@�T,�Ƅٿא���1�@Xb�G4@M��k�!?������@�T,�Ƅٿא���1�@Xb�G4@M��k�!?������@�T,�Ƅٿא���1�@Xb�G4@M��k�!?������@�T,�Ƅٿא���1�@Xb�G4@M��k�!?������@�T,�Ƅٿא���1�@Xb�G4@M��k�!?������@?i͗m�ٿ8����@���4@�\+/l�!?,����Q�@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@T�WF�ٿ-�ϳ��@]�un�4@u���!?������@U�h�9�ٿ��CM��@+F� g4@�sj
��!?[�Lp��@U�h�9�ٿ��CM��@+F� g4@�sj
��!?[�Lp��@U�h�9�ٿ��CM��@+F� g4@�sj
��!?[�Lp��@RvL>݀ٿ-�\�Bo�@�aQ�4@Bzw�!?�e����@RvL>݀ٿ-�\�Bo�@�aQ�4@Bzw�!?�e����@RvL>݀ٿ-�\�Bo�@�aQ�4@Bzw�!?�e����@RvL>݀ٿ-�\�Bo�@�aQ�4@Bzw�!?�e����@o_�v%~ٿ����m�@.׎�4@�i����!?i�,�с�@o_�v%~ٿ����m�@.׎�4@�i����!?i�,�с�@�$,[h~ٿ�XXJ�@��Z=?4@�QkRא!?&E�`�X�@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@URȌ��ٿC��#�@�:�:e4@������!?�n����@��8āٿiZB��A�@��Qo�4@/{)̊�!?��IJ���@]*|�ٿ�2V9T��@<��{4@���֐!?L��қr�@]*|�ٿ�2V9T��@<��{4@���֐!?L��қr�@��g0^�ٿJ���_�@�Ґ�4@y�~?�!?gro0��@��g0^�ٿJ���_�@�Ґ�4@y�~?�!?gro0��@��g0^�ٿJ���_�@�Ґ�4@y�~?�!?gro0��@nj+=ƊٿZ�� ͐�@0(��U4@կɎ��!?᧞�I�@nj+=ƊٿZ�� ͐�@0(��U4@կɎ��!?᧞�I�@nj+=ƊٿZ�� ͐�@0(��U4@կɎ��!?᧞�I�@��+3�ٿ�³?\�@?��t4@�?��)�!?Q�� +y�@�NY9X|ٿk@�7��@��4@����!?�M<����@��a'�ٿ�gE��@Kp�.4@�b�t��!?�Xb�8�@��a'�ٿ�gE��@Kp�.4@�b�t��!?�Xb�8�@��a'�ٿ�gE��@Kp�.4@�b�t��!?�Xb�8�@��a'�ٿ�gE��@Kp�.4@�b�t��!?�Xb�8�@%��{�ٿ�*e�(Q�@���G�4@��CQ*�!?��= v�@%��{�ٿ�*e�(Q�@���G�4@��CQ*�!?��= v�@%��{�ٿ�*e�(Q�@���G�4@��CQ*�!?��= v�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@_���!�ٿ��#G��@����]�3@Zb	�!?�N?>YJ�@�sDT~ٿSU�AY�@X7���4@�T���!?W����:�@�sDT~ٿSU�AY�@X7���4@�T���!?W����:�@�sDT~ٿSU�AY�@X7���4@�T���!?W����:�@�sDT~ٿSU�AY�@X7���4@�T���!?W����:�@8Kf�"�ٿ,�_(&��@<���	4@"n�4�!?� :�;P�@8Kf�"�ٿ,�_(&��@<���	4@"n�4�!?� :�;P�@[4���ٿQ"+�f�@1��4@8&v�!?�K)���@[4���ٿQ"+�f�@1��4@8&v�!?�K)���@[4���ٿQ"+�f�@1��4@8&v�!?�K)���@[4���ٿQ"+�f�@1��4@8&v�!?�K)���@[4���ٿQ"+�f�@1��4@8&v�!?�K)���@S~���ٿ-�Y�@e��w� 4@�xox�!?��Q5W�@S~���ٿ-�Y�@e��w� 4@�xox�!?��Q5W�@S~���ٿ-�Y�@e��w� 4@�xox�!?��Q5W�@O ����ٿQ�[hJ�@h�2��4@��(��!?A�=���@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@Qdu�܍ٿV�5����@?�)G�4@}"�2ߐ!?�K"�w�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@@g͆ٿ^�_]�B�@I����4@5�u+��!?f��k�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@�`G�ٿ�c��^�@�.�g�4@�gW�Đ!?ýx �;�@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@xp���ٿ2������@��ӆ�4@�og���!?���\���@���Q�ٿ���Mu�@���(4@A�%,��!?�M�����@���Q�ٿ���Mu�@���(4@A�%,��!?�M�����@���Q�ٿ���Mu�@���(4@A�%,��!?�M�����@�ЦI`�ٿcK&�N�@��́4@�ۓ��!?&<����@�ЦI`�ٿcK&�N�@��́4@�ۓ��!?&<����@�ЦI`�ٿcK&�N�@��́4@�ۓ��!?&<����@�ЦI`�ٿcK&�N�@��́4@�ۓ��!?&<����@V�(�G�ٿ����m�@���4@ �L��!?����"i�@�o�L�ٿ[X���@���#�4@b,�P|�!?�ܶ)́�@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@��،�ٿ4���-�@����T4@9�ξ�!?�2M�K��@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@z���O�ٿ@���@���04@.W枱�!?��tc;Z�@�?�ϳ�ٿGBQ��@zA��4@\��aѐ!?���Pt�@�WM�j�ٿ���ë��@�`��4@��&��!?.�8���@��I�ނٿ����A�@�Vpx4@���	�!?�*�9�U�@��I�ނٿ����A�@�Vpx4@���	�!?�*�9�U�@��I�ނٿ����A�@�Vpx4@���	�!?�*�9�U�@^2ZIl�ٿ!���Ya�@m���4@ɓ�颐!?�'��j��@^2ZIl�ٿ!���Ya�@m���4@ɓ�颐!?�'��j��@^2ZIl�ٿ!���Ya�@m���4@ɓ�颐!?�'��j��@^2ZIl�ٿ!���Ya�@m���4@ɓ�颐!?�'��j��@�o��H�ٿu���I�@�@k4@�����!?iR�_��@�o��H�ٿu���I�@�@k4@�����!?iR�_��@�o��H�ٿu���I�@�@k4@�����!?iR�_��@�o��H�ٿu���I�@�@k4@�����!?iR�_��@7��
L�ٿ7ѡ/h/�@��r�4@,ʵ�!?-�	A�@7��
L�ٿ7ѡ/h/�@��r�4@,ʵ�!?-�	A�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@Ҫ��$�ٿ5
�ie��@'s�HY4@	��F��!?*HIxc�@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@%mK<��ٿE-͢���@�-�J�4@S��G�!?��P~��@�3܎�ٿ�.T�ԝ�@��{d�4@����V�!? �WA�P�@ζ�K�ٿ�W�j��@L����
4@��w���!? ��o�@ζ�K�ٿ�W�j��@L����
4@��w���!? ��o�@ζ�K�ٿ�W�j��@L����
4@��w���!? ��o�@ζ�K�ٿ�W�j��@L����
4@��w���!? ��o�@ΰ@�l�ٿwP�[���@&�Ǿ	4@���+��!?$�9��f�@ΰ@�l�ٿwP�[���@&�Ǿ	4@���+��!?$�9��f�@ΰ@�l�ٿwP�[���@&�Ǿ	4@���+��!?$�9��f�@�����ٿ��Ţ@�@	4@%�j��!?����R�@�����ٿ��Ţ@�@	4@%�j��!?����R�@�����ٿ��Ţ@�@	4@%�j��!?����R�@�����ٿ��Ţ@�@	4@%�j��!?����R�@�V����ٿhH�l��@����4@��!?0|�j��@�V����ٿhH�l��@����4@��!?0|�j��@V�.˩�ٿn��'�@iߍ�n4@&}���!?��U�mZ�@V�.˩�ٿn��'�@iߍ�n4@&}���!?��U�mZ�@��;�ٿ�a�f6�@͠�1�4@�G���!?R��̚�@�u�x�ٿ��'K�(�@j�D�4@q;�tڐ!?]������@�u�x�ٿ��'K�(�@j�D�4@q;�tڐ!?]������@�u�x�ٿ��'K�(�@j�D�4@q;�tڐ!?]������@�u�x�ٿ��'K�(�@j�D�4@q;�tڐ!?]������@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@^�ѵ!�ٿ�ew���@n��.o4@(�<�W�!?�X2J�_�@.ݥxÈٿw�����@u��! 4@���yƐ!?������@>II��ٿ8Y^h2>�@.uv��3@Ȯ{�!?������@>II��ٿ8Y^h2>�@.uv��3@Ȯ{�!?������@>II��ٿ8Y^h2>�@.uv��3@Ȯ{�!?������@�*�(��ٿ�n'+c��@�����4@�.~� �!?�hey�#�@�*�(��ٿ�n'+c��@�����4@�.~� �!?�hey�#�@�*�(��ٿ�n'+c��@�����4@�.~� �!?�hey�#�@��K���ٿГ�Zo�@'q�L�3@�{�'&�!?SG�Pn��@��K���ٿГ�Zo�@'q�L�3@�{�'&�!?SG�Pn��@��K���ٿГ�Zo�@'q�L�3@�{�'&�!?SG�Pn��@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�״��ٿ/��R��@���=�3@$oi71�!?(P����@�X���ٿx챑�^�@(ll��4@�Rf/H�!?��P�@�X���ٿx챑�^�@(ll��4@�Rf/H�!?��P�@�X���ٿx챑�^�@(ll��4@�Rf/H�!?��P�@�X���ٿx챑�^�@(ll��4@�Rf/H�!?��P�@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@A�kim�ٿ� ܯ�@8`�4@	��0b�!?�c����@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@3I�8D�ٿ�{v	��@��[u�4@X<��!?<ڍ�!��@\G���ٿ��[W>�@�qTذ4@=���!?G2�?V�@\G���ٿ��[W>�@�qTذ4@=���!?G2�?V�@\G���ٿ��[W>�@�qTذ4@=���!?G2�?V�@\G���ٿ��[W>�@�qTذ4@=���!?G2�?V�@������ٿQ�+��@9IhTW4@��tq��!?�᩶!��@������ٿQ�+��@9IhTW4@��tq��!?�᩶!��@������ٿQ�+��@9IhTW4@��tq��!?�᩶!��@������ٿQ�+��@9IhTW4@��tq��!?�᩶!��@�,[�o�ٿ�~����@��u�4@c�nJ�!?V�ߑ$F�@�,[�o�ٿ�~����@��u�4@c�nJ�!?V�ߑ$F�@�,[�o�ٿ�~����@��u�4@c�nJ�!?V�ߑ$F�@�,[�o�ٿ�~����@��u�4@c�nJ�!?V�ߑ$F�@=��a�ٿ����S�@&��4@V��2$�!?j�j�b��@=��a�ٿ����S�@&��4@V��2$�!?j�j�b��@�V+aw�ٿ�s�T�U�@d�
��4@���1�!?:
��)�@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@S��}�ٿ3��t>�@k%��84@�ڠ�}�!?0@�
i��@�cz�ٿ�_���@Q�Bi�	4@B�mV͐!?����L�@�cz�ٿ�_���@Q�Bi�	4@B�mV͐!?����L�@�cz�ٿ�_���@Q�Bi�	4@B�mV͐!?����L�@�cz�ٿ�_���@Q�Bi�	4@B�mV͐!?����L�@�cz�ٿ�_���@Q�Bi�	4@B�mV͐!?����L�@`2 ��ٿ�ILjeh�@����3@oķ�!?����@`2 ��ٿ�ILjeh�@����3@oķ�!?����@`2 ��ٿ�ILjeh�@����3@oķ�!?����@`2 ��ٿ�ILjeh�@����3@oķ�!?����@�X����ٿ���U9S�@Is��4@G�kX��!?UV�)��@�X����ٿ���U9S�@Is��4@G�kX��!?UV�)��@�X����ٿ���U9S�@Is��4@G�kX��!?UV�)��@@�V�ٿx�sx��@����.4@6�7�ɐ!?j�oq���@^xp"z�ٿY?����@��o�4@u?�+��!?ȁ��U�@^xp"z�ٿY?����@��o�4@u?�+��!?ȁ��U�@^xp"z�ٿY?����@��o�4@u?�+��!?ȁ��U�@��B�s�ٿ$���F�@L��4@�usjO�!?�ݩ1���@��B�s�ٿ$���F�@L��4@�usjO�!?�ݩ1���@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@T��^yٿ@�[,�@��=LW4@OkӐ!?y�j��@�d��~ٿ?S����@ld&�4@8�,B�!?;�{L��@�d��~ٿ?S����@ld&�4@8�,B�!?;�{L��@z�,���ٿ �P`�@�.�n4@Ha�Gs�!?��0���@z�,���ٿ �P`�@�.�n4@Ha�Gs�!?��0���@z�,���ٿ �P`�@�.�n4@Ha�Gs�!?��0���@z�,���ٿ �P`�@�.�n4@Ha�Gs�!?��0���@z�,���ٿ �P`�@�.�n4@Ha�Gs�!?��0���@�ee�#{ٿn����@�� N_4@� �ې!?���KN�@�ee�#{ٿn����@�� N_4@� �ې!?���KN�@��m܁ٿ�F�#0�@jD�U4@ň|�!?��A�¬�@��m܁ٿ�F�#0�@jD�U4@ň|�!?��A�¬�@��m܁ٿ�F�#0�@jD�U4@ň|�!?��A�¬�@��m܁ٿ�F�#0�@jD�U4@ň|�!?��A�¬�@��m܁ٿ�F�#0�@jD�U4@ň|�!?��A�¬�@����[�ٿ�)�XT��@�z|{I4@�����!?:\2ʄ]�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@��Z��ٿ��f����@5�E-t	4@��~v��!?�Z�;"�@B\��ٿ�s�����@k����4@2�'Ɛ!?-������@B\��ٿ�s�����@k����4@2�'Ɛ!?-������@B\��ٿ�s�����@k����4@2�'Ɛ!?-������@B\��ٿ�s�����@k����4@2�'Ɛ!?-������@B\��ٿ�s�����@k����4@2�'Ɛ!?-������@�=���ٿ Ѡo��@;���A4@���T�!?��Q]���@i��ٿ��ce�@K�;�
4@=�xӐ!?zՒlO�@i��ٿ��ce�@K�;�
4@=�xӐ!?zՒlO�@i��ٿ��ce�@K�;�
4@=�xӐ!?zՒlO�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@��ٿ6t� � �@E��	4@�I�l��!?�++ua�@�.ܓ��ٿ�a��n��@����4@�aÞ��!?p�W���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@ک ��ٿ/�ч��@w�z�O4@s�D�!?�Ӎ���@�R��ٿ�T��_��@�E)�{4@%�����!?�&(t�@�R��ٿ�T��_��@�E)�{4@%�����!?�&(t�@�R��ٿ�T��_��@�E)�{4@%�����!?�&(t�@�R��ٿ�T��_��@�E)�{4@%�����!?�&(t�@�R��ٿ�T��_��@�E)�{4@%�����!?�&(t�@Hx��ٿ�k�po^�@�o�4@�v�ސ!?�n�{\��@]f~��ٿ
��_u��@�ږ��4@-QE���!?����G�@]f~��ٿ
��_u��@�ږ��4@-QE���!?����G�@]f~��ٿ
��_u��@�ږ��4@-QE���!?����G�@]f~��ٿ
��_u��@�ږ��4@-QE���!?����G�@]f~��ٿ
��_u��@�ږ��4@-QE���!?����G�@�%pz �ٿ��EV"2�@n�4@l����!? �8�s5�@�%pz �ٿ��EV"2�@n�4@l����!? �8�s5�@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@x�0�ٿ�a��@_*��4@ƭ5�А!??>ȥJ��@pIv��ٿe@U�H��@b_ҋ4@����֐!?:��EÑ�@pIv��ٿe@U�H��@b_ҋ4@����֐!?:��EÑ�@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�z"NÄٿB%��t��@F�~� 4@�]�Dڐ!?��c~b��@�1����ٿ��f�9�@��R�� 4@0	��!?��ڹ���@�1����ٿ��f�9�@��R�� 4@0	��!?��ڹ���@"���ٿúi,���@�7�Q'4@c�1t��!?�mw���@"���ٿúi,���@�7�Q'4@c�1t��!?�mw���@"���ٿúi,���@�7�Q'4@c�1t��!?�mw���@"���ٿúi,���@�7�Q'4@c�1t��!?�mw���@>U�f9�ٿ��!�@�}A�4@�+�Ő!?X(���@>U�f9�ٿ��!�@�}A�4@�+�Ő!?X(���@>U�f9�ٿ��!�@�}A�4@�+�Ő!?X(���@]:'�Ňٿ����.	�@Tb�� 4@��w�ɐ!?��O�M��@�	}�h�ٿ����"�@ͥ�t 4@�'0���!?����+�@�	}�h�ٿ����"�@ͥ�t 4@�'0���!?����+�@߂�	�ٿc�Y&�@��:ǐ4@;rW��!?���i��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@ץv�ٿ���6�@)�(�4@���ǐ!?�>�c��@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��õ��ٿj�D���@9���o4@K��ܐ!?��u�I�@��-;݆ٿ�LKi���@b<獥4@Lq�)�!?`�r��@��-;݆ٿ�LKi���@b<獥4@Lq�)�!?`�r��@��-;݆ٿ�LKi���@b<獥4@Lq�)�!?`�r��@��^��ٿ�"#�%�@��@6� 4@��ȥ�!?�k@�x��@��^��ٿ�"#�%�@��@6� 4@��ȥ�!?�k@�x��@��^��ٿ�"#�%�@��@6� 4@��ȥ�!?�k@�x��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@�M��(�ٿ��=��@�����4@����!?Z  ��@5)����ٿB��@�mK�4@�~��%�!? ����@5)����ٿB��@�mK�4@�~��%�!? ����@5)����ٿB��@�mK�4@�~��%�!? ����@5)����ٿB��@�mK�4@�~��%�!? ����@5)����ٿB��@�mK�4@�~��%�!? ����@5)����ٿB��@�mK�4@�~��%�!? ����@��Zv��ٿL �߮X�@�*�u� 4@<�E*,�!?�;�.���@r&+�5�ٿh٬��@�K|��4@��5�)�!?2�����@�ä8U�ٿ�a$�@��xd4@�j���!?ˊ�
i��@��8���ٿ3��m*�@�О4@������!?�>����@��8���ٿ3��m*�@�О4@������!?�>����@��8���ٿ3��m*�@�О4@������!?�>����@��Q�|ٿ��
���@岒�4@�����!?�X����@��Q�|ٿ��
���@岒�4@�����!?�X����@��Q�|ٿ��
���@岒�4@�����!?�X����@��Q�|ٿ��
���@岒�4@�����!?�X����@��Q�|ٿ��
���@岒�4@�����!?�X����@��Q�|ٿ��
���@岒�4@�����!?�X����@8'`�F�ٿ�%=��@ 	9�1�3@\Ѵ���!?����x��@	��d�ٿoImr���@��I��3@A��*v�!?!Qv����@��o��ٿ�)?W�"�@;�U��3@�}����!?���Y�@��o��ٿ�)?W�"�@;�U��3@�}����!?���Y�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�ZE_&�ٿ���4��@r�BH�4@�y���!?�(,V,Z�@�����ٿJ<|_A��@�[Zo,4@���a�!?Ak	A��@�����ٿJ<|_A��@�[Zo,4@���a�!?Ak	A��@�����ٿJ<|_A��@�[Zo,4@���a�!?Ak	A��@�����ٿJ<|_A��@�[Zo,4@���a�!?Ak	A��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@��΄�ٿ�4����@��dmN4@�~��!?�ҌY��@z���|�ٿ�e�A?��@1і��4@3Ϣ?ݐ!?J�����@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@��*��ٿ�h����@��C�4@�n���!?�M���@�@0�?��ٿ
���w�@*A\�4@g���!?�SL��@�8Ϻ�ٿ���^+��@��4@���ܦ�!?�/����@�8Ϻ�ٿ���^+��@��4@���ܦ�!?�/����@��e[ �ٿ�����@,E�ڿ4@!aA/Ɛ!?�D�b��@wR>Xd�ٿ2ר��@�ξB4@ ����!?�㊾���@wR>Xd�ٿ2ר��@�ξB4@ ����!?�㊾���@wR>Xd�ٿ2ר��@�ξB4@ ����!?�㊾���@wR>Xd�ٿ2ר��@�ξB4@ ����!?�㊾���@wR>Xd�ٿ2ר��@�ξB4@ ����!?�㊾���@�{�Մ�ٿd4�����@ŉ��
4@����ڐ!?�\\��@�����ٿ`�#�M"�@/[O64@F�py�!?�`W��@�����ٿ`�#�M"�@/[O64@F�py�!?�`W��@�����ٿ`�#�M"�@/[O64@F�py�!?�`W��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�{/�ٿU�ua)#�@��4@m�6Ő!?Eqk�,��@�|��ٿB�Gѣ�@��Z��4@-�{���!?N�~�@�|��ٿB�Gѣ�@��Z��4@-�{���!?N�~�@�|��ٿB�Gѣ�@��Z��4@-�{���!?N�~�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@~t'��ٿ�u���@�`���4@d����!?0P�.�@��ѓ�ٿԷ�ŝ6�@�Z]�4@�0}͐!?Ur[��@`��ٿ1MVYV)�@ҰZ�4@E�'��!?/��b�@�,�/ٿ���!�@�>7�4@�[�Ր!?��g�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@�����ٿkw�s�9�@k�	��4@�0k�!?��3�[�@+���g�ٿ�����@b�U�64@�����!?ʤ�?<w�@+���g�ٿ�����@b�U�64@�����!?ʤ�?<w�@�����|ٿ�uċ���@���4@�C��!?��g9h�@�����|ٿ�uċ���@���4@�C��!?��g9h�@�����|ٿ�uċ���@���4@�C��!?��g9h�@�����|ٿ�uċ���@���4@�C��!?��g9h�@�_��j{ٿL�����@쨔�4@�W��!?q1�3}�@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@X32�~ٿ��^Z��@xM�4@��*���!?��y��@�6�g��ٿ�R��j��@[�_H;4@U+�l�!?���M׫�@�6�g��ٿ�R��j��@[�_H;4@U+�l�!?���M׫�@�6�g��ٿ�R��j��@[�_H;4@U+�l�!?���M׫�@�6�g��ٿ�R��j��@[�_H;4@U+�l�!?���M׫�@�6�g��ٿ�R��j��@[�_H;4@U+�l�!?���M׫�@=J+<H�ٿ�@V!Y}�@��e\4@>�nJ��!?���`��@=J+<H�ٿ�@V!Y}�@��e\4@>�nJ��!?���`��@=J+<H�ٿ�@V!Y}�@��e\4@>�nJ��!?���`��@"��_�ٿ�*j,��@���C�4@�x�^��!?�y�e:`�@�'��ٿ-C@�r�@$��&4@`ީx�!?��)ҽ�@���b�ٿ��Lֹ�@��/��4@�!N�!?�FlZ�_�@���b�ٿ��Lֹ�@��/��4@�!N�!?�FlZ�_�@���b�ٿ��Lֹ�@��/��4@�!N�!?�FlZ�_�@���b�ٿ��Lֹ�@��/��4@�!N�!?�FlZ�_�@���b�ٿ��Lֹ�@��/��4@�!N�!?�FlZ�_�@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@Ǳo�5�ٿ�N���@����4@D��9��!?3��r��@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@dA$資ٿ��B�\��@{����4@���!?QA;�,�@RΓ�#�ٿ K�ha��@]�hs(4@ӳX���!?�W�"��@v%�]c�ٿ̒_ż	�@)���4@�D�U�!?�"V��@s�u�ٿZL^��X�@_t;�
4@�ш�Ӑ!?u(����@s�u�ٿZL^��X�@_t;�
4@�ш�Ӑ!?u(����@s�u�ٿZL^��X�@_t;�
4@�ш�Ӑ!?u(����@s�u�ٿZL^��X�@_t;�
4@�ш�Ӑ!?u(����@s�u�ٿZL^��X�@_t;�
4@�ш�Ӑ!?u(����@e�S��ٿ���`IV�@-���4@�����!?"�w+�<�@�b���ٿ�ki��:�@M����4@g�Ұ��!?��}���@�b���ٿ�ki��:�@M����4@g�Ұ��!?��}���@�b���ٿ�ki��:�@M����4@g�Ұ��!?��}���@<<%���ٿ����V�@H!���4@C˿iՐ!?K��+��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@�8H��ٿW� ���@S?n�4@�yd��!?9{��@V��x�ٿ��`�9��@51r��3@(,�k��!?���B��@�[d�ЅٿY�U��@Uλ��4@���!�!?lµX��@�����{ٿ�)�9���@`��`G�3@c�q��!?�`��C��@�����{ٿ�)�9���@`��`G�3@c�q��!?�`��C��@�����{ٿ�)�9���@`��`G�3@c�q��!?�`��C��@�����{ٿ�)�9���@`��`G�3@c�q��!?�`��C��@�����{ٿ�)�9���@`��`G�3@c�q��!?�`��C��@��r;~ٿ��D�@�ű�g�3@@�`��!?_�z���@��r;~ٿ��D�@�ű�g�3@@�`��!?_�z���@�¨�|ٿ��PQ���@
�� _�3@64%�֐!?��H|�@�¨�|ٿ��PQ���@
�� _�3@64%�֐!?��H|�@r.��ׄٿ�G��O�@:�����3@�t��!?L��R�@SқI\�ٿr��<a��@gmY� 4@s�
�!?���'�\�@SқI\�ٿr��<a��@gmY� 4@s�
�!?���'�\�@SқI\�ٿr��<a��@gmY� 4@s�
�!?���'�\�@SқI\�ٿr��<a��@gmY� 4@s�
�!?���'�\�@�$wV}ٿ<W%�l��@�$��4@@�b���!?
(���@`3��ٿ��<]T/�@����	4@�H ސ!?�*�S���@`3��ٿ��<]T/�@����	4@�H ސ!?�*�S���@��l�ٿ���v)�@�"H�	4@�G���!?c��i$��@��l�ٿ���v)�@�"H�	4@�G���!?c��i$��@e1I!h�ٿ=�-�j�@%���	4@���4Ӑ!?v��P��@��J�ٿr�*V�@�N�34@���!?��t�KX�@��J�ٿr�*V�@�N�34@���!?��t�KX�@��J�ٿr�*V�@�N�34@���!?��t�KX�@��J�ٿr�*V�@�N�34@���!?��t�KX�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@����ٿ�Q�*i��@#�lb4@���	��!?�괨*�@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@7=׎��ٿ*��X���@6o�}=4@
��ː!?�y<I��@�Sex�ٿ�:�D>��@�5��4@ �+���!?Z�J��@�Sex�ٿ�:�D>��@�5��4@ �+���!?Z�J��@��]i݂ٿ�>֝� �@2�l]l4@<���!?0cm���@��]i݂ٿ�>֝� �@2�l]l4@<���!?0cm���@��]i݂ٿ�>֝� �@2�l]l4@<���!?0cm���@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@2Z%F��ٿs��� �@�η�k4@��=A��!?���@!�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@����J�ٿ&\��G��@��F�Q4@�S	��!??*�oci�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@Ĝ��ٿǅm[���@��֣4@zq܈��!?��s�T�@��Q��ٿ|�:[m��@\!��4@n����!?g��k���@��Q��ٿ|�:[m��@\!��4@n����!?g��k���@��Q��ٿ|�:[m��@\!��4@n����!?g��k���@Z	��ٿSW���@Bugx4@��x�i�!?�V��M��@Z	��ٿSW���@Bugx4@��x�i�!?�V��M��@Z	��ٿSW���@Bugx4@��x�i�!?�V��M��@�:�^{�ٿL�
����@����4@ѻ*;��!?�in<�@�:�^{�ٿL�
����@����4@ѻ*;��!?�in<�@�,��	�ٿŎ���@6�[j�4@#��v2�!?�K�-pC�@���ԋٿ��bgV{�@��:� 4@��ń�!?�_p�>�@���ԋٿ��bgV{�@��:� 4@��ń�!?�_p�>�@R��{f�ٿe��u�=�@���4@^�.b�!?�<T3�u�@R��{f�ٿe��u�=�@���4@^�.b�!?�<T3�u�@R��{f�ٿe��u�=�@���4@^�.b�!?�<T3�u�@R��{f�ٿe��u�=�@���4@^�.b�!?�<T3�u�@'����{ٿ��mf3p�@z(�N�4@��펕�!?���l�@'����{ٿ��mf3p�@z(�N�4@��펕�!?���l�@'����{ٿ��mf3p�@z(�N�4@��펕�!?���l�@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@��G�}ٿ������@Z�b4@�����!?�ڛuv��@j'^�ٿ�a�$m�@yjkB�4@������!?2����o�@j'^�ٿ�a�$m�@yjkB�4@������!?2����o�@j'^�ٿ�a�$m�@yjkB�4@������!?2����o�@j'^�ٿ�a�$m�@yjkB�4@������!?2����o�@�U7v	�ٿO��d�@1�m�4@��.鑐!?���Y��@�U7v	�ٿO��d�@1�m�4@��.鑐!?���Y��@�U7v	�ٿO��d�@1�m�4@��.鑐!?���Y��@In��P�ٿ.~����@�@Am4@��׿��!?�4�U��@In��P�ٿ.~����@�@Am4@��׿��!?�4�U��@In��P�ٿ.~����@�@Am4@��׿��!?�4�U��@In��P�ٿ.~����@�@Am4@��׿��!?�4�U��@In��P�ٿ.~����@�@Am4@��׿��!?�4�U��@�"0�{~ٿdن�.��@uq�4@�w�j�!?��A�@�"0�{~ٿdن�.��@uq�4@�w�j�!?��A�@�m���ٿ7��$�@N���4@F󰘐�!?){��j�@�m���ٿ7��$�@N���4@F󰘐�!?){��j�@�m���ٿ7��$�@N���4@F󰘐�!?){��j�@�m���ٿ7��$�@N���4@F󰘐�!?){��j�@�m���ٿ7��$�@N���4@F󰘐�!?){��j�@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�l���ٿ$K/���@�y�}I4@ �8!?[�v�L��@�(I�5�ٿ�a�S���@�jQ��4@vh��!?��o��Y�@�(I�5�ٿ�a�S���@�jQ��4@vh��!?��o��Y�@�(I�5�ٿ�a�S���@�jQ��4@vh��!?��o��Y�@�(I�5�ٿ�a�S���@�jQ��4@vh��!?��o��Y�@�(I�5�ٿ�a�S���@�jQ��4@vh��!?��o��Y�@�Iÿ�ٿ�n�J3��@��Rrd4@���.D�!?��Ql���@�Iÿ�ٿ�n�J3��@��Rrd4@���.D�!?��Ql���@�Iÿ�ٿ�n�J3��@��Rrd4@���.D�!?��Ql���@=����ٿD�'�n�@�w�4@ڧn�ϐ!?jU n
�@����ٿ@%���3�@61|*4@����!?W�+� ��@�<e9��ٿۯ�M�@���z�4@g$��!?�����7�@k�&���ٿ�j�z��@��94@��|���!?X��t�@щ���ٿE�kE�@,4@>'���!?/��{�@щ���ٿE�kE�@,4@>'���!?/��{�@щ���ٿE�kE�@,4@>'���!?/��{�@&g���ٿ��s�7��@���4@A��T��!?���C"X�@&g���ٿ��s�7��@���4@A��T��!?���C"X�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@A_Bm�ٿ*�7tP�@5��"4@�����!?!I�q[�@�kP�]�ٿ00���@��b)4@�x��!?��b���@�kP�]�ٿ00���@��b)4@�x��!?��b���@�kP�]�ٿ00���@��b)4@�x��!?��b���@�kP�]�ٿ00���@��b)4@�x��!?��b���@�kP�]�ٿ00���@��b)4@�x��!?��b���@�kP�]�ٿ00���@��b)4@�x��!?��b���@���=��ٿOa[2��@��X
4@՞D��!?��C 4�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@���š�ٿ��d�I�@��h�W4@�;)ؐ!?yYT�Y�@:ݠኊٿ�%���@�8�#4@�DD��!?��#f{�@:ݠኊٿ�%���@�8�#4@�DD��!?��#f{�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@(8��ٿC-Z�a��@�)�4@�?�!?J7fɰ�@��X�ٿ�d!>�@�$�9�4@����!?$<����@��X�ٿ�d!>�@�$�9�4@����!?$<����@��X�ٿ�d!>�@�$�9�4@����!?$<����@��X�ٿ�d!>�@�$�9�4@����!?$<����@��ve�ٿQ2��8�@؁l4@t��!?��z��@��ve�ٿQ2��8�@؁l4@t��!?��z��@��ve�ٿQ2��8�@؁l4@t��!?��z��@��ve�ٿQ2��8�@؁l4@t��!?��z��@hЀE�ٿ0�%���@WMQ�	4@�f֪�!?<#d�y��@�G�z΂ٿ�oR���@�Xn4@C����!?��y]3�@�G�z΂ٿ�oR���@�Xn4@C����!?��y]3�@�G�z΂ٿ�oR���@�Xn4@C����!?��y]3�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@{EͿ�ٿt'ZW���@�ݾ�K4@*$��!?��	&�@\�IHC�ٿΏD����@�q���4@3��A��!?��Q��@��j�U�ٿE��	���@A��f^4@W7w:��!?��3_7�@��j�U�ٿE��	���@A��f^4@W7w:��!?��3_7�@��j�U�ٿE��	���@A��f^4@W7w:��!?��3_7�@��j�U�ٿE��	���@A��f^4@W7w:��!?��3_7�@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@�;�G�ٿ
�A��@]�~��4@��.�Đ!?�h�����@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��>V�ٿ�z#v9x�@0m��4@�7�2z�!?c�W�q��@��^�ٿ�`Դ��@d�z�4@�)���!?��(!���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@��@�ٿ�2�����@�3�E��3@�Y��ʐ!?��� ���@�e�2�ٿ�#~`�@�|vN�4@'�d���!?��[��@�e�2�ٿ�#~`�@�|vN�4@'�d���!?��[��@�e�2�ٿ�#~`�@�|vN�4@'�d���!?��[��@��PP�ٿ�'t�a�@)��^�4@ ��ݐ!?dM}�R�@��PP�ٿ�'t�a�@)��^�4@ ��ݐ!?dM}�R�@��PP�ٿ�'t�a�@)��^�4@ ��ݐ!?dM}�R�@��PP�ٿ�'t�a�@)��^�4@ ��ݐ!?dM}�R�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��!Cp�ٿL<����@�R��4@x����!?����EG�@��\�P�ٿ:/)��@�b�4@��N���!?�s]_��@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@l�8R��ٿE�|�Br�@�Iߣ�4@��O�ѐ!?�9d|���@A8�ٿ�\�(��@�䴿�4@~�6�Ð!?�#�O���@A8�ٿ�\�(��@�䴿�4@~�6�Ð!?�#�O���@A8�ٿ�\�(��@�䴿�4@~�6�Ð!?�#�O���@��<���ٿ�S*��@�*�0�4@Ĵ�&�!?͹r����@��<���ٿ�S*��@�*�0�4@Ĵ�&�!?͹r����@��<���ٿ�S*��@�*�0�4@Ĵ�&�!?͹r����@��<���ٿ�S*��@�*�0�4@Ĵ�&�!?͹r����@��<���ٿ�S*��@�*�0�4@Ĵ�&�!?͹r����@����zٿ���]��@Z��.�4@{��6��!?��>oe!�@����zٿ���]��@Z��.�4@{��6��!?��>oe!�@*�rwٿ���&��@�\���4@�M%��!?M[����@*�rwٿ���&��@�\���4@�M%��!?M[����@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�!�ٿw6��F��@�s��4@�2��7�!?��-~��@�o#�ٿ2�d�{�@����4@a��FH�!?8�|�}�@�����ٿY�P���@�2�S~4@���l�!?6��+ź�@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@< w�l�ٿ�����@��Vw&4@��;��!?<�>e��@��cD��ٿ]����@�G0�b4@s�0v�!?ߝ&���@��cD��ٿ]����@�G0�b4@s�0v�!?ߝ&���@��cD��ٿ]����@�G0�b4@s�0v�!?ߝ&���@��cD��ٿ]����@�G0�b4@s�0v�!?ߝ&���@��cD��ٿ]����@�G0�b4@s�0v�!?ߝ&���@>x拗�ٿ��'q)(�@d�u4@!�O��!?p���S�@>x拗�ٿ��'q)(�@d�u4@!�O��!?p���S�@ww�ٿz�G0���@�N&J4@)0����!?9�T���@ �/�ٿ	Fw� �@�Q�&4@F=e�!?��K{��@ �/�ٿ	Fw� �@�Q�&4@F=e�!?��K{��@ �/�ٿ	Fw� �@�Q�&4@F=e�!?��K{��@ �/�ٿ	Fw� �@�Q�&4@F=e�!?��K{��@pz���ٿSϒϐ�@�)D4@�М�!?8v�0&�@pz���ٿSϒϐ�@�)D4@�М�!?8v�0&�@�p��ٿ�75����@��e�4@��\�Ɛ!?�Lc����@m'����ٿ�b�v���@��K@4@��7Đ!?[u͉�E�@m'����ٿ�b�v���@��K@4@��7Đ!?[u͉�E�@�j[���ٿ�y��<i�@�2O+4@�G�(�!?AB���\�@3w�PW�ٿ2r�[�(�@	��� 4@���!?b*T|��@3w�PW�ٿ2r�[�(�@	��� 4@���!?b*T|��@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@%��8�ٿ��λЂ�@�����4@ĝr=ߐ!?� �tDn�@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@�Tj<��ٿA�&�u�@ZE$�4@��X9��!?��J�9 �@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@en�]�ٿ��.���@��>�4@�AGН�!?b ֊��@�:ʃٿ�ȶ�?��@��E��4@푍���!?>1��W��@�:ʃٿ�ȶ�?��@��E��4@푍���!?>1��W��@�:ʃٿ�ȶ�?��@��E��4@푍���!?>1��W��@�:ʃٿ�ȶ�?��@��E��4@푍���!?>1��W��@q-��ٿ$��'V��@����Q 4@�Q���!?L?��M.�@q-��ٿ$��'V��@����Q 4@�Q���!?L?��M.�@q-��ٿ$��'V��@����Q 4@�Q���!?L?��M.�@���W{�ٿUrǔ��@;�s%4@�n�Ȑ!?&}�����@���W{�ٿUrǔ��@;�s%4@�n�Ȑ!?&}�����@�G�<�ٿ (����@�C⽄4@_?U	�!?ԍ�}�u�@�G�<�ٿ (����@�C⽄4@_?U	�!?ԍ�}�u�@�G�<�ٿ (����@�C⽄4@_?U	�!?ԍ�}�u�@�G�<�ٿ (����@�C⽄4@_?U	�!?ԍ�}�u�@�G�<�ٿ (����@�C⽄4@_?U	�!?ԍ�}�u�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@eq��k�ٿgG�i�o�@=�O��4@6j�ڐ!?��M�@R�?v�ٿ�
jL�T�@��#4@��j�!?��+�G�@R�?v�ٿ�
jL�T�@��#4@��j�!?��+�G�@R�?v�ٿ�
jL�T�@��#4@��j�!?��+�G�@R�?v�ٿ�
jL�T�@��#4@��j�!?��+�G�@�A�O�ٿ��Q0���@�^Ȱn4@�����!?�'�&P�@^�����ٿw�1��k�@��3�4@$��Ӑ!?M%�p
>�@^�����ٿw�1��k�@��3�4@$��Ӑ!?M%�p
>�@��kJ��ٿ�ɮ�F�@�����4@} �gӐ!?��^��M�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@ŝG
�ٿ빟aI�@B]��
4@��ܐ!?��@�@��J�ٿ�=E���@��a��4@d�w��!?W����@��J�ٿ�=E���@��a��4@d�w��!?W����@��J�ٿ�=E���@��a��4@d�w��!?W����@(=ӛ��ٿǮ��E�@�n��s4@�9���!?Ԇ����@(=ӛ��ٿǮ��E�@�n��s4@�9���!?Ԇ����@(=ӛ��ٿǮ��E�@�n��s4@�9���!?Ԇ����@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@�u3'%�ٿ�`2����@����c4@ �Ӑ!?g�c+��@f�Ib�ٿ�Sh%?�@h]QWP4@�Aϩ�!?��R���@f�Ib�ٿ�Sh%?�@h]QWP4@�Aϩ�!?��R���@5'���ٿ��.��@l{D��4@��v�!?#-��T��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@ۼ�E]�ٿ#<�k��@.�%��4@�V䯐!?���Y-��@�4���ٿɽ�c��@N]�^�4@#v���!?��
$@�@�4���ٿɽ�c��@N]�^�4@#v���!?��
$@�@�}��g�ٿv���l�@-�p�4@�n��!?Ĉ�y� �@���dL�ٿ�ScJ���@כ�p 4@�>hŐ!?���X�@���dL�ٿ�ScJ���@כ�p 4@�>hŐ!?���X�@���dL�ٿ�ScJ���@כ�p 4@�>hŐ!?���X�@���dL�ٿ�ScJ���@כ�p 4@�>hŐ!?���X�@���Td�ٿdND��@�\��4@�ܔ
�!?��H�C��@���Td�ٿdND��@�\��4@�ܔ
�!?��H�C��@���Td�ٿdND��@�\��4@�ܔ
�!?��H�C��@��ȉ/�ٿ��6Ro�@gzF�4@����!?� !A�@��ȉ/�ٿ��6Ro�@gzF�4@����!?� !A�@ '�d}ٿ���0��@��uv4@my���!?~}���@ '�d}ٿ���0��@��uv4@my���!?~}���@�~�аyٿ�l��J�@��i4@:��Ŷ�!?K�����@�~�аyٿ�l��J�@��i4@:��Ŷ�!?K�����@�ul!	�ٿ�ҙ㳔�@9M��{4@}����!?F]��� �@�ul!	�ٿ�ҙ㳔�@9M��{4@}����!?F]��� �@�ul!	�ٿ�ҙ㳔�@9M��{4@}����!?F]��� �@�ul!	�ٿ�ҙ㳔�@9M��{4@}����!?F]��� �@�RAyb�ٿK�9�j�@"��	4@�VDʹ�!?�v����@�IP�H�ٿ�m�/IQ�@��J��4@�'�k̐!?���Ʈ:�@�IP�H�ٿ�m�/IQ�@��J��4@�'�k̐!?���Ʈ:�@�IP�H�ٿ�m�/IQ�@��J��4@�'�k̐!?���Ʈ:�@�IP�H�ٿ�m�/IQ�@��J��4@�'�k̐!?���Ʈ:�@�IP�H�ٿ�m�/IQ�@��J��4@�'�k̐!?���Ʈ:�@���Fr�ٿ+Q��W�@B���4@���Q��!?7��i���@���Fr�ٿ+Q��W�@B���4@���Q��!?7��i���@���Fr�ٿ+Q��W�@B���4@���Q��!?7��i���@���Fr�ٿ+Q��W�@B���4@���Q��!?7��i���@ހ�9S�ٿ�;�L>�@ 9�*"4@��^֐!?J�����@�.1%7�ٿĖ;����@r:F0.4@Å �֐!?D�M`�@�.1%7�ٿĖ;����@r:F0.4@Å �֐!?D�M`�@�rf��ٿ�����@���hJ4@:����!?8V�Q�	�@�rf��ٿ�����@���hJ4@:����!?8V�Q�	�@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@�����ٿCgđ�[�@Ƽt�4@�J�ݐ!?K�Q����@��Y�ٿ�Ƙ�W\�@�V���4@z�)Ր!?�X��O�@��Y�ٿ�Ƙ�W\�@�V���4@z�)Ր!?�X��O�@�@򌃁ٿ�%O�@*b���4@	��F �!?N<�k)*�@�@򌃁ٿ�%O�@*b���4@	��F �!?N<�k)*�@�@򌃁ٿ�%O�@*b���4@	��F �!?N<�k)*�@�@򌃁ٿ�%O�@*b���4@	��F �!?N<�k)*�@�@򌃁ٿ�%O�@*b���4@	��F �!?N<�k)*�@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@�[IjӈٿB�D�M�@�&̇�4@��6�Ɛ!?������@r�F�o�ٿ�S�q�@cԖ4"4@��R|��!?Mt���T�@r�F�o�ٿ�S�q�@cԖ4"4@��R|��!?Mt���T�@r�F�o�ٿ�S�q�@cԖ4"4@��R|��!?Mt���T�@r�F�o�ٿ�S�q�@cԖ4"4@��R|��!?Mt���T�@r�F�o�ٿ�S�q�@cԖ4"4@��R|��!?Mt���T�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@�@;�ʉٿ1e����@�)�P4@2b�Ґ!? �IWZ�@$����ٿ���pً�@�*���4@��@�!?�P2kh��@$����ٿ���pً�@�*���4@��@�!?�P2kh��@$����ٿ���pً�@�*���4@��@�!?�P2kh��@$����ٿ���pً�@�*���4@��@�!?�P2kh��@$����ٿ���pً�@�*���4@��@�!?�P2kh��@$����ٿ���pً�@�*���4@��@�!?�P2kh��@|���@�ٿ||�П�@Q*�N4@r*�Ȑ!?�Yp,J��@|���@�ٿ||�П�@Q*�N4@r*�Ȑ!?�Yp,J��@ڑL�ٿ�J/I��@�#��Q4@ �|Tڐ!?�o�&��@ڑL�ٿ�J/I��@�#��Q4@ �|Tڐ!?�o�&��@��wt��ٿ�3}����@� {�W4@rNh���!?쨒����@��wt��ٿ�3}����@� {�W4@rNh���!?쨒����@v�[���ٿ1P�Ȯ��@+�Ư�4@v��8��!?�'��{��@v�[���ٿ1P�Ȯ��@+�Ư�4@v��8��!?�'��{��@K[�-�ٿ���A���@d���4@¾7�Ð!?|鞅sE�@j�2�ςٿ˯ʫ�M�@�%*�s	4@�&Qߐ!?B��ߏ�@j�2�ςٿ˯ʫ�M�@�%*�s	4@�&Qߐ!?B��ߏ�@j�2�ςٿ˯ʫ�M�@�%*�s	4@�&Qߐ!?B��ߏ�@j�2�ςٿ˯ʫ�M�@�%*�s	4@�&Qߐ!?B��ߏ�@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@�'��Q�ٿP��ep*�@�֜3�4@d�����!?[>o ���@ V
͟�ٿ�߽�S��@�:|�n4@�-G� �!?W�&u�-�@����~ٿbd�� �@Ŵ�L�4@�;���!?�4�E+�@����~ٿbd�� �@Ŵ�L�4@�;���!?�4�E+�@����~ٿbd�� �@Ŵ�L�4@�;���!?�4�E+�@�눌��ٿ�����2�@�(�Z(4@�;C���!?CAh��@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@�;U��ٿ�Տ�C�@��^�4@A����!?P���]�@%��ٿ�"��@�{�� 4@� OtÐ!?:j��@��@%��ٿ�"��@�{�� 4@� OtÐ!?:j��@��@<u)�ٿ���E%w�@6�7Ύ4@�=yX��!?+x ֪�@Y7'R��ٿ�N*(�@W��� 4@��9��!?cC�r��@�$֔�ٿO��@;[]��4@��%��!?2��8��@�$֔�ٿO��@;[]��4@��%��!?2��8��@�$֔�ٿO��@;[]��4@��%��!?2��8��@�$֔�ٿO��@;[]��4@��%��!?2��8��@y�o{��ٿ>�����@K$Pι4@f��p��!?7U��-�@y�o{��ٿ>�����@K$Pι4@f��p��!?7U��-�@,�-��ٿy����@�93��4@�G�D�!?�įѩ��@,�-��ٿy����@�93��4@�G�D�!?�įѩ��@,�-��ٿy����@�93��4@�G�D�!?�įѩ��@,�-��ٿy����@�93��4@�G�D�!?�įѩ��@T$aH�}ٿ���!��@)@J�4@�ǯa|�!?�	�b��@T$aH�}ٿ���!��@)@J�4@�ǯa|�!?�	�b��@f#�5j�ٿ�BȨ�v�@#컖4@��g��!?�	�?`�@y��<��ٿ�$�:���@po��4@�HjȐ!?Bx��0�@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@�U���ٿ3���Z��@�#܊F�3@���oՐ!?a��G��@C�H��ٿ�Bf���@$b��3@���א!?	���@����ٿ�&���@a�[m 4@��?�!?��mt��@�F��O}ٿ�H�aq��@��I{4@Wlj���!?�h��j�@�F��O}ٿ�H�aq��@��I{4@Wlj���!?�h��j�@�F��O}ٿ�H�aq��@��I{4@Wlj���!?�h��j�@�F��O}ٿ�H�aq��@��I{4@Wlj���!?�h��j�@�F��O}ٿ�H�aq��@��I{4@Wlj���!?�h��j�@F/�n�ٿ�W`��@h~�@F4@^Ϝa�!?n���"��@C����ٿ�x!20��@BƂ��4@9�3O��!?����ۂ�@C����ٿ�x!20��@BƂ��4@9�3O��!?����ۂ�@���번ٿ)�X�f�@"��.4@��Tˇ�!?�ui�5/�@���번ٿ)�X�f�@"��.4@��Tˇ�!?�ui�5/�@���번ٿ)�X�f�@"��.4@��Tˇ�!?�ui�5/�@���번ٿ)�X�f�@"��.4@��Tˇ�!?�ui�5/�@���번ٿ)�X�f�@"��.4@��Tˇ�!?�ui�5/�@�Jc|�ٿ�ё����@&X?B4@V�x��!?>�En)�@�Jc|�ٿ�ё����@&X?B4@V�x��!?>�En)�@�Jc|�ٿ�ё����@&X?B4@V�x��!?>�En)�@;�SŏٿÒ.1�@����4@��>_�!?�b�N�@�����ٿ��?���@����4@����!?D��6���@�����ٿ��?���@����4@����!?D��6���@�����ٿ��?���@����4@����!?D��6���@�����ٿ��?���@����4@����!?D��6���@��暅ٿ��s�8�@C�ޛ�4@{��>@�!?9�w�]�@��暅ٿ��s�8�@C�ޛ�4@{��>@�!?9�w�]�@��暅ٿ��s�8�@C�ޛ�4@{��>@�!?9�w�]�@��暅ٿ��s�8�@C�ޛ�4@{��>@�!?9�w�]�@��暅ٿ��s�8�@C�ޛ�4@{��>@�!?9�w�]�@;ES��ٿ�P�5��@L-d�84@ZLK�c�!?]�8���@;ES��ٿ�P�5��@L-d�84@ZLK�c�!?]�8���@;ES��ٿ�P�5��@L-d�84@ZLK�c�!?]�8���@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�����ٿQi���S�@��G}�4@��8d�!?�������@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�D�-�ٿ��p =�@�ko�4@�g� �!?�}�w�@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�-{a?�ٿUdH�2U�@�9�+�4@��􂧐!?��$���@�[j��ٿ�a�\"�@a����4@�a���!?ӌ�����@�[j��ٿ�a�\"�@a����4@�a���!?ӌ�����@�[j��ٿ�a�\"�@a����4@�a���!?ӌ�����@�[j��ٿ�a�\"�@a����4@�a���!?ӌ�����@"]<ٿ��u7'�@\�ݳ�4@�T  �!?G����@"]<ٿ��u7'�@\�ݳ�4@�T  �!?G����@��63N�ٿ� � ��@_)j�4@�����!?����x
�@��63N�ٿ� � ��@_)j�4@�����!?����x
�@��S�ٿs�A�P�@����4@�`tD��!?��ž��@�ę���ٿCO��e��@��W�S4@���͐!?B�E=���@�ę���ٿCO��e��@��W�S4@���͐!?B�E=���@�ę���ٿCO��e��@��W�S4@���͐!?B�E=���@�ę���ٿCO��e��@��W�S4@���͐!?B�E=���@P��P�ٿ�Dٸk�@�z�O�4@Qx�ې!?@�1��"�@dWEDK�ٿ���%��@J�G�4@�����!?���#��@dWEDK�ٿ���%��@J�G�4@�����!?���#��@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@K�xF�ٿL��#��@�?]94@G���!?�r���4�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@�N��v�ٿJ�&�Y�@{��4@�1o��!?��r/k�@AC��8�ٿ�HȘQ��@��H=B4@+\s�k�!?�F�7a}�@AC��8�ٿ�HȘQ��@��H=B4@+\s�k�!?�F�7a}�@�N���ٿ�e�-3�@���jt4@t�=`�!?s�e�s��@�N���ٿ�e�-3�@���jt4@t�=`�!?s�e�s��@�Ay�d�ٿ}i��Z�@�Z�"� 4@�k(>��!?�m�uof�@���ŏٿ�04_d��@Q/�I@4@�j�ڹ�!?S��~��@����ٿ،P���@�L?�4@1�!?��j4�@�u�ٿ߀����@�wB��4@[��:�!?�vЖz�@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@���鏃ٿm�֓��@�RL1�4@�7��ߐ!?�!��@�ȁ�ٿ!#x���@�c�
4@���3Ґ!?���Ϊ�@�ȁ�ٿ!#x���@�c�
4@���3Ґ!?���Ϊ�@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@�̖C:{ٿQSF����@OӨ�4@{�E���!?�s#����@��&���ٿ� �MR&�@E9�e4@5@��ѐ!?�Q
F7`�@��&���ٿ� �MR&�@E9�e4@5@��ѐ!?�Q
F7`�@��&���ٿ� �MR&�@E9�e4@5@��ѐ!?�Q
F7`�@��&���ٿ� �MR&�@E9�e4@5@��ѐ!?�Q
F7`�@��&���ٿ� �MR&�@E9�e4@5@��ѐ!?�Q
F7`�@�
�TU�ٿ��}��C�@g�?4@���~ڐ!?��g�U�@�
�TU�ٿ��}��C�@g�?4@���~ڐ!?��g�U�@^#�Cv�ٿ
�A�)��@���R"4@d�V��!?��
,��@^#�Cv�ٿ
�A�)��@���R"4@d�V��!?��
,��@^#�Cv�ٿ
�A�)��@���R"4@d�V��!?��
,��@^#�Cv�ٿ
�A�)��@���R"4@d�V��!?��
,��@^#�Cv�ٿ
�A�)��@���R"4@d�V��!?��
,��@�N\�ٿ��!S�@�?0~4@������!?����@�@�N\�ٿ��!S�@�?0~4@������!?����@�@�N\�ٿ��!S�@�?0~4@������!?����@�@�N\�ٿ��!S�@�?0~4@������!?����@�@}�A��ٿ�/D�F��@�ڀ&�4@�,p���!?�zK����@}�A��ٿ�/D�F��@�ڀ&�4@�,p���!?�zK����@}�A��ٿ�/D�F��@�ڀ&�4@�,p���!?�zK����@R�J��ٿYX����@�*�4@�����!?&�u���@R�J��ٿYX����@�*�4@�����!?&�u���@R�J��ٿYX����@�*�4@�����!?&�u���@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@��f�@�ٿq���5��@m4�K}4@h{9t�!?��	k��@�ޕ���ٿX�#
��@�q]Aa4@��J��!?�}��7�@�ޕ���ٿX�#
��@�q]Aa4@��J��!?�}��7�@�ޕ���ٿX�#
��@�q]Aa4@��J��!?�}��7�@�ޕ���ٿX�#
��@�q]Aa4@��J��!?�}��7�@`J!���ٿ�_�cζ�@�{E=;4@D���!?�Xn���@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@Kag��ٿ_�P��@���w4@�w!ː!?�M,Y-�@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@������ٿ#���Ӟ�@�>!�4@��۷Ґ!?���P���@.����ٿ;J�=��@W.��?4@��o��!?���S���@.����ٿ;J�=��@W.��?4@��o��!?���S���@d0q��ٿTH�:W�@JS��]	4@�_�mϐ!?^w#�|��@d0q��ٿTH�:W�@JS��]	4@�_�mϐ!?^w#�|��@�Lc�/�ٿ �����@����4@?�P˿�!?������@�Lc�/�ٿ �����@����4@?�P˿�!?������@�Lc�/�ٿ �����@����4@?�P˿�!?������@�Lc�/�ٿ �����@����4@?�P˿�!?������@�Lc�/�ٿ �����@����4@?�P˿�!?������@���=�ٿ�5�f�@�r�!4@s�
�ߐ!?���nO��@���=�ٿ�5�f�@�r�!4@s�
�ߐ!?���nO��@#"�̶�ٿ��'��@�y��(4@�
���!? 0M�7_�@#"�̶�ٿ��'��@�y��(4@�
���!? 0M�7_�@#"�̶�ٿ��'��@�y��(4@�
���!? 0M�7_�@#"�̶�ٿ��'��@�y��(4@�
���!? 0M�7_�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@��.|�ٿ�q�J�@�#�!�4@�V}>��!?�F�!�@ ~1N׏ٿ������@݀��4@Ey�ᢐ!?n�n*P��@ ~1N׏ٿ������@݀��4@Ey�ᢐ!?n�n*P��@ ~1N׏ٿ������@݀��4@Ey�ᢐ!?n�n*P��@ ~1N׏ٿ������@݀��4@Ey�ᢐ!?n�n*P��@w��Տٿ+a��,��@�<�k4@����!?��J��-�@w��Տٿ+a��,��@�<�k4@����!?��J��-�@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@WQ��ȁٿ����fB�@)T1l4@��Ѕ��!?����v��@6]�6Ѕٿ�\�q���@� �ٕ4@���b�!?أ$��@�6�.1�ٿ��B���@��{G�4@h�!<v�!?�Pr�@�6�.1�ٿ��B���@��{G�4@h�!<v�!?�Pr�@�|���ٿ���~��@o��n4@م	a��!? P�q�@�|���ٿ���~��@o��n4@م	a��!? P�q�@�|���ٿ���~��@o��n4@م	a��!? P�q�@T}n��ٿl��2uP�@ЂM@4@i����!?g"�1y�@T}n��ٿl��2uP�@ЂM@4@i����!?g"�1y�@T}n��ٿl��2uP�@ЂM@4@i����!?g"�1y�@T5̏ٿ[j^6��@
�Cj?4@k��Ԯ�!?!�����@T5̏ٿ[j^6��@
�Cj?4@k��Ԯ�!?!�����@T5̏ٿ[j^6��@
�Cj?4@k��Ԯ�!?!�����@T5̏ٿ[j^6��@
�Cj?4@k��Ԯ�!?!�����@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@P̱�+�ٿ�}s���@qYx�4@٫�	��!?��!Z�'�@Y6�o�ٿ@/v �Y�@Jh���4@o#��!?~���b��@Y6�o�ٿ@/v �Y�@Jh���4@o#��!?~���b��@Y6�o�ٿ@/v �Y�@Jh���4@o#��!?~���b��@Y6�o�ٿ@/v �Y�@Jh���4@o#��!?~���b��@�Y�ٿ�Փ1��@�pP{:4@�~2�!?_��<�6�@�Y�ٿ�Փ1��@�pP{:4@�~2�!?_��<�6�@�Y�ٿ�Փ1��@�pP{:4@�~2�!?_��<�6�@�Y�ٿ�Փ1��@�pP{:4@�~2�!?_��<�6�@�tх��ٿ�����@�ΠN44@ q���!?��A�&�@t�Sָ�ٿ0�2��@iO�
W4@���Ȑ!?1�D׻��@��+6�ٿ�ᩴ���@z��"�4@_P)�w�!?i�2+��@��+6�ٿ�ᩴ���@z��"�4@_P)�w�!?i�2+��@��+6�ٿ�ᩴ���@z��"�4@_P)�w�!?i�2+��@��+6�ٿ�ᩴ���@z��"�4@_P)�w�!?i�2+��@��+6�ٿ�ᩴ���@z��"�4@_P)�w�!?i�2+��@S8Î]�ٿ��a���@*#<)�4@�9e��!?������@��ˌ͊ٿA�XX!��@�$��'4@՘#�!?�8�P�@>���ٿ��+W9�@@*7��4@v���<�!?O&�h��@�;�⮇ٿA�.���@9�Y�4@�+��6�!?@S]���@�;�⮇ٿA�.���@9�Y�4@�+��6�!?@S]���@w2�tU�ٿe��_?�@z�5�4@iLz��!?�d��b�@w2�tU�ٿe��_?�@z�5�4@iLz��!?�d��b�@w2�tU�ٿe��_?�@z�5�4@iLz��!?�d��b�@w2�tU�ٿe��_?�@z�5�4@iLz��!?�d��b�@w2�tU�ٿe��_?�@z�5�4@iLz��!?�d��b�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�̮ٜ�ٿ������@��"44@�n(��!?�G��0�@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�fO�ٿ���_�@���ַ4@!f*ڐ!?��AU��@�I��L�ٿc�!���@I�}2�
4@��5�l�!?�x:[=��@�I��L�ٿc�!���@I�}2�
4@��5�l�!?�x:[=��@�I��L�ٿc�!���@I�}2�
4@��5�l�!?�x:[=��@X���g�ٿ�p�Ku��@D���z
4@�汐!?C�;���@X���g�ٿ�p�Ku��@D���z
4@�汐!?C�;���@X���g�ٿ�p�Ku��@D���z
4@�汐!?C�;���@X���g�ٿ�p�Ku��@D���z
4@�汐!?C�;���@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@������ٿ     ��@      4@�t><K�!?S����+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�v�+�ٿĺ�����@ݸ�� 4@����9�!?8S�u�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@�U��ٿ�e}~���@+(����3@��sUs�!?��XY�+�@���o��ٿ1�ry���@&> 4@�1���!?;X5�+�@���o��ٿ1�ry���@&> 4@�1���!?;X5�+�@���o��ٿ1�ry���@&> 4@�1���!?;X5�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@������ٿs�\���@��U 4@��~���!?�Vo<�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@9�q?��ٿ_�KM���@�V�� 4@!e�ק�!?^]B�+�@Ǭ�6˙ٿ�K�8���@��B 4@8s�x\�!? 9�C�+�@Ǭ�6˙ٿ�K�8���@��B 4@8s�x\�!? 9�C�+�@��șٿ���@���@c�U 4@y⿛&�!?��E�+�@�=�Ιٿ�4�:���@�<� 4@ؠ�R��!?Ĳ�R�+�@�=�Ιٿ�4�:���@�<� 4@ؠ�R��!?Ĳ�R�+�@>]̙ٿ��D���@�� 4@__I���!?��K�+�@>]̙ٿ��D���@�� 4@__I���!?��K�+�@�$Ιٿ�4j#���@���� 4@��?h�!?�%B�+�@Q��˙ٿV�&���@�y� 4@��W�!?�m�;�+�@Q��˙ٿV�&���@�y� 4@��W�!?�m�;�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@�Epbԙٿ�M�,���@;[oh 4@�F8�א!?��3�+�@���֙ٿ��9���@�(�� 4@L#~j!?�&?�+�@���֙ٿ��9���@�(�� 4@L#~j!?�&?�+�@Lx��ՙٿ��n2���@�ۛ9 4@`�U"m�!?)�@�+�@|V��ՙٿA��3���@} �� 4@j]x��!?H|>@�+�@|V��ՙٿA��3���@} �� 4@j]x��!?H|>@�+�@|V��ՙٿA��3���@} �� 4@j]x��!?H|>@�+�@��@̙ٿ}6�7���@��y� 4@��!?,�@�+�@��@̙ٿ}6�7���@��y� 4@��!?,�@�+�@w����ٿU�<���@�<� 4@�;�V��!?���A�+�@w����ٿU�<���@�<� 4@�;�V��!?���A�+�@Ů1@��ٿ9ː>���@�\ 4@�:p�!?V��M�+�@Ů1@��ٿ9ː>���@�\ 4@�:p�!?V��M�+�@Ů1@��ٿ9ː>���@�\ 4@�:p�!?V��M�+�@�-6���ٿ�˾L���@ޏ�� 4@����~�!?��M�+�@첬2��ٿ-��Q���@R��� 4@�Z��!?�^YO�+�@o^s��ٿ�
�L���@
s�} 4@ph�֐!?k^N�+�@o^s��ٿ�
�L���@
s�} 4@ph�֐!?k^N�+�@o^s��ٿ�
�L���@
s�} 4@ph�֐!?k^N�+�@o^s��ٿ�
�L���@
s�} 4@ph�֐!?k^N�+�@��K鯙ٿ��iS���@G�� 4@X����!?���O�+�@��K鯙ٿ��iS���@G�� 4@X����!?���O�+�@l��f��ٿB��]���@��Q� 4@��Reؐ!?�|�U�+�@��A��ٿ��[���@���� 4@����̐!?�n]T�+�@��A��ٿ��[���@���� 4@����̐!?�n]T�+�@��A��ٿ��[���@���� 4@����̐!?�n]T�+�@��A��ٿ��[���@���� 4@����̐!?�n]T�+�@�O����ٿ�ܳ^���@��X
 4@��İې!?���R�+�@�O����ٿ�ܳ^���@��X
 4@��İې!?���R�+�@HBZ��ٿO�,T���@uT� 4@i�XPt�!?���Q�+�@�3?��ٿn��T���@�X�o 4@ϟ��~�!?yM�T�+�@��~��ٿ��ON���@�պ 4@�Z���!?�C�T�+�@9����ٿ�F���@�p�R 4@�Q5f��!?L�R�+�@��힑�ٿ��.Q���@t��� 4@�[���!?���Q�+�@��힑�ٿ��.Q���@t��� 4@�[���!?���Q�+�@��힑�ٿ��.Q���@t��� 4@�[���!?���Q�+�@R��䑙ٿ��[���@!�� 4@f�ԅ�!?!ƀT�+�@��;h��ٿ���Y���@綧 4@D��~�!?��S�+�@��;h��ٿ���Y���@綧 4@D��~�!?��S�+�@��;h��ٿ���Y���@綧 4@D��~�!?��S�+�@]A~��ٿ���V���@!y�� 4@� ��֐!?�]N�+�@���ٿ*v�V���@r��' 4@L�%_]�!?��4M�+�@j2`h��ٿgV���@$� 4@�#l�G�!?@�MK�+�@a\���ٿ�~HQ���@�Y� 4@t��
�!?.b I�+�@gl�ٿXҦL���@�d� 4@��<u��!?��G�+�@��΀�ٿ���P���@ɏ 4@��UՐ!?=v J�+�@�c!��ٿ���N���@$Ⴏ 4@yc�Đ!?�/xL�+�@�c!��ٿ���N���@$Ⴏ 4@yc�Đ!?�/xL�+�@�c!��ٿ���N���@$Ⴏ 4@yc�Đ!?�/xL�+�@�c!��ٿ���N���@$Ⴏ 4@yc�Đ!?�/xL�+�@n��-|�ٿ$|FO���@F`�L 4@/W���!?�M�+�@�M�u�ٿ�HZS���@��yK	 4@|���Ő!?�O�+�@���$n�ٿHX���@����	 4@�l~&�!?U�V�+�@���$n�ٿHX���@����	 4@�l~&�!?U�V�+�@���$n�ٿHX���@����	 4@�l~&�!?U�V�+�@e��t�ٿ�|W���@��*�	 4@�����!?�єT�+�@e��t�ٿ�|W���@��*�	 4@�����!?�єT�+�@bF7�x�ٿ�+j[���@n�:� 4@�+M/��!?o�uU�+�@�_ Ji�ٿ���X���@Q�	 4@W
Qy�!?��[X�+�@-�WAk�ٿ��P���@Ũ��	 4@��qː!?��kZ�+�@�[�m�ٿ؍5P���@�z��	 4@(DD�ݐ!?�%�W�+�@����i�ٿ��8R���@��M	 4@-1
�!?¦�W�+�@����i�ٿ��8R���@��M	 4@-1
�!?¦�W�+�@����i�ٿ��8R���@��M	 4@-1
�!?¦�W�+�@����i�ٿ��8R���@��M	 4@-1
�!?¦�W�+�@����i�ٿ��8R���@��M	 4@-1
�!?¦�W�+�@c^��v�ٿ�^�S���@��۞ 4@u26\�!?��jO�+�@"/�i�ٿgY�S���@<�s� 4@mE���!?�6�N�+�@ ��^�ٿ�3+O���@{��	 4@��;Ր!?;��R�+�@ ��^�ٿ�3+O���@{��	 4@��;Ր!?;��R�+�@��E�a�ٿB
R���@�T�u	 4@/����!?�sR�+�@��E�a�ٿB
R���@�T�u	 4@/����!?�sR�+�@\�_�ٿ�L���@�x"d	 4@��H���!?mR�+�@���W_�ٿF8P���@J���	 4@��"�
�!?�#JT�+�@C�+'[�ٿ\\�I���@_��	 4@�O)�!?�OP�+�@C�+'[�ٿ\\�I���@_��	 4@�O)�!?�OP�+�@��W�ٿ��RK���@<��	 4@9A�!?�^�T�+�@����c�ٿ�oH���@���C	 4@qY1�"�!?:��V�+�@����c�ٿ�oH���@���C	 4@qY1�"�!?:��V�+�@Fz9 j�ٿ'k�L���@�~�T	 4@����!?v/FU�+�@����j�ٿ?��S���@.��� 4@s)�|L�!?�T�+�@V�h�j�ٿ�3K���@@z�� 4@�m�1q�!?㚻T�+�@�~Y�x�ٿ��&S���@�t�n 4@ĸ܁T�!?���Q�+�@�~Y�x�ٿ��&S���@�t�n 4@ĸ܁T�!?���Q�+�@%I�n�ٿ���S���@FE�� 4@��&C�!?�GqW�+�@%I�n�ٿ���S���@FE�� 4@��&C�!?�GqW�+�@���m�ٿ]�:V���@�K9� 4@���|}�!?ds�Y�+�@�$q�ٿT|U���@9%C� 4@0j�ޘ�!?�Z*W�+�@�$q�ٿT|U���@9%C� 4@0j�ޘ�!?�Z*W�+�@{1�2h�ٿ�2�H���@��� 4@�͌�!?��V�+�@Dəg�ٿ鋶F���@w�� 4@���g�!?؀ Y�+�@Dəg�ٿ鋶F���@w�� 4@���g�!?؀ Y�+�@��h�ٿ%�A���@���� 4@�9S���!?��bS�+�@�V��b�ٿ`��9���@͞�	 4@Su��Ő!?)_nT�+�@\��e�ٿ���7���@%F� 4@�"�̐!?#��T�+�@���hW�ٿox�;���@����	 4@�V�Q�!?%��W�+�@1�TL�ٿZYF5���@�ymc
 4@`7��!?N��[�+�@����@�ٿ�"�,���@��� 4@x]���!?�U�]�+�@����@�ٿ�"�,���@��� 4@x]���!?�U�]�+�@�ACdG�ٿA2�1���@��
 4@$_�\ݐ!?H,�Z�+�@��p�X�ٿ�OD:���@�4<
 4@��[��!?�qY�+�@�1X�ٿ5��=���@.��'
 4@��L$��!?B��\�+�@�4c�ٿ�'�<���@m��	 4@�.X^��!?��V�+�@�+�e�ٿԠ6���@�C�	 4@:��e��!?��XS�+�@�+�e�ٿԠ6���@�C�	 4@:��e��!?��XS�+�@�+�e�ٿԠ6���@�C�	 4@:��e��!?��XS�+�@�+�e�ٿԠ6���@�C�	 4@:��e��!?��XS�+�@��Q%^�ٿ���4���@���	 4@N0�h��!?��Q�+�@�[r�ٿ/�4���@s�g 4@"�ǐ!?�{M�+�@�[r�ٿ/�4���@s�g 4@"�ǐ!?�{M�+�@A��x�ٿ��m5���@]+�E 4@��Ӑ!?O�R�+�@V�'u�ٿIe�-���@��  4@���Ɛ!?O6AU�+�@��@�f�ٿ:�;���@�索	 4@�i	Uܐ!?q �Z�+�@��@�f�ٿ:�;���@�索	 4@�i	Uܐ!?q �Z�+�@��@�f�ٿ:�;���@�索	 4@�i	Uܐ!?q �Z�+�@��yy�ٿ �?@���@�Ŕ 4@L���!?�	W�+�@Vm��w�ٿ���:���@Y#�� 4@�)N��!?�^T�+�@̾{j��ٿcŬ@���@sW�i 4@���!?��Q�+�@?�[B��ٿǄK���@���) 4@������!?�^DM�+�@?�[B��ٿǄK���@���) 4@������!?�^DM�+�@�)걮�ٿ�gIG���@�/�� 4@�ė��!?,�
L�+�@_�s}��ٿږ�D���@���� 4@!��Ր!?r��S�+�@+�t.��ٿ���G���@�d 4@3����!?P�U�+�@��y��ٿ��P���@��� 4@�AЗ�!?萞R�+�@:����ٿ=�EN���@��u 4@���!?�ӌO�+�@w��_��ٿ~z�[���@���� 4@Cd,k��!?�P9M�+�@������ٿ�f�Q���@5�@� 4@�u����!?��R�+�@�s�n��ٿ��O���@��47 4@L�\��!?_�S�+�@�p�D��ٿ��Q���@��� 4@$�aŐ!?���T�+�@#y�$��ٿ�.�S���@�a� 4@ֻ򧅐!?:��T�+�@��x(��ٿ�8�\���@��� 4@��/���!?�6W�+�@�qϛ��ٿ�	h_���@Z�� 4@���p�!?]W�+�@oH(q��ٿhwb���@�|�� 4@�"����!?֟:S�+�@f�;���ٿO�Ja���@���� 4@5�rѐ!?)��R�+�@H�&ᣙٿY.hZ���@h��6 4@�ça��!?nDX�+�@G"U���ٿ.`U���@�b@ 4@lv�C#�!?��$W�+�@/�����ٿ&X���@Y%h. 4@��љǐ!?�%�R�+�@/�����ٿ&X���@Y%h. 4@��љǐ!?�%�R�+�@9#���ٿi*hO���@��R� 4@�#-���!?S�+�@�'֕��ٿy��a���@O� 4@�;9>��!?j>V�+�@�'֕��ٿy��a���@O� 4@�;9>��!?j>V�+�@g�vR��ٿX�c���@�f@� 4@�λΐ!?���V�+�@)�8@��ٿ��X���@7�Y 4@�VQȐ!?��2S�+�@�\���ٿ3�nV���@w1�� 4@��� �!?��R�+�@ԛJ��ٿjDX���@��# 4@7�@��!?e��N�+�@��z��ٿ�-N���@Y˿� 4@�n1� �!?�9DM�+�@���?��ٿ)�J���@�
�( 4@x�9�!?!9PO�+�@���?��ٿ)�J���@�
�( 4@x�9�!?!9PO�+�@E�Dٿ�U�B���@�9�� 4@���{�!?T�P�+�@a�TәٿhM[���@�kW 4@{S����!?�C�P�+�@a�TәٿhM[���@�kW 4@{S����!?�C�P�+�@�n��ٿ;M�f���@�+2e 4@���j`�!?#E�Q�+�@�,A�ߙٿ���f���@5U� 4@�5 �K�!?���R�+�@��ٿ�b���@�L� 4@�h��t�!?�2%P�+�@��ٿ�b���@�L� 4@�h��t�!?�2%P�+�@��ٿ�b���@�L� 4@�h��t�!?�2%P�+�@��ٿ�b���@�L� 4@�h��t�!?�2%P�+�@��ٿ�b���@�L� 4@�h��t�!?�2%P�+�@4���ٿS��l���@��8 4@�� �D�!?/��T�+�@4���ٿS��l���@��8 4@�� �D�!?/��T�+�@4���ٿS��l���@��8 4@�� �D�!?/��T�+�@�����ٿ:-v���@Q�M� 4@� g.�!?� T�+�@�����ٿ:-v���@Q�M� 4@� g.�!?� T�+�@�����ٿ:-v���@Q�M� 4@� g.�!?� T�+�@�?��ٿ��`}���@dw� 4@�����!?��|U�+�@{�5�͙ٿn�Mk���@O<� 4@A�W3��!?!�V�+�@{�5�͙ٿn�Mk���@O<� 4@A�W3��!?!�V�+�@��~�ٿ��(n���@H�� 4@953�W�!?p�=[�+�@	#�7��ٿ�><d���@��� 4@ٴ����!?�!�_�+�@	#�7��ٿ�><d���@��� 4@ٴ����!?�!�_�+�@va�K�ٿ�h�G���@QJ�	 4@���!?#a�+�@�V�Y��ٿ_m�Q���@��	� 4@� ����!?NI]�+�@�V�Y��ٿ_m�Q���@��	� 4@� ����!?NI]�+�@]�F��ٿ��7\���@��h 4@��Ӳϐ!?d��]�+�@���j}�ٿ���S���@�s� 4@s��!?��0h�+�@W�L�@�ٿ�56@���@_2�(	 4@��
w�!?��:f�+�@�"B�ޘٿa
����@��sX 4@(?���!?g�Kk�+�@�"B�ޘٿa
����@��sX 4@(?���!?g�Kk�+�@e�.��ٿ0E����@7n�� 4@+�ˬ��!?��zi�+�@&)�Ęٿ��O���@i�� 4@�-��Ȑ!?���o�+�@�_L�˘ٿP ����@�� � 4@���b�!?�� o�+�@�k��ۘٿC+���@@� 4@:6��F�!?��p�+�@�k��ۘٿC+���@@� 4@:6��F�!?��p�+�@�k��ۘٿC+���@@� 4@:6��F�!?��p�+�@����ٿ������@^�+H 4@�����!?dKLu�+�@����ٿ������@^�+H 4@�����!?dKLu�+�@�oټH�ٿ,������@N��^ 4@��~;��!?�	��+�@�oټH�ٿ,������@N��^ 4@��~;��!?�	��+�@�oټH�ٿ,������@N��^ 4@��~;��!?�	��+�@UD�@u�ٿ�ȏ����@Vkϊ 4@�(^W��!?�؃�+�@p��z\�ٿf�u����@�	�� 4@�s�q�!?�j3��+�@p��z\�ٿf�u����@�	�� 4@�s�q�!?�j3��+�@H@*\��ٿ#����@���? 4@�ay'��!?�@(|�+�@���ٿ�m����@��' 4@�G���!?3V���+�@x$�֗ٿ�s�����@Ĺ�� 4@�G�ͅ�!?�@-��+�@B���p�ٿ3�����@��N 4@!]�⊐!?ͦ�v�+�@B���p�ٿ3�����@��N 4@!]�⊐!?ͦ�v�+�@B���p�ٿ3�����@��N 4@!]�⊐!?ͦ�v�+�@�� � �ٿ�)�����@ޘ� 4@�Ҋ�~�!?�x�+�@�;��\�ٿ@������@=E� 4@��6]�!?�ͯ��+�@�1�i
�ٿ!�q���@�`�� 4@�Ktb�!?6+I��+�@��p��ٿ�������@ +�� 4@������!?�=7��+�@�`S�;�ٿ�=�e���@��� 4@g�;ϐ!?��ǌ�+�@�`S�;�ٿ�=�e���@��� 4@g�;ϐ!?��ǌ�+�@�FU,l�ٿ�����@Zð 4@`p�3�!?��6��+�@�W#ѕٿ)%7����@��E�  4@Ć�qO�!?�O��+�@�W#ѕٿ)%7����@��E�  4@Ć�qO�!?�O��+�@��'��ٿD�����@ s�! 4@Y[�i�!?����+�@#�u���ٿ"�N����@�C�' 4@���?�!?F5��+�@�h�(�ٿX<b���@�+�� 4@7��)��!?�iG��+�@�h�(�ٿX<b���@�+�� 4@7��)��!?�iG��+�@ԓ-3��ٿ�H���@���0 4@��Ɛ!?J.���+�@�ܡؓٿ*��)���@��1�. 4@�Y���!?(���+�@�ܡؓٿ*��)���@��1�. 4@�Y���!?(���+�@Ng�Q�ٿ�C�U���@�A:u+ 4@�;e�!?����+�@Ng�Q�ٿ�C�U���@�A:u+ 4@�;e�!?����+�@Ng�Q�ٿ�C�U���@�A:u+ 4@�;e�!?����+�@Ng�Q�ٿ�C�U���@�A:u+ 4@�;e�!?����+�@��_�ٿ1+����@����& 4@n-��!?pC*��+�@>�����ٿӄYx���@@�@+ 4@逘!�!?JO���+�@>�����ٿӄYx���@@�@+ 4@逘!�!?JO���+�@����t�ٿk�2���@ט�X 4@G$GS��!?�:��+�@����t�ٿk�2���@ט�X 4@G$GS��!?�:��+�@W��XƖٿ�?zB���@]��< 4@���ʐ!?oF'��+�@W��XƖٿ�?zB���@]��< 4@���ʐ!?oF'��+�@W��XƖٿ�?zB���@]��< 4@���ʐ!?oF'��+�@PNx�Q�ٿ��w���@�� 4@-����!?C���+�@PNx�Q�ٿ��w���@�� 4@-����!?C���+�@F��I�ٿR���@F� 4@�M���!?M�g��+�@���Ȗٿ�.]1���@��� 4@���o��!?0�Ğ�+�@���Ȗٿ�.]1���@��� 4@���o��!?0�Ğ�+�@�Mx� �ٿ&�����@2�h& 4@7#���!?�g ��+�@�ʁ��ٿ�j����@u�% 4@2B<���!?6,ϴ�+�@�o��8�ٿH�����@$�{$ 4@ �d���!?��q��+�@��\�ٿ1;n����@�%ܲ2 4@-�$�!?K��+�@B�k6��ٿvF����@N��3 4@x#V��!?����+�@��D���ٿ�����@�30 4@�]�f�!??����+�@Lh�ZG�ٿ���1���@4=C? 4@��D�!?�^��+�@`�΁ٿ���G���@�=AQ 4@(�+��!?�!WV�+�@H	�7n�ٿ��U����@��\E 4@�CR/�!?.+�0�+�@H	�7n�ٿ��U����@��\E 4@�CR/�!?.+�0�+�@H	�7n�ٿ��U����@��\E 4@�CR/�!?.+�0�+�@H	�7n�ٿ��U����@��\E 4@�CR/�!?.+�0�+�@nKhߌٿ�;����@l#)�] 4@���2�!?��Q��+�@?�P�ٿ������@lŖ)^ 4@��.�!?����+�@�bǼ;�ٿ,�(T���@Ҁ�b 4@tpPA��!?Ba��+�@Z^�u�ٿ�طY���@���^ 4@��z��!?��t��+�@�tQzY�ٿ�����@�Wf� 4@�~c�ސ!?{�=�+�@��@�̅ٿp������@G�� 4@�C���!?�5Y�+�@��@�̅ٿp������@G�� 4@�C���!?�5Y�+�@��@�̅ٿp������@G�� 4@�C���!?�5Y�+�@�Fc�2�ٿ��ğ���@��� 4@x�c��!?��r]�+�@�Fc�2�ٿ��ğ���@��� 4@x�c��!?��r]�+�@NX4l��ٿ-�#���@�ZtM� 4@�{w�k�!?��{?�+�@NX4l��ٿ-�#���@�ZtM� 4@�{w�k�!?��{?�+�@NX4l��ٿ-�#���@�ZtM� 4@�{w�k�!?��{?�+�@�$��:�ٿ:�����@&f๰ 4@�⚵��!?Tu��+�@�$��:�ٿ:�����@&f๰ 4@�⚵��!?Tu��+�@��zTK�ٿa�$���@b��s 4@X�t
��!?�g���+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@���T]�ٿ$c���@LTΦr 4@.Rwr�!?�EX��+�@�7j�ٿ��>B���@J�_ 4@���㘐!?�db��+�@�7j�ٿ��>B���@J�_ 4@���㘐!?�db��+�@�7j�ٿ��>B���@J�_ 4@���㘐!?�db��+�@�7j�ٿ��>B���@J�_ 4@���㘐!?�db��+�@�7j�ٿ��>B���@J�_ 4@���㘐!?�db��+�@�C0ЊٿK[����@��;�k 4@g����!?7��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@H�;R��ٿ��
4���@p;�� 4@���!?�|��+�@�L=��ٿAV�����@����� 4@��u���!?xlI��+�@�L=��ٿAV�����@����� 4@��u���!?xlI��+�@�a�
߂ٿ�>����@��V�� 4@"�U���!?�Z���+�@����Ҋٿ�b����@��l 4@���Ґ!?-Ծ�+�@����Ҋٿ�b����@��l 4@���Ґ!?-Ծ�+�@��s^<�ٿ�W#����@��"z� 4@�F�א!?!A���+�@��s^<�ٿ�W#����@��"z� 4@�F�א!?!A���+�@��s^<�ٿ�W#����@��"z� 4@�F�א!?!A���+�@��s^<�ٿ�W#����@��"z� 4@�F�א!?!A���+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@wgL$�ٿ�
����@c���i 4@�{P؇�!?��Ҷ�+�@����d�ٿ���U���@��H_ 4@\�q_m�!?/v���+�@�\>nl�ٿ�?����@W�U� 4@�3Ca`�!?���+�@)v����ٿ�%~���@��Iij 4@�^n�!?0e���+�@)v����ٿ�%~���@��Iij 4@�^n�!?0e���+�@��0�ٿ)H�����@U�Ã 4@��ɐ!?3��+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@w�MIɇٿû�����@�e҄ 4@�i[�!?K�b.�+�@v@�ٿ�������@�Y�� 4@��=]Ɛ!?�z��+�@v@�ٿ�������@�Y�� 4@��=]Ɛ!?�z��+�@v@�ٿ�������@�Y�� 4@��=]Ɛ!?�z��+�@v@�ٿ�������@�Y�� 4@��=]Ɛ!?�z��+�@Xf�Y�ٿ)z9���@V�>L� 4@�����!?Y%o��+�@'�q�ʊٿ�yq���@�Hv 4@��y�!?�7���+�@'�q�ʊٿ�yq���@�Hv 4@��y�!?�7���+�@'�q�ʊٿ�yq���@�Hv 4@��y�!?�7���+�@'�q�ʊٿ�yq���@�Hv 4@��y�!?�7���+�@�X�ۃٿ4_Up���@��V/� 4@�?|���!?��\��+�@�C��ٿ�1�~���@%��u� 4@_��?̐!?��g��+�@��0��ٿ��Y���@����� 4@:��}ǐ!?�&��+�@3�CvK�ٿ�Zg����@#kG�y 4@�q���!?�D�+�@�A�ҍٿ������@QlP�m 4@�M�ې!?Bo8��+�@�A�ҍٿ������@QlP�m 4@�M�ې!?Bo8��+�@�%���}ٿ���"���@��qz� 4@��U��!?3�JR�+�@�n���{ٿLo+A��@R� � 4@�����!? >{[�+�@���H&xٿ�N	��@���� 4@��wo	�!?5	���+�@�`�sٿJ���@6��4@�9!	�!?����+�@k�+RPvٿ�;TH��@�'�4@t�Z7��!?E4���+�@�cyw�wٿz8���@���4@��Cm��!?f�/�+�@hƜM�|ٿO�r����@��%� 4@�.`�z�!?4�<��+�@hƜM�|ٿO�r����@��%� 4@�.`�z�!?4�<��+�@Vm ���ٿ��)���@���� 4@)1�b�!?���+�@���5�ٿ4��{���@Y!�I� 4@�]�A�!?ʤt8�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@#�á�ٿ������@�\�)� 4@B%sa�!?ӻt'�+�@�|��׌ٿE��w���@�{��y 4@��>���!?�����+�@�|��׌ٿE��w���@�{��y 4@��>���!?�����+�@,�Ԙ�ٿ��E���@*��� 4@�,XH�!?�E�I�+�@,�Ԙ�ٿ��E���@*��� 4@�,XH�!?�E�I�+�@��I��ٿY}s2���@jᭃ 4@��$\�!?��2,�+�@��I��ٿY}s2���@jᭃ 4@��$\�!?��2,�+�@��I��ٿY}s2���@jᭃ 4@��$\�!?��2,�+�@��I��ٿY}s2���@jᭃ 4@��$\�!?��2,�+�@��I��ٿY}s2���@jᭃ 4@��$\�!?��2,�+�@��T�ٿ�/����@
�\� 4@��&���!?��4�+�@��T�ٿ�/����@
�\� 4@��&���!?��4�+�@��T�ٿ�/����@
�\� 4@��&���!?��4�+�@��$[�ٿ�:����@ ۽� 4@'�!翐!?ur�-�+�@-³�
�ٿ	Z�!���@l��pD 4@�O_X�!?�u.!�+�@-³�
�ٿ	Z�!���@l��pD 4@�O_X�!?�u.!�+�@-³�
�ٿ	Z�!���@l��pD 4@�O_X�!?�u.!�+�@-³�
�ٿ	Z�!���@l��pD 4@�O_X�!?�u.!�+�@s�/e�ٿ�:�I���@7=��� 4@��h��!?�c��+�@s�/e�ٿ�:�I���@7=��� 4@��h��!?�c��+�@s�/e�ٿ�:�I���@7=��� 4@��h��!?�c��+�@ԁ�҄ٿ�ZO����@�P�G� 4@�"Z��!?OZXc�+�@ԁ�҄ٿ�ZO����@�P�G� 4@�"Z��!?OZXc�+�@��G;��ٿ�n���@�h5� 4@:��μ�!?��g�+�@|��<�ٿ�v����@]��i� 4@�(��!? ����+�@|��<�ٿ�v����@]��i� 4@�(��!? ����+�@d���ٿ�o�y���@�0�� 4@D'�א!?��)�+�@C�J{��ٿ�����@��Dљ 4@e/ Ő!?��[7�+�@C�J{��ٿ�����@��Dљ 4@e/ Ő!?��[7�+�@AΉ��ٿ5|���@�
G�4@������!?��{��+�@�r�戀ٿT!Η���@j9K� 4@��H���!?�7�b�+�@�p��ٿ�vy-���@x�9Բ 4@��ܐ!?���+�@�p��ٿ�vy-���@x�9Բ 4@��ܐ!?���+�@�p��ٿ�vy-���@x�9Բ 4@��ܐ!?���+�@�p��ٿ�vy-���@x�9Բ 4@��ܐ!?���+�@�p��ٿ�vy-���@x�9Բ 4@��ܐ!?���+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@�o𞏄ٿ8p����@s��� 4@���ᤐ!?k��:�+�@=�d��ٿ@7����@��D�� 4@���ފ�!?�@��+�@=�d��ٿ@7����@��D�� 4@���ފ�!?�@��+�@y���ٿ�����@�M�t� 4@����֐!?�zD�+�@*�I�ٿp�{���@`�@�� 4@K\7���!?��2��+�@��m�ٿ�	۰���@t�*�O 4@M�U��!?�r# �+�@��m�ٿ�	۰���@t�*�O 4@M�U��!?�r# �+�@(	=���ٿȠ�����@�8�uq 4@vD#Ǧ�!?��c_�+�@(	=���ٿȠ�����@�8�uq 4@vD#Ǧ�!?��c_�+�@�;��jٿ��~d���@V��� 4@!��{��!?��B��+�@�Ld��ٿ�5����@ě�� 4@��wА!?|O���+�@SHm�P�ٿp�}���@@3a4@�����!?yAB��+�@SHm�P�ٿp�}���@@3a4@�����!?yAB��+�@�N�P��ٿ~����@�F�u�4@=�<d�!?�M6�+�@���5>�ٿ������@�E<�,4@�ɵ:�!?E�΀�+�@���5>�ٿ������@�E<�,4@�ɵ:�!?E�΀�+�@���5>�ٿ������@�E<�,4@�ɵ:�!?E�΀�+�@���5>�ٿ������@�E<�,4@�ɵ:�!?E�΀�+�@���5>�ٿ������@�E<�,4@�ɵ:�!?E�΀�+�@a%\5��ٿ,�@Y���@�L�_4@lw:�!?�j�J�+�@a%\5��ٿ,�@Y���@�L�_4@lw:�!?�j�J�+�@a%\5��ٿ,�@Y���@�L�_4@lw:�!?�j�J�+�@a%\5��ٿ,�@Y���@�L�_4@lw:�!?�j�J�+�@���ٿO��e���@2[��� 4@4����!?[����+�@�q0#��ٿG����@i:h6� 4@��c9��!?���+�@�q0#��ٿG����@i:h6� 4@��c9��!?���+�@'�����ٿa�j����@�sL��3@�_���!?�$c��+�@'�����ٿa�j����@�sL��3@�_���!?�$c��+�@_���I�ٿ�����@�i��g 4@�"B�!?����+�@;�\s��ٿ�.���@����8 4@��.4��!?� ��+�@)�L�)�ٿ������@2J�#4@g`J��!?�����+�@)�L�)�ٿ������@2J�#4@g`J��!?�����+�@)�L�)�ٿ������@2J�#4@g`J��!?�����+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�*�L2�ٿ�d:����@���0� 4@f"߳Đ!?(�F��+�@�%�ދ�ٿ//�O���@Q���� 4@��&��!?_��+�@�%�ދ�ٿ//�O���@Q���� 4@��&��!?_��+�@�%�ދ�ٿ//�O���@Q���� 4@��&��!?_��+�@������ٿ:+4-���@����� 4@>�P�ϐ!?л�/�+�@qf�d@�ٿ0����@4�SH� 4@���ʐ!?Q��j�+�@��:P1�ٿK]5� ��@P���4@=�aʐ!?8-���+�@��:P1�ٿK]5� ��@P���4@=�aʐ!?8-���+�@��:P1�ٿK]5� ��@P���4@=�aʐ!?8-���+�@e��gR�ٿ�^����@@ �~ 4@�<̈́��!?���K�+�@��,���ٿ��1���@Db&D4@bl$��!?��#�+�@��,���ٿ��1���@Db&D4@bl$��!?��#�+�@��,���ٿ��1���@Db&D4@bl$��!?��#�+�@��,���ٿ��1���@Db&D4@bl$��!?��#�+�@��,���ٿ��1���@Db&D4@bl$��!?��#�+�@���/�ٿ���@0P��4@1�0Ð!?�Z��+�@���/�ٿ���@0P��4@1�0Ð!?�Z��+�@���;3�ٿ>�a��@����4@�,����!?Hۡ��+�@���;3�ٿ>�a��@����4@�,����!?Hۡ��+�@���;3�ٿ>�a��@����4@�,����!?Hۡ��+�@���;3�ٿ>�a��@����4@�,����!?Hۡ��+�@1u8␇ٿ%~����@k�W5j4@Om�b�!?����+�@1u8␇ٿ%~����@k�W5j4@Om�b�!?����+�@1u8␇ٿ%~����@k�W5j4@Om�b�!?����+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@��f�ٿ��/���@�p���4@��*�T�!?z�h��+�@����ٿd`�!��@T/��4@1XQ"��!?�)�+�@��pe!�ٿ9��@+�*+24@*3f�!?����+�@퉯�ٿN����@�%$ZX4@BB���!?�:x�+�@l�iiυٿ趦���@M���V4@|�՝�!?6�@�+�@l�iiυٿ趦���@M���V4@|�՝�!?6�@�+�@e��=�ٿM� w%��@�}m3g4@�v� ��!?��@+�+�@e��=�ٿM� w%��@�}m3g4@�v� ��!?��@+�+�@e��=�ٿM� w%��@�}m3g4@�v� ��!?��@+�+�@e��=�ٿM� w%��@�}m3g4@�v� ��!?��@+�+�@e��=�ٿM� w%��@�}m3g4@�v� ��!?��@+�+�@$�X?�ٿ�q�z��@n�'4@5��C��!?��W��+�@$�X?�ٿ�q�z��@n�'4@5��C��!?��W��+�@$�X?�ٿ�q�z��@n�'4@5��C��!?��W��+�@$�X?�ٿ�q�z��@n�'4@5��C��!?��W��+�@���{�ٿ]ב/��@Y��(4@$��͐!?����+�@���{�ٿ]ב/��@Y��(4@$��͐!?����+�@���{�ٿ]ב/��@Y��(4@$��͐!?����+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@25A��ٿNO�*4��@�4���4@,f(袐!?�&���+�@��{F��ٿ.���@�v��4@)g�+	�!?�����+�@��{F��ٿ.���@�v��4@)g�+	�!?�����+�@�MIe��ٿ�Z���@��J=4@G����!?	?�U�+�@�MIe��ٿ�Z���@��J=4@G����!?	?�U�+�@�MIe��ٿ�Z���@��J=4@G����!?	?�U�+�@��Q��ٿ�A���@�5�G4@�x�ݐ!?�2_��+�@��Q��ٿ�A���@�5�G4@�x�ݐ!?�2_��+�@-�.;H�ٿ$#8���@b�n�4@�����!?ъ�+�@-�.;H�ٿ$#8���@b�n�4@�����!?ъ�+�@-�.;H�ٿ$#8���@b�n�4@�����!?ъ�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@ʂ"�(ٿ�^���@�M���4@�@Q���!?�u�8�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@��"��ٿ}��l*��@xW�4@��dݐ!?��B�+�@����ٿd=,C��@"�I=�4@fDW��!?"�Q9�+�@����ٿd=,C��@"�I=�4@fDW��!?"�Q9�+�@�N���ٿ��O��@���:4@��ِ!?V���+�@�N���ٿ��O��@���:4@��ِ!?V���+�@�N���ٿ��O��@���:4@��ِ!?V���+�@Q�I�ٿd� ��@�Łq4@�U�/��!?�4��+�@Q�I�ٿd� ��@�Łq4@�U�/��!?�4��+�@Q�I�ٿd� ��@�Łq4@�U�/��!?�4��+�@Q�I�ٿd� ��@�Łq4@�U�/��!?�4��+�@�)��ٿ]�r&��@=��9{4@����ݐ!?�* w�+�@�)��ٿ]�r&��@=��9{4@����ݐ!?�* w�+�@�)��ٿ]�r&��@=��9{4@����ݐ!?�* w�+�@���<I�ٿ[Qj:��@����4@����!?M��+�@�x�)��ٿ7�|q��@�f�k4@�+�{�!?�95��+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@��0�ٿr�H��@wys(l
4@w@��!?z%K�+�@�JUw��ٿ�,�K2��@2��*4@5���!?+�3��+�@�JUw��ٿ�,�K2��@2��*4@5���!?+�3��+�@��RU��ٿ����5��@��s�F	4@(~�-��!?�@��+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�$(}ٿ5�!O��@	��m4@��Uΐ!?]�e�+�@�0ӂx�ٿ�C� 2��@~�Ee64@ρe~�!?	��+�@Zb��݁ٿ⥇j!��@���g4@+���!?.��+�@�	_O�ٿ7��7��@�yPK	4@�l�ț�!?�W�P�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@	5~�y�ٿ:����@1��-c4@�:m��!?�yJ�+�@��*�ٿMT;����@�`Y34@}�4��!?�f���+�@��*�ٿMT;����@�`Y34@}�4��!?�f���+�@��nt�ٿ !�Z��@�8bO�4@KJ2���!?/�v�+�@��nt�ٿ !�Z��@�8bO�4@KJ2���!?/�v�+�@��nt�ٿ !�Z��@�8bO�4@KJ2���!?/�v�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@��A�wٿ�����@ev�\q4@���ڐ!?BR�+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@+�ܗ��ٿ�-���@�BN4@Ռ�'��!?��+�@Q�UN�ٿ�eb2��@��Z��4@_�ŋ�!?��+�@Q�UN�ٿ�eb2��@��Z��4@_�ŋ�!?��+�@Q�UN�ٿ�eb2��@��Z��4@_�ŋ�!?��+�@����ٿ���@2f���3@Y����!?b��k�+�@����ٿ���@2f���3@Y����!?b��k�+�@����ٿ���@2f���3@Y����!?b��k�+�@���ӵ�ٿ;�3�ۇ�@Ǭ� 4@9U���!?^`@x�+�@����ٿ( q���@I"�)4@,
C��!?un���+�@����ٿ( q���@I"�)4@,
C��!?un���+�@$�?ʇٿ��6Z��@���u$4@3��!?{C��+�@�!�<O�ٿF�2��@A�_�4@��1�!?v�D|�+�@�!�<O�ٿF�2��@A�_�4@��1�!?v�D|�+�@�!�<O�ٿF�2��@A�_�4@��1�!?v�D|�+�@&y�Ѐٿ�b4��@Z�?�4@ۑ;6�!?r��F�+�@�{��`�ٿ��-�*��@,�\4@����!?y���+�@�{��`�ٿ��-�*��@,�\4@����!?y���+�@�{��`�ٿ��-�*��@,�\4@����!?y���+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@���ٿr�43��@�XVDT4@��B��!?�@B��+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@6QWY:�ٿ�5n���@a�D4@�P�G�!?�#���+�@5��k�|ٿT�����@s/<l4@�_��!?�U�+�@�Ә�}ٿ�
��ч�@2O�:�4@����!?���6�+�@�Ә�}ٿ�
��ч�@2O�:�4@����!?���6�+�@�Ә�}ٿ�
��ч�@2O�:�4@����!?���6�+�@�Ә�}ٿ�
��ч�@2O�:�4@����!?���6�+�@�Ә�}ٿ�
��ч�@2O�:�4@����!?���6�+�@8����zٿ�f-f���@(��4@���ː!?�i�ة+�@8����zٿ�f-f���@(��4@���ː!?�i�ة+�@���~�ٿ:�����@��1�	4@"9u~�!?�ݱ+�@�DӸB�ٿ5U����@'�`��4@�`sH��!?!p�+�@�DӸB�ٿ5U����@'�`��4@�`sH��!?!p�+�@�DӸB�ٿ5U����@'�`��4@�`sH��!?!p�+�@�DӸB�ٿ5U����@'�`��4@�`sH��!?!p�+�@R��{ٿ�h��u��@"�;�64@*����!? ��o+�@;���jٿ�����@U?=a�4@w_����!?��37�+�@;���jٿ�����@U?=a�4@w_����!?��37�+�@���&ٿ�V �@jb��	4@�m�ؐ!?�=��d+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@m�q�ٿ��Չ���@
���4@�7����!?M;�Wh+�@Ez��/�ٿ}��!���@�B�4@}�&��!?��"}�+�@P67�ٿ������@vs�4@d���!?���s�+�@P67�ٿ������@vs�4@d���!?���s�+�@P67�ٿ������@vs�4@d���!?���s�+�@P67�ٿ������@vs�4@d���!?���s�+�@�~m�W�ٿ� ��:��@�B6�4@�d��!?�8�{;+�@�~m�W�ٿ� ��:��@�B6�4@�d��!?�8�{;+�@�~m�W�ٿ� ��:��@�B6�4@�d��!?�8�{;+�@�~m�W�ٿ� ��:��@�B6�4@�d��!?�8�{;+�@�~m�W�ٿ� ��:��@�B6�4@�d��!?�8�{;+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@W���ٿ"�wj��@:�>�\4@�w�!?Pj8�h+�@���t��ٿ�$�(r��@J�=o4@)��=��!?JͿ�\+�@Q>=��ٿ��|���@�S+684@�C���!?9�-�+�@Q>=��ٿ��|���@�S+684@�C���!?9�-�+�@Q>=��ٿ��|���@�S+684@�C���!?9�-�+�@�1��ٿ�S����@��p�C	4@F�ߴ�!? �:�+�@�1��ٿ�S����@��p�C	4@F�ߴ�!? �:�+�@�1��ٿ�S����@��p�C	4@F�ߴ�!? �:�+�@����ٿJ~�ѧ��@�:�K4@�9�g��!?
��N,�@y�2T|ٿ�Z��ڈ�@g�S�M	4@n�W��!?S�kr,�@y�2T|ٿ�Z��ڈ�@g�S�M	4@n�W��!?S�kr,�@ ����ٿp����@?��4@��1���!?�C�f,�@ ����ٿp����@?��4@��1���!?�C�f,�@ ����ٿp����@?��4@��1���!?�C�f,�@ ����ٿp����@?��4@��1���!?�C�f,�@ ����ٿp����@?��4@��1���!?�C�f,�@O�t�ٿ�IU���@0��|�4@���Ő!?A�J��+�@O�t�ٿ�IU���@0��|�4@���Ő!?A�J��+�@]ʹ�ˏٿ�&�%(��@~f��14@#te��!?O��
�,�@]ʹ�ˏٿ�&�%(��@~f��14@#te��!?O��
�,�@뛉�_�ٿ��u��@z@�	4@,�-��!?��u,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@ ��B+�ٿ�Lêb��@����4@��m��!?����,�@�%~�R}ٿ<Q����@��<�4@?X<iܐ!?E��Uf-�@�%~�R}ٿ<Q����@��<�4@?X<iܐ!?E��Uf-�@��C0�ٿD�'X���@���4@Ha��!?�'X6V,�@��C0�ٿD�'X���@���4@Ha��!?�'X6V,�@��C0�ٿD�'X���@���4@Ha��!?�'X6V,�@��C0�ٿD�'X���@���4@Ha��!?�'X6V,�@�$`�ٿ��n�ԉ�@���;4@�*���!?F�A-�@�$`�ٿ��n�ԉ�@���;4@�*���!?F�A-�@�$`�ٿ��n�ԉ�@���;4@�*���!?F�A-�@�$`�ٿ��n�ԉ�@���;4@�*���!?F�A-�@�$`�ٿ��n�ԉ�@���;4@�*���!?F�A-�@JRd�ٿx��D��@QM�A.4@��Ѿ�!?�Ba��-�@JRd�ٿx��D��@QM�A.4@��Ѿ�!?�Ba��-�@JRd�ٿx��D��@QM�A.4@��Ѿ�!?�Ba��-�@�L ⴏٿp��QO��@]��\4@�a��ɐ!?�� ,�@ʙ�do�ٿ(1����@��Qb4@��9���!?��0&f,�@ʙ�do�ٿ(1����@��Qb4@��9���!?��0&f,�@_̌��ٿ����1��@ץ�.	4@"}nm9�!?���,�@W���ؑٿ�pbw|��@r�h4@[8Y�!?a�s�\+�@W���ؑٿ�pbw|��@r�h4@[8Y�!?a�s�\+�@W���ؑٿ�pbw|��@r�h4@[8Y�!?a�s�\+�@��[؂ٿ�Yzr��@��\4@Q�|��!?�
U�j+�@��[؂ٿ�Yzr��@��\4@Q�|��!?�
U�j+�@��[؂ٿ�Yzr��@��\4@Q�|��!?�
U�j+�@��[؂ٿ�Yzr��@��\4@Q�|��!?�
U�j+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@�tC��ٿ�*U���@Y�OJ34@��ӥ�!?�K바+�@K�U�/�ٿ�&�(���@�w�&4@2����!?����*�@K�U�/�ٿ�&�(���@�w�&4@2����!?����*�@K�U�/�ٿ�&�(���@�w�&4@2����!?����*�@K�U�/�ٿ�&�(���@�w�&4@2����!?����*�@�@���ٿ4-bV���@��s�(�3@}����!?�|Lۥ+�@�@���ٿ4-bV���@��s�(�3@}����!?�|Lۥ+�@�@���ٿ4-bV���@��s�(�3@}����!?�|Lۥ+�@�@���ٿ4-bV���@��s�(�3@}����!?�|Lۥ+�@���r�ٿX�p��@�c��3@&���!?�\��-�@���r�ٿX�p��@�c��3@&���!?�\��-�@��RTFٿR3m���@R��W4@�Vn�!?��6��.�@��RTFٿR3m���@R��W4@�Vn�!?��6��.�@��RTFٿR3m���@R��W4@�Vn�!?��6��.�@��RTFٿR3m���@R��W4@�Vn�!?��6��.�@�{#Ɇٿ|�
Id��@b��t4@FmKҐ!?=�Ӄ.�@�{#Ɇٿ|�
Id��@b��t4@FmKҐ!?=�Ӄ.�@�{#Ɇٿ|�
Id��@b��t4@FmKҐ!?=�Ӄ.�@�{#Ɇٿ|�
Id��@b��t4@FmKҐ!?=�Ӄ.�@֩�r�ٿ�FY�g��@���f�4@+�Sl��!?�@4C�/�@֩�r�ٿ�FY�g��@���f�4@+�Sl��!?�@4C�/�@֩�r�ٿ�FY�g��@���f�4@+�Sl��!?�@4C�/�@֩�r�ٿ�FY�g��@���f�4@+�Sl��!?�@4C�/�@֩�r�ٿ�FY�g��@���f�4@+�Sl��!?�@4C�/�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@�hέy�ٿ�Qʈ��@� �ء 4@Ɵ�}�!?���0�@"H�;��ٿ���Ш��@�fǛ4@�x��^�!?��.�W3�@"H�;��ٿ���Ш��@�fǛ4@�x��^�!?��.�W3�@"H�;��ٿ���Ш��@�fǛ4@�x��^�!?��.�W3�@"H�;��ٿ���Ш��@�fǛ4@�x��^�!?��.�W3�@�!�%k�ٿz��ő�@r��� 4@������!?E�X03�@�!�%k�ٿz��ő�@r��� 4@������!?E�X03�@�!�%k�ٿz��ő�@r��� 4@������!?E�X03�@�!�%k�ٿz��ő�@r��� 4@������!?E�X03�@>����ٿ����ƕ�@ce���4@!=E�!?��e��6�@�L��ٿ/����@�	�/ 4@ ����!?��h�3�@�L��ٿ/����@�	�/ 4@ ����!?��h�3�@�L��ٿ/����@�	�/ 4@ ����!?��h�3�@�L��ٿ/����@�	�/ 4@ ����!?��h�3�@�L��ٿ/����@�	�/ 4@ ����!?��h�3�@�[ζ�ٿj�ڽ��@�,�9�3@�m����!?���/`0�@�[ζ�ٿj�ڽ��@�,�9�3@�m����!?���/`0�@D���ƅٿ���ʑ�@͡��3@�j��!?&���3�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@كVAŉٿ�z\
;��@�ѽ4@����$�!?G��0�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@�+*Ǎٿ�d����@�|ES4@���%�!?x&��}7�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@K�}p�ٿ��ea��@F3[�+4@S�X���!?m�E��1�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@`��
�ٿ
O{A���@��D4@�Z��&�!?Sl��6�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@-�փٿ-�Ka?��@ى��4@0�v�!?f
_$Z<�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�����}ٿ���b��@wR�+�4@x��!?w�i�;�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�7w�Åٿ��	��@�SUDy4@�֟��!?��ť�,�@�l�юٿ;	�+��@+'�� 4@S��Ȑ!?�´�(�@�l�юٿ;	�+��@+'�� 4@S��Ȑ!?�´�(�@�l�юٿ;	�+��@+'�� 4@S��Ȑ!?�´�(�@�l�юٿ;	�+��@+'�� 4@S��Ȑ!?�´�(�@�l�юٿ;	�+��@+'�� 4@S��Ȑ!?�´�(�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@{G���{ٿ�
��D��@0Yr�E4@�Fw���!?�d5�A�@u�l`Vٿ��}����@9)�W^4@��&��!?H)P�2�@���{ٿ+'ܶx��@7ЬM�4@1��p�!?��V.�@���{ٿ+'ܶx��@7ЬM�4@1��p�!?��V.�@N���ٿ6?9QRr�@a|��4@��.��!?�v8a��@N���ٿ6?9QRr�@a|��4@��.��!?�v8a��@O+��r�ٿ�,~�@'�\54@��5�ǐ!?n3��#$�@O+��r�ٿ�,~�@'�\54@��5�ǐ!?n3��#$�@O+��r�ٿ�,~�@'�\54@��5�ǐ!?n3��#$�@��鿉ٿ/=8�^s�@�ɍ4@f�#�!?�Z����@��鿉ٿ/=8�^s�@�ɍ4@f�#�!?�Z����@��鿉ٿ/=8�^s�@�ɍ4@f�#�!?�Z����@��鿉ٿ/=8�^s�@�ɍ4@f�#�!?�Z����@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@Q�kS�ٿsP,�df�@�`�V�	4@qFâڐ!?ȈZ��@b+10ٿ�e��z�@�}zM		4@>�|�ǐ!?R��!�@b+10ٿ�e��z�@�}zM		4@>�|�ǐ!?R��!�@b+10ٿ�e��z�@�}zM		4@>�|�ǐ!?R��!�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@B����ٿ`�&��h�@:a��^4@�H�@�!?"��\�@cp��ގٿ�LV�@��� 4@��3�!?f��D��@cp��ގٿ�LV�@��� 4@��3�!?f��D��@8og���ٿ�[	�i�@A�dE4@�9���!?��&�@8og���ٿ�[	�i�@A�dE4@�9���!?��&�@8og���ٿ�[	�i�@A�dE4@�9���!?��&�@8og���ٿ�[	�i�@A�dE4@�9���!?��&�@��멕ٿ.T����@w�hv4@�h͏Ӑ!?9�i3���@��멕ٿ.T����@w�hv4@�h͏Ӑ!?9�i3���@��멕ٿ.T����@w�hv4@�h͏Ӑ!?9�i3���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@����ٿ��^į�@�kx��4@� R��!?}~Wp���@� ���ٿ�}`I���@���2_4@���8��!?mɶ(��@~�}f=�ٿu"�����@�Tq�g	4@ݫw�Y�!?B�f΁�@~�}f=�ٿu"�����@�Tq�g	4@ݫw�Y�!?B�f΁�@~�}f=�ٿu"�����@�Tq�g	4@ݫw�Y�!?B�f΁�@(σ�_�ٿ>��l��@�b���4@c�K���!?R�C^�b�@(σ�_�ٿ>��l��@�b���4@c�K���!?R�C^�b�@(σ�_�ٿ>��l��@�b���4@c�K���!?R�C^�b�@(σ�_�ٿ>��l��@�b���4@c�K���!?R�C^�b�@��|�~ٿ�� R��@K�� 4@8��R��!?��m_�@�APAقٿ4��˶�@���/]�3@*k_a��!?W{���@�����ٿRk�*��@�UW/Y4@��MM�!?�D�<И�@�����ٿRk�*��@�UW/Y4@��MM�!?�D�<И�@�����ٿRk�*��@�UW/Y4@��MM�!?�D�<И�@�����ٿRk�*��@�UW/Y4@��MM�!?�D�<И�@�����ٿRk�*��@�UW/Y4@��MM�!?�D�<И�@+��#��ٿ��FC,��@lĦ�4@S"��!?{��o��@+��#��ٿ��FC,��@lĦ�4@S"��!?{��o��@+��#��ٿ��FC,��@lĦ�4@S"��!?{��o��@+��#��ٿ��FC,��@lĦ�4@S"��!?{��o��@�b�e0�ٿ�k1���@E��T�3@Z�p���!?d��@�o蒃ٿ؍>)��@���4@��!��!?�ưg���@�o蒃ٿ؍>)��@���4@��!��!?�ưg���@�o蒃ٿ؍>)��@���4@��!��!?�ưg���@�o蒃ٿ؍>)��@���4@��!��!?�ưg���@��2"Q�ٿ�%����@ޥ@�w 4@���1��!?D�7>�a�@��2"Q�ٿ�%����@ޥ@�w 4@���1��!?D�7>�a�@��2"Q�ٿ�%����@ޥ@�w 4@���1��!?D�7>�a�@�g��ٿ��|��@t_h�4@��`=��!?Ґ���@�g��ٿ��|��@t_h�4@��`=��!?Ґ���@�g��ٿ��|��@t_h�4@��`=��!?Ґ���@�g��ٿ��|��@t_h�4@��`=��!?Ґ���@�����ٿ�j]h8�@ZVu4@&jL�!?]�a��@�����ٿ�j]h8�@ZVu4@&jL�!?]�a��@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@!�>��ٿΘ�!���@a�+<�4@@��(�!?R�����@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@ӧ$�|�ٿlN��{�@N\4@�a �!? 2�Z�@.Y�yٿp�Ё2��@PX6G�4@D�0&s�!?�3^��@.Y�yٿp�Ё2��@PX6G�4@D�0&s�!?�3^��@.Y�yٿp�Ё2��@PX6G�4@D�0&s�!?�3^��@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@%S=C�ٿr%��<��@�@��4@�W����!?խ�R���@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@d��X�ٿ����\�@ ��#�3@@M�ڐ!?�t\!C�@n�J�Z�ٿ�o�eq�@Ke�� 4@ۅi
��!?�>NS�@n�J�Z�ٿ�o�eq�@Ke�� 4@ۅi
��!?�>NS�@n�J�Z�ٿ�o�eq�@Ke�� 4@ۅi
��!?�>NS�@n�J�Z�ٿ�o�eq�@Ke�� 4@ۅi
��!?�>NS�@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@Wu�C��ٿ�<o��!�@ҥL� 4@ �W���!?s��@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�>�s��ٿs;>�ɿ�@�Rd�4@l9H�Ґ!?q����@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�֡%3�ٿ`�ٲ^+�@��B�3@C�F��!?�cٟ�@�ջl�ٿ��O���@�l�'��3@���~��!?I����@�ջl�ٿ��O���@�l�'��3@���~��!?I����@�ջl�ٿ��O���@�l�'��3@���~��!?I����@�ջl�ٿ��O���@�l�'��3@���~��!?I����@�ջl�ٿ��O���@�l�'��3@���~��!?I����@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@b��r��ٿE����N�@R��9+�3@A�%E�!?D�u�<8�@���i(�ٿZWد�@�c/4@�ܢ��!?�Ot����@���i(�ٿZWد�@�c/4@�ܢ��!?�Ot����@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@���-�ٿ�Ĥ7Q�@az�;�4@�p�4��!?g�ʶ��@E�R�ٿ������@�1y�f4@��1�ߐ!?){����@�q�͉ٿu��6��@kb��4@�a�z�!?����@�q�͉ٿu��6��@kb��4@�a�z�!?����@x�C��ٿB����@z����4@�g��!?��sy���@x�C��ٿB����@z����4@�g��!?��sy���@x�C��ٿB����@z����4@�g��!?��sy���@��qP~ٿ��c�,@�@A��4@���FU�!?�i9��,�@�C"xٿe�[�6��@Z+��4@R��^�!?�)1ϛl�@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@_Oѵ�}ٿ<��S���@=^H �3@�c�E+�!?��͡��@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@x R+�ٿ��{�P��@
�z�4@{8�B�!?��~~�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�c�2�ٿ�' �i�@:��=�3@Xէ�!?f$n�L�@�Ҕ�A�ٿ��h��M�@�9�;~�3@u.�80�!?��|�47�@.���'�ٿ�5	�<��@�d6<��3@K��^�!?*S��]��@.���'�ٿ�5	�<��@�d6<��3@K��^�!?*S��]��@.���'�ٿ�5	�<��@�d6<��3@K��^�!?*S��]��@.���'�ٿ�5	�<��@�d6<��3@K��^�!?*S��]��@���ٿ�t�wA��@�,��3@�4CY\�!?K��,���@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@_�>3�ٿt�L�݊�@[�Ӗ4@�
��V�!?'��f�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�k%\�ٿ�R�\x��@bN��4@_xf�
�!?�P�m~�@�%�1�ٿ��.V��@Y���4@9ި,�!?�w)���@�%�1�ٿ��.V��@Y���4@9ި,�!?�w)���@�%�1�ٿ��.V��@Y���4@9ި,�!?�w)���@�%�1�ٿ��.V��@Y���4@9ި,�!?�w)���@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@�р)̅ٿ`:b�>b�@�C���3@��7ߐ!?��Qk>G�@��WA��ٿ��\Lkl�@��4�@ 4@VI���!?��ryO�@��WA��ٿ��\Lkl�@��4�@ 4@VI���!?��ryO�@��WA��ٿ��\Lkl�@��4�@ 4@VI���!?��ryO�@��WA��ٿ��\Lkl�@��4�@ 4@VI���!?��ryO�@��WA��ٿ��\Lkl�@��4�@ 4@VI���!?��ryO�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�lCp��ٿ�ώ�`�@���v� 4@>e�}!?�M*wF�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�˓�ٿ�^�z�@��4@���Ð!?�_¯Y�@�.uԈٿ�dHCJ�@nމ�4@���!?|,�'�4�@�.uԈٿ�dHCJ�@nމ�4@���!?|,�'�4�@�.uԈٿ�dHCJ�@nމ�4@���!?|,�'�4�@�.uԈٿ�dHCJ�@nމ�4@���!?|,�'�4�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@d�ЉB�ٿ��?��@�����4@ת�Ր!?�e�@�r�æ�ٿ�dj*H��@O�TQ4@!S���!?�4�`��@�g����ٿ[tb���@s\��4@5����!?6��r���@�g����ٿ[tb���@s\��4@5����!?6��r���@�g����ٿ[tb���@s\��4@5����!?6��r���@�g����ٿ[tb���@s\��4@5����!?6��r���@p�D��ٿ��m�_�@���S4@�+�-�!?���TE�@p�D��ٿ��m�_�@���S4@�+�-�!?���TE�@p�D��ٿ��m�_�@���S4@�+�-�!?���TE�@p�D��ٿ��m�_�@���S4@�+�-�!?���TE�@p�D��ٿ��m�_�@���S4@�+�-�!?���TE�@y���\�ٿ,��T���@0���3@&�2vI�!?-�O�D��@y���\�ٿ,��T���@0���3@&�2vI�!?-�O�D��@y���\�ٿ,��T���@0���3@&�2vI�!?-�O�D��@y���\�ٿ,��T���@0���3@&�2vI�!?-�O�D��@y���\�ٿ,��T���@0���3@&�2vI�!?-�O�D��@l��(b�ٿ^��_D��@E��% 4@��^_ِ!?뤲@���@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@��Vٗ�ٿ.�.��@l���4@��JӐ!?��rF��@�7���ٿ ��@��*H4@���*��!?B��:
�@����?�ٿ��ILw�@�/�K!4@!�͟��!?d���_��@����?�ٿ��ILw�@�/�K!4@!�͟��!?d���_��@����?�ٿ��ILw�@�/�K!4@!�͟��!?d���_��@����?�ٿ��ILw�@�/�K!4@!�͟��!?d���_��@����?�ٿ��ILw�@�/�K!4@!�͟��!?d���_��@���Z��ٿ�za6���@n�#@4@��n��!?����Z��@-�H�l�ٿy�e1�@�� �X4@�����!?S5��)!�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@J���ٿ�gn�<w�@���#4@�C��ݐ!?�a��W�@��n�ٿ���Wj�@l�X��3@��IĐ!?.�&�M�@��n�ٿ���Wj�@l�X��3@��IĐ!?.�&�M�@��n�ٿ���Wj�@l�X��3@��IĐ!?.�&�M�@��n�ٿ���Wj�@l�X��3@��IĐ!?.�&�M�@����h�ٿ���3��@��=�O4@NV��!?��6e��@����h�ٿ���3��@��=�O4@NV��!?��6e��@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@4;�Ђٿ8V$�ԇ�@�9�04@B=ۤ�!?�/Ƣ�d�@
妆;�ٿ�9�$��@�>܉�4@'����!?�N`�@
妆;�ٿ�9�$��@�>܉�4@'����!?�N`�@
妆;�ٿ�9�$��@�>܉�4@'����!?�N`�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@"�A�ٿ�"7m�:�@���4@��א!?U���(�@����ٿ5w����@Wa��4@h�|Ȑ!?�����@��eC[�ٿIj1����@	�&�t4@1��ِ!?����i�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�b{ț�ٿ�,��'D�@
]O�4@������!?<Ś�/�@�s`��ٿ"�B"�W�@Qҩ24@��p�̐!?\Ԁs>�@�s`��ٿ"�B"�W�@Qҩ24@��p�̐!?\Ԁs>�@��~�ٿr��$4�@���[4@RA�!?l����@��~�ٿr��$4�@���[4@RA�!?l����@��~�ٿr��$4�@���[4@RA�!?l����@��~�ٿr��$4�@���[4@RA�!?l����@C���]�ٿ��B�L�@�-v�4@��{dz�!?�m4�\6�@C���]�ٿ��B�L�@�-v�4@��{dz�!?�m4�\6�@ ��4��ٿt��G@��@;����4@�D���!?�*gz��@ ��4��ٿt��G@��@;����4@�D���!?�*gz��@�dRKR�ٿ5�4��4�@��i���3@Mz����!?��7XV#�@�dRKR�ٿ5�4��4�@��i���3@Mz����!?��7XV#�@�dRKR�ٿ5�4��4�@��i���3@Mz����!?��7XV#�@�dRKR�ٿ5�4��4�@��i���3@Mz����!?��7XV#�@nÂ�5�ٿ9+�FR�@23�<� 4@51%B��!?cebf�9�@>����ٿ|����@�v�Q� 4@ۋ�{y�!?��Ҕs	�@P�/�:�ٿ���<z��@ˮ�6�4@�Ʉ���!?~� ���@P�/�:�ٿ���<z��@ˮ�6�4@�Ʉ���!?~� ���@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@�)�Z�|ٿvE��@�@�!� =4@��a��!?F`y,�@���ٿ�Ғ�#�@v��4@z^��!?�[L�#�@��z�ٿ^I��"�@�0�I�4@�3��!?sN�Ҍ�@��z�ٿ^I��"�@�0�I�4@�3��!?sN�Ҍ�@F���ٿ�g=����@�V;,�4@��*_�!?[��Ɣ�@�%�ٿ��PK{��@�#Ҳ4@7߼ϐ!?�1�:��@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@���X|ٿ�j�`�@e�qH�4@�W��!?�ۀ�E�@�nֻ�ٿTj�*�K�@� ��4@�k���!?�δ�6�@������ٿ�J��k�@�1j04@�P��!?�1�1fN�@������ٿ�J��k�@�1j04@�P��!?�1�1fN�@Ĩ�!�ٿ�Fɇ�`�@Uό�4@�ץ�ؐ!?����EF�@Ĩ�!�ٿ�Fɇ�`�@Uό�4@�ץ�ؐ!?����EF�@Ĩ�!�ٿ�Fɇ�`�@Uό�4@�ץ�ؐ!?����EF�@5�U l�ٿ$T�|?�@jz�4@�b��!??��d�,�@5�U l�ٿ$T�|?�@jz�4@�b��!??��d�,�@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@�lυٿݾо���@ƞ�e4@�����!?��)o��@!z�_L�ٿ�����@��t]4@�:�Ӑ!?W��t�{�@!z�_L�ٿ�����@��t]4@�:�Ӑ!?W��t�{�@!z�_L�ٿ�����@��t]4@�:�Ӑ!?W��t�{�@!z�_L�ٿ�����@��t]4@�:�Ӑ!?W��t�{�@!z�_L�ٿ�����@��t]4@�:�Ӑ!?W��t�{�@ԡ�B�ٿrNMF�@ݘ��4@K��!?�`�n&1�@ԡ�B�ٿrNMF�@ݘ��4@K��!?�`�n&1�@ԡ�B�ٿrNMF�@ݘ��4@K��!?�`�n&1�@ԡ�B�ٿrNMF�@ݘ��4@K��!?�`�n&1�@ԡ�B�ٿrNMF�@ݘ��4@K��!?�`�n&1�@	�a�]�ٿ 7�0a�@Vz6�4@��L~��!?�xs��D�@	�a�]�ٿ 7�0a�@Vz6�4@��L~��!?�xs��D�@	�a�]�ٿ 7�0a�@Vz6�4@��L~��!?�xs��D�@	�a�]�ٿ 7�0a�@Vz6�4@��L~��!?�xs��D�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@�.�Fn�ٿ��m	�=�@1��K��3@u��5ɐ!?��a>)�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@����;�ٿ������@�(��N4@�\K�ʐ!?�;Њa�@�N�d�ٿ���W�@��_z4@�R����!?�f�i<�@{E���ٿuQO�I�@g;-4@AP�Ƕ�!?b�����@��DT�ٿ'"��7��@o���4@�3<��!?x�[��@��DT�ٿ'"��7��@o���4@�3<��!?x�[��@��DT�ٿ'"��7��@o���4@�3<��!?x�[��@��DT�ٿ'"��7��@o���4@�3<��!?x�[��@��?�ٿ'�����@=����3@�����!?\�����@��?�ٿ'�����@=����3@�����!?\�����@��?�ٿ'�����@=����3@�����!?\�����@�"X��ٿ^p��&N�@�$���4@�j�80�!?�W��{8�@��@�ٿ�6�0��@����I4@�����!?��S��x�@DM/$�ٿ��S#7�@.�)�4@�w%��!?5Ϗ�4%�@DM/$�ٿ��S#7�@.�)�4@�w%��!?5Ϗ�4%�@DM/$�ٿ��S#7�@.�)�4@�w%��!?5Ϗ�4%�@DM/$�ٿ��S#7�@.�)�4@�w%��!?5Ϗ�4%�@DM/$�ٿ��S#7�@.�)�4@�w%��!?5Ϗ�4%�@�(�^�ٿ��[K�@��a�'4@k u�!?��qϨ4�@�(�^�ٿ��[K�@��a�'4@k u�!?��qϨ4�@�(�^�ٿ��[K�@��a�'4@k u�!?��qϨ4�@�(�^�ٿ��[K�@��a�'4@k u�!?��qϨ4�@�(�^�ٿ��[K�@��a�'4@k u�!?��qϨ4�@[˵�U�ٿ�_�����@�ک� 4@�	'7ې!?([�Wy�@��ٿ�ևQ�r�@�%_�-4@K�^�!?C���Q�@=hԯ��ٿ��$���@M�ó� 4@�*����!?�{���k�@=hԯ��ٿ��$���@M�ó� 4@�*����!?�{���k�@=hԯ��ٿ��$���@M�ó� 4@�*����!?�{���k�@2\�V�ٿj�F���@�P�0�4@����!?KW�r��@f׭�ٿ�]�V�@}
�C�3@:����!?�I[\<�@f׭�ٿ�]�V�@}
�C�3@:����!?�I[\<�@f׭�ٿ�]�V�@}
�C�3@:����!?�I[\<�@���T-�ٿ�[@S��@{Yt� 4@>�'B��!?<mѰ���@���T-�ٿ�[@S��@{Yt� 4@>�'B��!?<mѰ���@.�Y���ٿ�5tF��@,���4@fne+�!?B�`�k��@���9�ٿLd8��X�@sM��4@������!?��C9�=�@]B���ٿH�$�i��@�W�Rq4@à�纐!?���`+w�@�m�5�ٿ�8#��f�@�d50A4@�1ʌ�!?V,=P�K�@�m�5�ٿ�8#��f�@�d50A4@�1ʌ�!?V,=P�K�@�m�5�ٿ�8#��f�@�d50A4@�1ʌ�!?V,=P�K�@�m�5�ٿ�8#��f�@�d50A4@�1ʌ�!?V,=P�K�@�m�5�ٿ�8#��f�@�d50A4@�1ʌ�!?V,=P�K�@~����ٿn\��x5�@��js?4@e.I�Ő!?*��yS#�@~����ٿn\��x5�@��js?4@e.I�Ő!?*��yS#�@~����ٿn\��x5�@��js?4@e.I�Ő!?*��yS#�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@��-�o�ٿ3_�!���@���m�4@�� Ґ!?pUsk�n�@�n.�n�ٿP_(H�o�@\�c&4@HXV�ߐ!?G-�N�@�n.�n�ٿP_(H�o�@\�c&4@HXV�ߐ!?G-�N�@����b�ٿ!��MZh�@Ů4@��9a}�!?J
:]�G�@����b�ٿ!��MZh�@Ů4@��9a}�!?J
:]�G�@����;�ٿJh
����@/51E4@�+���!?�z^l�@��!�ٿ����W�@_�)�4@��Tl��!?�%J^�6�@��!�ٿ����W�@_�)�4@��Tl��!?�%J^�6�@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@�2v�P�ٿ'������@����� 4@ēꀐ!?�����@K� D��ٿ��b�D�@��T4@��<x�!?�*i��"�@K� D��ٿ��b�D�@��T4@��<x�!?�*i��"�@K� D��ٿ��b�D�@��T4@��<x�!?�*i��"�@K� D��ٿ��b�D�@��T4@��<x�!?�*i��"�@K� D��ٿ��b�D�@��T4@��<x�!?�*i��"�@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@=͔/t�ٿ6Gq40�@����24@�-|��!?������@�:X�|ٿ�Y}��@9��P�4@S����!?�϶����@�:X�|ٿ�Y}��@9��P�4@S����!?�϶����@�:X�|ٿ�Y}��@9��P�4@S����!?�϶����@���2+�ٿͣ��mn�@��0$��3@�dW�!?48Ik�I�@���2+�ٿͣ��mn�@��0$��3@�dW�!?48Ik�I�@�N�yٿr���#�@����4@)��ī�!?-���H�@!��$�ٿ�*����@)Ţ0h�3@a���А!?��=���@6w��*�ٿRw0��@�;f4@?s�!?��@6w��*�ٿRw0��@�;f4@?s�!?��@6w��*�ٿRw0��@�;f4@?s�!?��@6w��*�ٿRw0��@�;f4@?s�!?��@�^\�ٿ�m�.Z=�@a���94@��v��!?:���,�@�^\�ٿ�m�.Z=�@a���94@��v��!?:���,�@�����ٿ��In�O�@��p��4@�����!?����@�@�����ٿ��In�O�@��p��4@�����!?����@�@�����ٿ��In�O�@��p��4@�����!?����@�@�����ٿ��In�O�@��p��4@�����!?����@�@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@��\J��ٿ�tY�\�@k���4@��`j�!?������@�~�䗈ٿ�g��3N�@WY��m4@�B�iP�!?y�NxH�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@O�^��ٿ�E�,Z�@c���4@rO^F��!?reA �G�@��-Q%�ٿd��t���@��i4@!u���!?����}�@��-Q%�ٿd��t���@��i4@!u���!?����}�@�[�z;~ٿp.uD�@��b��4@AE�ې!?�+�(+�@�[�z;~ٿp.uD�@��b��4@AE�ې!?�+�(+�@�[�z;~ٿp.uD�@��b��4@AE�ې!?�+�(+�@���
#�ٿʹ���@��4�. 4@UXMB�!?����<��@7  �Q�ٿ�ɐ��@�J���4@v���!?EG2V
�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@�S�`n�ٿA��L�@Zn�4@W$�V�!?�'!]�D�@?��P7�ٿg�H��@OJ�4@e��mŐ!?� �ZQ_�@?��P7�ٿg�H��@OJ�4@e��mŐ!?� �ZQ_�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I��fh�ٿ�4��p�@��9.4@�V��j�!?���S<�@I�L�;�ٿ#�̥�@aE�m4@��Hʐ!?�%*�
[�@I�L�;�ٿ#�̥�@aE�m4@��Hʐ!?�%*�
[�@I�L�;�ٿ#�̥�@aE�m4@��Hʐ!?�%*�
[�@I�L�;�ٿ#�̥�@aE�m4@��Hʐ!?�%*�
[�@���cj�ٿ1N~+��@P���&4@O\R��!?fp�U�@���cj�ٿ1N~+��@P���&4@O\R��!?fp�U�@���cj�ٿ1N~+��@P���&4@O\R��!?fp�U�@�!T�M�ٿ+�*Rxh�@JL��� 4@��T�h�!?��%Z�@�!T�M�ٿ+�*Rxh�@JL��� 4@��T�h�!?��%Z�@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@{��ٿ���
�O�@��>64@ 𲵐!?�B/r���@�!�8߂ٿ;�n�i�@j|U�;4@���А!?�i�6���@����ٿ�N�f��@�=�4@�Y�pϐ!?]��r��@����ٿ�N�f��@�=�4@�Y�pϐ!?]��r��@����ٿ�N�f��@�=�4@�Y�pϐ!?]��r��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�r !�ٿ��3�҉�@��;K�4@a{z��!?��.ɔ��@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�W�#�|ٿ�O�a��@�ʓ�4@��N`��!?4'9b�@�w��C�ٿ�p)
��@O��X4@[�a5��!?߈��3�@�w��C�ٿ�p)
��@O��X4@[�a5��!?߈��3�@�t�yC�ٿIk+�X-�@�Ў
4@!DN1��!?��:R��@�t�yC�ٿIk+�X-�@�Ў
4@!DN1��!?��:R��@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@vO�T�ٿ�Q[~���@���͞4@p9�"q�!??�<�@�@��M�	�ٿoT?�I��@�;"o� 4@����!?
i{C-I�@��M�	�ٿoT?�I��@�;"o� 4@����!?
i{C-I�@��M�	�ٿoT?�I��@�;"o� 4@����!?
i{C-I�@��M�	�ٿoT?�I��@�;"o� 4@����!?
i{C-I�@:l��~ٿ�8�����@�O���4@Z��#��!?h�hw���@:l��~ٿ�8�����@�O���4@Z��#��!?h�hw���@:l��~ٿ�8�����@�O���4@Z��#��!?h�hw���@Y���Áٿʁ?࣍�@��a 4@r���q�!?zԓ6�@Y���Áٿʁ?࣍�@��a 4@r���q�!?zԓ6�@Y���Áٿʁ?࣍�@��a 4@r���q�!?zԓ6�@Y���Áٿʁ?࣍�@��a 4@r���q�!?zԓ6�@ ��'�ٿy���J�@��U�4@��I���!?�^�m_�@ ��'�ٿy���J�@��U�4@��I���!?�^�m_�@ ��'�ٿy���J�@��U�4@��I���!?�^�m_�@<�-�ٿ�;o. ��@��}#? 4@I�$I��!?"���*�@�� �ҋٿ�BU��
�@:���� 4@�*�	x�!?2<�	/�@Q�(�F�ٿ��I�@�	��;4@:W����!?�k��~��@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@$=�ŋٿh��Mx��@�1�p4@��5�u�!?ø*f6�@���[�ٿ�H����@K=�?4@8�_�W�!?~��Lb�@���[�ٿ�H����@K=�?4@8�_�W�!?~��Lb�@���[�ٿ�H����@K=�?4@8�_�W�!?~��Lb�@�ԉ~�ٿ�vD�q��@��l>[4@ҡ�b�!?���}��@�ԉ~�ٿ�vD�q��@��l>[4@ҡ�b�!?���}��@�ԉ~�ٿ�vD�q��@��l>[4@ҡ�b�!?���}��@�ԉ~�ٿ�vD�q��@��l>[4@ҡ�b�!?���}��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@ђ�JI�ٿ#��gf�@����
4@y����!?r��ԣ��@�AO��ٿ���+�@P�b�4@#J0�!?�ei!�@U5�Z�ٿ�c=(�_�@-s�i	4@H�o0�!?�wF� 2�@U5�Z�ٿ�c=(�_�@-s�i	4@H�o0�!?�wF� 2�@U5�Z�ٿ�c=(�_�@-s�i	4@H�o0�!?�wF� 2�@�4����ٿ�I�,��@�O#84@8w��&�!?�]�t���@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@!T\��}ٿ��!���@��1�4@o�Ր!?�����@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@WP�ٿo��~�@f��7�4@�YE���!?����6V�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�3�g�ٿ��i�Z��@�6��x4@&��Ӑ!?����8�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�~M`�ٿ�n��@�`	�4@>�׭�!?��Ҙ�@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@�IXt�ٿԊ�p�@�J�4@G<����!?�Q�
T��@5�ǰy�ٿ������@�em��4@��b��!?K�:y�@5�ǰy�ٿ������@�em��4@��b��!?K�:y�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@Ǧ�ꆍٿ�Fg|�@=���4@4&3�j�!?k��0�@�D��ٿ"|�;�v�@� ,e4@ǫ�m!?��0w��@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��
P}ٿ����@s�1ku4@0���!?٦�`�u�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@��k߻�ٿ�ҧ�XQ�@��F4@*���ؐ!?�x~��O�@Rvfσٿ�8%����@�iy�4@����!?9vj�R��@
��ևٿ��)q��@��+��4@#O����!?�u �[��@
��ևٿ��)q��@��+��4@#O����!?�u �[��@� �d�ٿD�����@� V�4@��s��!?�&�R;�@� �d�ٿD�����@� V�4@��s��!?�&�R;�@� �d�ٿD�����@� V�4@��s��!?�&�R;�@� �d�ٿD�����@� V�4@��s��!?�&�R;�@� �d�ٿD�����@� V�4@��s��!?�&�R;�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@XH�8�ٿ��Fƍ��@9�'a��3@;���!?��&n�M�@������ٿ{%H�I�@��3��4@�1�Ǩ�!??��2�b�@IޟDx�ٿ���B,�@�ڪ��4@�8�Ɛ!?��%2E��@IޟDx�ٿ���B,�@�ڪ��4@�8�Ɛ!?��%2E��@Q���ٿ)���*��@�"��4@d��!?����u�@Q���ٿ)���*��@�"��4@d��!?����u�@Q���ٿ)���*��@�"��4@d��!?����u�@Q���ٿ)���*��@�"��4@d��!?����u�@Q���ٿ)���*��@�"��4@d��!?����u�@Q���ٿ)���*��@�"��4@d��!?����u�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@@��"��ٿ������@���� 4@ShM0ɐ!?Wֱ�@��nVуٿ>n�)�P�@DY9~4@�O?ː!?m_5}���@��nVуٿ>n�)�P�@DY9~4@�O?ː!?m_5}���@��nVуٿ>n�)�P�@DY9~4@�O?ː!?m_5}���@��nVуٿ>n�)�P�@DY9~4@�O?ː!?m_5}���@�?C�ٿ�ު7Y��@�&�\g 4@���ݐ!?[5�ǟ�@�?C�ٿ�ު7Y��@�&�\g 4@���ݐ!?[5�ǟ�@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@xM�L��ٿ���R��@!�[/Y4@����{�!?Щq���@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�a�;Ԓٿ��HV_��@�F㻝4@�Q��q�!?��d��@�D��\�ٿ]�d�~f�@u�N4@RI��!?A�r"��@�D��\�ٿ]�d�~f�@u�N4@RI��!?A�r"��@h8E�ƀٿ��a7�@��b
4@�0�!?.D��g��@h8E�ƀٿ��a7�@��b
4@�0�!?.D��g��@h8E�ƀٿ��a7�@��b
4@�0�!?.D��g��@��l�>�ٿ�=���@,y%���3@�����!?)K#� l�@��l�>�ٿ�=���@,y%���3@�����!?)K#� l�@��l�>�ٿ�=���@,y%���3@�����!?)K#� l�@��l�>�ٿ�=���@,y%���3@�����!?)K#� l�@��l�>�ٿ�=���@,y%���3@�����!?)K#� l�@����ٿ�]0�f��@l���}4@���qӐ!?��4���@0b)hz�ٿ�&����@m*��Y4@��2P��!?f�^/D��@0b)hz�ٿ�&����@m*��Y4@��2P��!?f�^/D��@0b)hz�ٿ�&����@m*��Y4@��2P��!?f�^/D��@����6�ٿ��p�1��@���4@��׼��!?e��v���@����6�ٿ��p�1��@���4@��׼��!?e��v���@����6�ٿ��p�1��@���4@��׼��!?e��v���@����6�ٿ��p�1��@���4@��׼��!?e��v���@����6�ٿ��p�1��@���4@��׼��!?e��v���@إ���ٿ�?N��@,(j�b4@C�}��!?v�P��@إ���ٿ�?N��@,(j�b4@C�}��!?v�P��@إ���ٿ�?N��@,(j�b4@C�}��!?v�P��@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@F�N��ٿ���p/��@�n��4@�x)֐!?G��Z�@��T�U�ٿ��t��@$<.�;4@:A9��!?v'q�:��@��T�U�ٿ��t��@$<.�;4@:A9��!?v'q�:��@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@��wPٿ�A��ٻ�@��4@�3���!?����3�@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@�]���ٿ��}kEr�@�ʷ�4@�,ے�!?�p�N���@q�����ٿ����T�@Τ΁�4@���_��!?*�y��@q�����ٿ����T�@Τ΁�4@���_��!?*�y��@q�����ٿ����T�@Τ΁�4@���_��!?*�y��@q�����ٿ����T�@Τ΁�4@���_��!?*�y��@���$�ٿ��N��b�@���[�4@��k!Ӑ!?\���"�@���$�ٿ��N��b�@���[�4@��k!Ӑ!?\���"�@c���1�ٿ�s2ߥt�@1kޚT4@:9ѐ!?(�\����@c���1�ٿ�s2ߥt�@1kޚT4@:9ѐ!?(�\����@c���1�ٿ�s2ߥt�@1kޚT4@:9ѐ!?(�\����@c���1�ٿ�s2ߥt�@1kޚT4@:9ѐ!?(�\����@c���1�ٿ�s2ߥt�@1kޚT4@:9ѐ!?(�\����@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@4�vl��ٿrM}���@��pd�4@��+2�!?�2��C�@���рٿ5�r���@���"4@�����!?��f���@q�x�k�ٿU���p��@�����4@�e8��!?BH��@q�x�k�ٿU���p��@�����4@�e8��!?BH��@q�x�k�ٿU���p��@�����4@�e8��!?BH��@q�x�k�ٿU���p��@�����4@�e8��!?BH��@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@@��o��ٿ9=�2��@pL�T4@2M�{А!?m��ɛ�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@a���M�ٿ�FM����@��d&^4@�ӷĐ!?XH���m�@Ӭ��׉ٿ�t��*�@�eUM�4@�vĺא!?�^��c�@����I�ٿ2�
�l�@<�$�Q4@�r��א!?^�(M��@����I�ٿ2�
�l�@<�$�Q4@�r��א!?^�(M��@��]Z�ٿ�[w���@�Pp4@5��� �!?Q�0���@��]Z�ٿ�[w���@�Pp4@5��� �!?Q�0���@O#�[߄ٿ5��J���@Y��x�4@j�/�!?�����@f.�Q	�ٿ",�Y��@�V��4@Ô�ؐ!?$�ƅ���@�˹T-�ٿ@gv���@�[�54@\��;��!?�( 7e�@w�z��ٿ�B{����@�xX�4@|�_Y�!?U��쏡�@w�z��ٿ�B{����@�xX�4@|�_Y�!?U��쏡�@w�z��ٿ�B{����@�xX�4@|�_Y�!?U��쏡�@w�z��ٿ�B{����@�xX�4@|�_Y�!?U��쏡�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@U'�S�ٿD�7�'b�@ju'��4@<�o؜�!?��M)�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@�CE�ٿyB�4�e�@��E>�4@4_�>��!?�]��Ɲ�@C�5H�ٿ��b%��@u���|4@B����!?�b��p�@C�5H�ٿ��b%��@u���|4@B����!?�b��p�@E-�#I�ٿ8�檷��@ź{"g4@x�輐!?2��&�@�S�{��ٿ�{��4�@��94@�!??����@�S�{��ٿ�{��4�@��94@�!??����@�S�{��ٿ�{��4�@��94@�!??����@�S�{��ٿ�{��4�@��94@�!??����@�S�{��ٿ�{��4�@��94@�!??����@Ո�Ćٿ�q[@�n�@�Ǔ�@4@/�2@ǐ!?73�s��@Ո�Ćٿ�q[@�n�@�Ǔ�@4@/�2@ǐ!?73�s��@�z�T
�ٿ���G
��@Qmm5�4@X*��Ր!?��_\�a�@�z�T
�ٿ���G
��@Qmm5�4@X*��Ր!?��_\�a�@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�5	`�ٿ_�=�@�Duy�4@7��y�!?ѩG���@�ʒ�ٿ��v�@J��34@�e\��!?A���ݜ�@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@�OW1�ٿ�1aIY�@�[5��4@�D*)ݐ!?��]��@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@AF�w�ٿg�G��@��{3�4@}؆uː!?E A�\E�@��y�ٿ�����@>mi L4@���-�!?E@ݸr.�@��y�ٿ�����@>mi L4@���-�!?E@ݸr.�@�ְ�ދٿ9�:4�!�@Y�ZlG4@���
�!?4��|.�@�ְ�ދٿ9�:4�!�@Y�ZlG4@���
�!?4��|.�@n,Ǚהٿ�� ��@7�fE�4@��Ր!?����S��@��>T�ٿ"��ɂ^�@iv�^�4@��HpӐ!?��8�4�@��>T�ٿ"��ɂ^�@iv�^�4@��HpӐ!?��8�4�@��>T�ٿ"��ɂ^�@iv�^�4@��HpӐ!?��8�4�@i~_vx�ٿ�%� ���@%���Y4@�\�^��!?�>����@i~_vx�ٿ�%� ���@%���Y4@�\�^��!?�>����@i~_vx�ٿ�%� ���@%���Y4@�\�^��!?�>����@i~_vx�ٿ�%� ���@%���Y4@�\�^��!?�>����@i~_vx�ٿ�%� ���@%���Y4@�\�^��!?�>����@x�#�ٿ^�/����@˅_�4@8����!?��9on�@��'�ـٿ�!��/��@Ud�o4@9d"���!?���f�'�@��'�ـٿ�!��/��@Ud�o4@9d"���!?���f�'�@��'�ـٿ�!��/��@Ud�o4@9d"���!?���f�'�@��'�ـٿ�!��/��@Ud�o4@9d"���!?���f�'�@S�e��ٿ�J���@���4@i�d��!?��_���@S�e��ٿ�J���@���4@i�d��!?��_���@S�e��ٿ�J���@���4@i�d��!?��_���@S�e��ٿ�J���@���4@i�d��!?��_���@=l�\��ٿj�X�]�@m��x�4@�����!?�v�́��@=l�\��ٿj�X�]�@m��x�4@�����!?�v�́��@=l�\��ٿj�X�]�@m��x�4@�����!?�v�́��@]�Z�+~ٿ����:��@���U.4@�x�J��!?�2F��@]�Z�+~ٿ����:��@���U.4@�x�J��!?�2F��@]�Z�+~ٿ����:��@���U.4@�x�J��!?�2F��@�$)�5�ٿ�a)� �@m9�)4@��B���!?�c�l�z�@�l�ٝ�ٿ(�P@A�@؎:��4@���zِ!?����Ö�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@�^�c�ٿN82X���@���4@Ш�Ɛ!?o�
ݲ�@��Z�ٿ!O���d�@*u�4@�_2��!?�|����@��Z�ٿ!O���d�@*u�4@�_2��!?�|����@MQ��_�ٿd�Y|T��@cb�)4@�T9�[�!?aLW"�@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@��Nߋٿ̫��>	�@���f�4@_��y�!?VӤ3 �@`ss��ٿ��_�!0�@�Ͱ�
4@l��<��!?����E�@`ss��ٿ��_�!0�@�Ͱ�
4@l��<��!?����E�@��/�D�ٿ �_���@�)���4@�"O/��!?�V]t��@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@E�#�ٿV�S���@*Ʃ��4@5"�Gِ!?�2R�-�@t��h�|ٿ�`VQ)�@���4@����!?a�ƕ�C�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@$�l�ٿ/���\�@⸄�� 4@�e��Ő!?e�p�#�@���v��ٿ�l�(u��@��8Am4@Mf+MŐ!?.P����@\Uy�O�ٿůY���@ox| 4@�:���!?��\���@jm��}ٿ	e����@d���_�3@3@�U��!?oR�~��@jm��}ٿ	e����@d���_�3@3@�U��!?oR�~��@bX1�o�ٿ�r�k��@�G�M��3@��`ç�!?t;��Z��@oH-�ٿ�2-Wk�@�`���3@q�oq�!? ��swY�@��N_�ٿ�tt�p�@1��4@�ѵ_Ԑ!?��N���@��N_�ٿ�tt�p�@1��4@�ѵ_Ԑ!?��N���@���Th�ٿ�`Ӗ�c�@�n�U4@: T{��!?#�!#`��@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@s�ڂ�ٿ��I=��@D�>'*4@��Ւ�!?u����@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@�ވ���ٿW�e����@`�}&4@� 묲�!?�~�g(�@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@`�KC�ٿ�6�I��@[��"�4@�ܯ_��!?�M���@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@z"�_��ٿ���i���@���tR4@�X�!?�O�)r�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@t�fJ�ٿz�+}�@Z��I4@G���!?�n��qJ�@C&��
�ٿ��g[��@�aA��4@��5ñ�!?�8�����@*��,��ٿg�Z
��@�����4@c���r�!?n�Ω���@c����ٿ��m6@��@�]i�j4@7��`�!?��ϗ��@�kM'�ٿZoy]��@��(9G4@b�v68�!?#�2���@�kM'�ٿZoy]��@��(9G4@b�v68�!?#�2���@I���H�ٿr/a���@�6S��4@Z��S2�!?8��GM�@I���H�ٿr/a���@�6S��4@Z��S2�!?8��GM�@I���H�ٿr/a���@�6S��4@Z��S2�!?8��GM�@I���H�ٿr/a���@�6S��4@Z��S2�!?8��GM�@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@��񌻃ٿ���q���@�5֠�4@��r{�!?	�#'C��@�����ٿK���{�@*�Va4@L5:���!?���r_��@�����ٿK���{�@*�Va4@L5:���!?���r_��@�]N���ٿs8r lv�@���c4@&���!?�~����@n�w{�ٿ�N �-�@k�)y�4@�S�&��!? �����@n�w{�ٿ�N �-�@k�)y�4@�S�&��!? �����@n�w{�ٿ�N �-�@k�)y�4@�S�&��!? �����@n�w{�ٿ�N �-�@k�)y�4@�S�&��!? �����@n�w{�ٿ�N �-�@k�)y�4@�S�&��!? �����@}�b�ٿ.t&q�@a�
�4@���.m�!?�� �[�@}�b�ٿ.t&q�@a�
�4@���.m�!?�� �[�@!dWևٿwQ�P%��@f�W4@�'n��!?��=:���@!dWևٿwQ�P%��@f�W4@�'n��!?��=:���@!dWևٿwQ�P%��@f�W4@�'n��!?��=:���@!dWևٿwQ�P%��@f�W4@�'n��!?��=:���@!dWևٿwQ�P%��@f�W4@�'n��!?��=:���@j�~�ٿno��E�@��Oex4@�!ΐ!?V�?�Z�@j�~�ٿno��E�@��Oex4@�!ΐ!?V�?�Z�@��x1܍ٿ��3�={�@��	4@D�d���!?�8R�G�@��W�R�ٿ� �K���@�{ǆ	4@JÍ��!?� ��	��@��W�R�ٿ� �K���@�{ǆ	4@JÍ��!?� ��	��@3�
Gw�ٿ�����o�@:x�T�4@�z���!?�DLi�@3�
Gw�ٿ�����o�@:x�T�4@�z���!?�DLi�@3�
Gw�ٿ�����o�@:x�T�4@�z���!?�DLi�@3�
Gw�ٿ�����o�@:x�T�4@�z���!?�DLi�@�)s<r�ٿp�����@�S1�4@Aeϭɐ!?J
�ބD�@+f�ɏٿ��,�A�@���H4@T�j9��!?�sw����@+f�ɏٿ��,�A�@���H4@T�j9��!?�sw����@+f�ɏٿ��,�A�@���H4@T�j9��!?�sw����@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@1B�+V�ٿx5��=�@��g�4@�1�a��!?�vZH7.�@��*	��ٿ��CI���@����u4@b�P헐!?ߐ&ut$�@��*	��ٿ��CI���@����u4@b�P헐!?ߐ&ut$�@�am~�ٿ�ڑř��@�Wc�4@	�4��!?~�M���@�am~�ٿ�ڑř��@�Wc�4@	�4��!?~�M���@�am~�ٿ�ڑř��@�Wc�4@	�4��!?~�M���@�am~�ٿ�ڑř��@�Wc�4@	�4��!?~�M���@�am~�ٿ�ڑř��@�Wc�4@	�4��!?~�M���@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@pi1�}ٿ�8����@%{��4@׎�lǐ!?�J�4�@ U�>ЄٿIa����@du�J4@whAÐ!?`�)b�@ U�>ЄٿIa����@du�J4@whAÐ!?`�)b�@ U�>ЄٿIa����@du�J4@whAÐ!?`�)b�@arD��ٿ���}�E�@�84@���ِ!?0�u���@arD��ٿ���}�E�@�84@���ِ!?0�u���@���
|ٿ����+��@�ߣ�4@|l|ѐ!?�������@���
|ٿ����+��@�ߣ�4@|l|ѐ!?�������@���
|ٿ����+��@�ߣ�4@|l|ѐ!?�������@���
|ٿ����+��@�ߣ�4@|l|ѐ!?�������@t��U.�ٿ"*U�s�@��\$ 4@���̐!?��2`�@�6R��ٿ<��с�@�L4@�ϋʳ�!?���'��@�6R��ٿ<��с�@�L4@�ϋʳ�!?���'��@�6R��ٿ<��с�@�L4@�ϋʳ�!?���'��@�6R��ٿ<��с�@�L4@�ϋʳ�!?���'��@�6R��ٿ<��с�@�L4@�ϋʳ�!?���'��@g�����ٿ�)D�H�@-��54@*�	�!?�[�sY�@b�Zφٿ)�ˑ��@V��	4@��Mtѐ!?��B�6��@��c�C�ٿ��Fxj!�@�k��4@ޯ,�א!?���<,j�@��c�C�ٿ��Fxj!�@�k��4@ޯ,�א!?���<,j�@��c�C�ٿ��Fxj!�@�k��4@ޯ,�א!?���<,j�@��u�~ٿ|������@t��`R	4@�(�!?��8���@��u�~ٿ|������@t��`R	4@�(�!?��8���@��u�~ٿ|������@t��`R	4@�(�!?��8���@\yO3��ٿ&���V�@���4@�Fσ�!?{��t�:�@\yO3��ٿ&���V�@���4@�Fσ�!?{��t�:�@�H`��ٿ월��C�@�!��4@�l0��!?����W�@�H`��ٿ월��C�@�!��4@�l0��!?����W�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@���^A�ٿ����5�@���4@8�q���!?�<u¨>�@E�K,a�ٿ&Z�&d�@���r4@B�Ɩ��!?�!24��@E�K,a�ٿ&Z�&d�@���r4@B�Ɩ��!?�!24��@A�z;��ٿ�ެب��@+�K4@2Y=ː!?��Й��@A�z;��ٿ�ެب��@+�K4@2Y=ː!?��Й��@A�z;��ٿ�ެب��@+�K4@2Y=ː!?��Й��@A�z;��ٿ�ެب��@+�K4@2Y=ː!?��Й��@A�z;��ٿ�ެب��@+�K4@2Y=ː!?��Й��@�"h�ٿz�z<J�@����4@Rt�Ӑ!?Iα[ �@�"h�ٿz�z<J�@����4@Rt�Ӑ!?Iα[ �@V�Ӿ^�ٿ5#_ h��@A��O�4@�DTԐ!?��̮&�@V�Ӿ^�ٿ5#_ h��@A��O�4@�DTԐ!?��̮&�@V�Ӿ^�ٿ5#_ h��@A��O�4@�DTԐ!?��̮&�@V�Ӿ^�ٿ5#_ h��@A��O�4@�DTԐ!?��̮&�@V�Ӿ^�ٿ5#_ h��@A��O�4@�DTԐ!?��̮&�@����~ٿ�o���2�@p�Cq%4@��|׻�!?\�:I�@��[A�ٿ&Ϳ����@�"sD�4@o���y�!?O���@��[A�ٿ&Ϳ����@�"sD�4@o���y�!?O���@��[A�ٿ&Ϳ����@�"sD�4@o���y�!?O���@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@#�_�ٿ�Y,1���@��/%�4@I;JL�!?3$N\�@~F�n��ٿ�g����@ˬ"�d4@�H�&a�!?�i���@	��ٿsX����@5?��8 4@+e�!?���E��@	��ٿsX����@5?��8 4@+e�!?���E��@	��ٿsX����@5?��8 4@+e�!?���E��@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@���<��ٿ��J3*��@��\�� 4@ئ?Y��!?�#�b���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@|��_�ٿ;�3�Z��@1��4@Q�F�!?�<���@lԁ1�ٿ�t7 �7�@��Gr�4@`�
��!?�ʭa���@lԁ1�ٿ�t7 �7�@��Gr�4@`�
��!?�ʭa���@lԁ1�ٿ�t7 �7�@��Gr�4@`�
��!?�ʭa���@lԁ1�ٿ�t7 �7�@��Gr�4@`�
��!?�ʭa���@m��B��ٿR���¯�@��J�j�3@/�"̐!?�[���N�@���&��ٿ=�����@���7B 4@��bF��!?�-&�[�@���&��ٿ=�����@���7B 4@��bF��!?�-&�[�@���&��ٿ=�����@���7B 4@��bF��!?�-&�[�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@�	<���ٿy� ޿�@$ۿ��4@b���ؐ!?�ĺ�&^�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@9
t?�}ٿ���h�q�@%c׬�4@
�-�!?�J-}�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@1S���ٿ�TP�K��@�;9�4@H ��!?�I�#O4�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@�G�w��ٿ	���dr�@T�@4@�jWv�!?�6WG|;�@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@y���ٿ�Q���@��V�� 4@%]Ӻ�!?S8zK��@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@��a��ٿ:���*�@Fe�4@"����!?6��!�(�@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@���<�ٿ��t��?�@����A4@�#��z�!?�,�,��@}��-ٿ&[����@���4@���&��!?�R�mU��@}��-ٿ&[����@���4@���&��!?�R�mU��@}��-ٿ&[����@���4@���&��!?�R�mU��@}��-ٿ&[����@���4@���&��!?�R�mU��@}��-ٿ&[����@���4@���&��!?�R�mU��@}��-ٿ&[����@���4@���&��!?�R�mU��@_=�U��ٿ�ո�3�@�5�4@d>S�!?NW�9��@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@H�H�Љٿ��T���@�)c4@�%CM�!?���2�@�!��_�ٿ��G�-��@�X�)4@g[���!?�R�4�@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@z��F�ٿ@�p��@�/��4@@�h�!?��+��@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@N��ˈٿsNM2��@����4@e��c��!?Z�����@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��ٿ)�!�β�@����4@��H�K�!?FZ+�2�@��3ڂ�ٿ���ԠR�@�N�OQ4@b��t�!?�*����@��3ڂ�ٿ���ԠR�@�N�OQ4@b��t�!?�*����@��3ڂ�ٿ���ԠR�@�N�OQ4@b��t�!?�*����@��3ڂ�ٿ���ԠR�@�N�OQ4@b��t�!?�*����@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@c����ٿ�O�YZ.�@��%�4@8#hs�!?���?U��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@�k�(�|ٿ�����Z�@&��4@�m�
�!?;�_�,��@Sh A|ٿ�A ����@o��c�4@�����!?ͬ�4�;�@Sh A|ٿ�A ����@o��c�4@�����!?ͬ�4�;�@Sh A|ٿ�A ����@o��c�4@�����!?ͬ�4�;�@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@���q^�ٿ�������@U	|4@ '����!?VH�<=��@8�)��ٿ������@�!��84@���
��!?�ƈ���@�"��M�ٿd�2���@�ҥ�D4@��Qg��!?s
'8��@�"��M�ٿd�2���@�ҥ�D4@��Qg��!?s
'8��@��T���ٿd6*b�@����f4@K���o�!?z�ҁ�@j�j%r�ٿ�=A�$2�@��߭4@���ߐ!?Jhj��@j�j%r�ٿ�=A�$2�@��߭4@���ߐ!?Jhj��@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@Ͳ�qX�ٿ#����@	J��4@�8餇�!?�u��|7�@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@�h勎ٿ�hM�.�@�(cG�4@�u�!?�^����@POŁo�ٿ_�G���@�'OG�4@)?f�Ր!?viH�_��@POŁo�ٿ_�G���@�'OG�4@)?f�Ր!?viH�_��@POŁo�ٿ_�G���@�'OG�4@)?f�Ր!?viH�_��@�9h@�}ٿ,W�^��@3�X4@A8{�!?��[���@�VU\�ٿ0^�f��@#�g�84@��&g�!?}U��u�@�VU\�ٿ0^�f��@#�g�84@��&g�!?}U��u�@PCi�B�ٿ��&����@��n�}4@�e�1u�!?�ٕzV�@PCi�B�ٿ��&����@��n�}4@�e�1u�!?�ٕzV�@h���ٿ��/��@�!1��4@�h�NS�!?�R좒b�@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@xVה�ٿ�.5�D��@�^с4@��5zn�!?�n+mF��@a�b5�ٿd������@�.2o 4@Й����!?<�|���@a�b5�ٿd������@�.2o 4@Й����!?<�|���@a�b5�ٿd������@�.2o 4@Й����!?<�|���@a�b5�ٿd������@�.2o 4@Й����!?<�|���@a�b5�ٿd������@�.2o 4@Й����!?<�|���@a�b5�ٿd������@�.2o 4@Й����!?<�|���@5Sp��~ٿYw�]m��@�P.A��3@�>���!?> {�%�@5Sp��~ٿYw�]m��@�P.A��3@�>���!?> {�%�@c��~ٿ��&���@���&4@���Z��!?��1����@c��~ٿ��&���@���&4@���Z��!?��1����@c��~ٿ��&���@���&4@���Z��!?��1����@FD��ٿ��e����@���+4@�:ʐ!?f��h��@FD��ٿ��e����@���+4@�:ʐ!?f��h��@FD��ٿ��e����@���+4@�:ʐ!?f��h��@FD��ٿ��e����@���+4@�:ʐ!?f��h��@��_�ٿ0���}�@�WA�4@� ,�ɐ!?�bq��p�@��_�ٿ0���}�@�WA�4@� ,�ɐ!?�bq��p�@���0؀ٿgS����@"W��4@?�*`Ր!?|8̨ۨ�@���0؀ٿgS����@"W��4@?�*`Ր!?|8̨ۨ�@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���ר�ٿ>�� ���@,�,�4@�luQ�!?��ծ��@���J�ٿ,y����@����4@+{"���!?m�a����@���J�ٿ,y����@����4@+{"���!?m�a����@���J�ٿ,y����@����4@+{"���!?m�a����@���J�ٿ,y����@����4@+{"���!?m�a����@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@[��x��ٿ�\!�@���k4@Ǖ~(|�!?��җѩ�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@z@(�l�ٿ\�c�s��@��� 4@G��E��!?�z]k�2�@ P�Z�ٿ���]��@���u�4@;�UW�!?�=�\�@ P�Z�ٿ���]��@���u�4@;�UW�!?�=�\�@ P�Z�ٿ���]��@���u�4@;�UW�!?�=�\�@ P�Z�ٿ���]��@���u�4@;�UW�!?�=�\�@ P�Z�ٿ���]��@���u�4@;�UW�!?�=�\�@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@#-=!�ٿ&��2�R�@�ӧ$�4@A@�"��!?�����@���ٿ{�"��K�@�C[4@	Q�k �!?3P���@µ�kH�ٿ5T�â�@p^W� 4@-�ډ�!?�XƄ�i�@µ�kH�ٿ5T�â�@p^W� 4@-�ډ�!?�XƄ�i�@µ�kH�ٿ5T�â�@p^W� 4@-�ډ�!?�XƄ�i�@zk���ٿ`�%�M��@B���4@��~!��!?�,�{�[�@zk���ٿ`�%�M��@B���4@��~!��!?�,�{�[�@zk���ٿ`�%�M��@B���4@��~!��!?�,�{�[�@zk���ٿ`�%�M��@B���4@��~!��!?�,�{�[�@zk���ٿ`�%�M��@B���4@��~!��!?�,�{�[�@P�X���ٿ���@\����4@x�ek+�!?f�&����@P�X���ٿ���@\����4@x�ek+�!?f�&����@P�X���ٿ���@\����4@x�ek+�!?f�&����@5)[�x�ٿ�c����@x���4@%�!�!?#_`����@5)[�x�ٿ�c����@x���4@%�!�!?#_`����@5)[�x�ٿ�c����@x���4@%�!�!?#_`����@5)[�x�ٿ�c����@x���4@%�!�!?#_`����@�RD��ٿX�	��@����4@%F�C�!?�&����@uk��هٿBb�26	�@���$4@Dې$�!?)�`o��@s���{�ٿ�Bܾt��@~���4@
�n��!?���bɟ�@�ʆ�~ٿ���+�@O�3y�4@��}�!?��$����@�ʆ�~ٿ���+�@O�3y�4@��}�!?��$����@�ʆ�~ٿ���+�@O�3y�4@��}�!?��$����@�ʆ�~ٿ���+�@O�3y�4@��}�!?��$����@Y�"x^{ٿ��"�}�@R�b�4@�L	p�!?f��f�@�Rd�yxٿ� �����@��2�_4@�(I���!?��6V���@�Rd�yxٿ� �����@��2�_4@�(I���!?��6V���@�Rd�yxٿ� �����@��2�_4@�(I���!?��6V���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@C�V��ٿ���8n�@�O�4@�1�g[�!?+�K���@4�Y�ٿm|b�ѣ�@�����4@���v��!?�Ey+���@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@�'�7U�ٿ]����@�u4LG 4@�I�g�!?.��G!�@͒�vX�ٿ�@G�@J�b���3@�ݮMɐ!?nj�2~��@���T�ٿ�8q>���@���Q54@4����!?�������@���T�ٿ�8q>���@���Q54@4����!?�������@���T�ٿ�8q>���@���Q54@4����!?�������@���T�ٿ�8q>���@���Q54@4����!?�������@���T�ٿ�8q>���@���Q54@4����!?�������@���T�ٿ�8q>���@���Q54@4����!?�������@g`b,�ٿ��, �@{��J� 4@gt���!?hV6B���@J�Y�w�ٿG�=2RV�@��iԾ4@�#�)�!?��Aޑa�@��(�Ȁٿv�xp�@?Z��� 4@�Wu(�!?��Π���@��(�Ȁٿv�xp�@?Z��� 4@�Wu(�!?��Π���@��(�Ȁٿv�xp�@?Z��� 4@�Wu(�!?��Π���@��(�Ȁٿv�xp�@?Z��� 4@�Wu(�!?��Π���@��Q��ٿ�;ǔŁ�@��G��4@`��$�!?LO�.��@��Q��ٿ�;ǔŁ�@��G��4@`��$�!?LO�.��@��Q��ٿ�;ǔŁ�@��G��4@`��$�!?LO�.��@��Q��ٿ�;ǔŁ�@��G��4@`��$�!?LO�.��@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@vyR��}ٿ-�����@��7?4@3�O2�!?xY�p�]�@AB����ٿ�|���@X��l4@�s��.�!?��J����@5L�)�ٿ'w�!g�@L,���4@�n��!?���F�~�@5L�)�ٿ'w�!g�@L,���4@�n��!?���F�~�@���(L�ٿev3=z~�@|��84@w��Cj�!?��r��M�@���(L�ٿev3=z~�@|��84@w��Cj�!?��r��M�@¼��ύٿ�M�`t��@�����4@��*��!?#�d����@¼��ύٿ�M�`t��@�����4@��*��!?#�d����@�@�t�ٿ��4=��@����4@�O�ǹ�!?o�cl��@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@]Q愂ٿ&�950/�@�N
C4@�^"���!?��seߙ�@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@����քٿ�D�/�@��	�Q4@�<$,��!?_FM��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@1���Q�ٿ�h�^��@`	��4@c��g��!?�-)��@hrZ�ٿ��GG¸�@&6o�4@���U~�!?�3-w�J�@hrZ�ٿ��GG¸�@&6o�4@���U~�!?�3-w�J�@�M�k�ٿ�:eB��@�3/:��3@�W�~�!?ы%����@4e�ڎ�ٿ��9h��@B�]�4@�b�\_�!?,*1����@4e�ڎ�ٿ��9h��@B�]�4@�b�\_�!?,*1����@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@��,5��ٿ2C���@��*t<4@�)4-��!?.���6��@9�+���ٿ��l&�@-Ov�4@����!?@ ��@$�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@T�=s�ٿmg�%���@�K��4@�+ِ!? ��Z�@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@1���-�ٿr}^���@��R��4@���l�!?�	��t��@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�lg\��ٿ���p�@?��j�4@�A�F�!?���	�@�DT��ٿN��X�p�@�yb��4@��ZK�!?CV_Y;�@�DT��ٿN��X�p�@�yb��4@��ZK�!?CV_Y;�@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@�:�\Z�ٿ��ñ���@K��\	4@��{'�!?�m+`M��@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@S�]��ٿv�Ѳ�@�Y�D*	4@#K׌ �!?)"u���@z����ٿ��u����@s���4@�{ː!?kџ�t2�@z����ٿ��u����@s���4@�{ː!?kџ�t2�@z����ٿ��u����@s���4@�{ː!?kџ�t2�@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@{"��ٿc�Y���@$aXi4@V�% b�!?��a���@Ȁ���ٿ?��d��@�ͣf� 4@��w"o�!?�����E�@Ȁ���ٿ?��d��@�ͣf� 4@��w"o�!?�����E�@Ȁ���ٿ?��d��@�ͣf� 4@��w"o�!?�����E�@Ȁ���ٿ?��d��@�ͣf� 4@��w"o�!?�����E�@Ȁ���ٿ?��d��@�ͣf� 4@��w"o�!?�����E�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@��9e�ٿ/��3.��@�ժ��4@X��?ܐ!?;���5�@x~�#H�ٿ�s����@�}V�4@t%��ސ!?��H��@x~�#H�ٿ�s����@�}V�4@t%��ސ!?��H��@x~�#H�ٿ�s����@�}V�4@t%��ސ!?��H��@x~�#H�ٿ�s����@�}V�4@t%��ސ!?��H��@x~�#H�ٿ�s����@�}V�4@t%��ސ!?��H��@<$0}ąٿ���2�@e�ﻅ 4@�X��ѐ!?�VS{9�@<$0}ąٿ���2�@e�ﻅ 4@�X��ѐ!?�VS{9�@<$0}ąٿ���2�@e�ﻅ 4@�X��ѐ!?�VS{9�@<$0}ąٿ���2�@e�ﻅ 4@�X��ѐ!?�VS{9�@n4̒��ٿU�]��@�^# 4@�%�RА!?I�?��J�@�<��ٿ@fm���@#͙F4@v�>$��!?F�U�)�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@c桉�ٿd��2�)�@q��7?4@Z%���!?���t�_�@v�+�ٿ�}�J��@��s�H4@�s����!?���c�@v�+�ٿ�}�J��@��s�H4@�s����!?���c�@v�+�ٿ�}�J��@��s�H4@�s����!?���c�@Hl���ٿe�nH��@�F���4@*�ђJ�!?���=^�@Hl���ٿe�nH��@�F���4@*�ђJ�!?���=^�@��晴ٿ�,S3W��@l�Y�4@2�脐!?�?�_�@��晴ٿ�,S3W��@l�Y�4@2�脐!?�?�_�@��晴ٿ�,S3W��@l�Y�4@2�脐!?�?�_�@-͓���ٿ�P���@�C
c4@���T�!?޶D|+�@-͓���ٿ�P���@�C
c4@���T�!?޶D|+�@-͓���ٿ�P���@�C
c4@���T�!?޶D|+�@0/�ٿm��x�@�zق}4@"�p�Q�!?�P!��@0/�ٿm��x�@�zق}4@"�p�Q�!?�P!��@0/�ٿm��x�@�zق}4@"�p�Q�!?�P!��@0/�ٿm��x�@�zق}4@"�p�Q�!?�P!��@�M�Q�ٿ.3�O�@N�j5�4@ֈ`��!?L�{l��@�M�Q�ٿ.3�O�@N�j5�4@ֈ`��!?L�{l��@�M�Q�ٿ.3�O�@N�j5�4@ֈ`��!?L�{l��@�M�Q�ٿ.3�O�@N�j5�4@ֈ`��!?L�{l��@M�$�6�ٿ�W� ���@e�J4@���2��!?,�>pB��@M�$�6�ٿ�W� ���@e�J4@���2��!?,�>pB��@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@Z#� �ٿ:����@FE3	4@l';�א!?|c�gW�@�Q���ٿ�N eP��@\[Z��4@
�����!?fq9gǖ�@wd�YL�ٿ���K�@�Ř�34@��u�ې!?P$c����@wd�YL�ٿ���K�@�Ř�34@��u�ې!?P$c����@=˛L��ٿ�;����@s>K+4@$7�6��!?q�ma��@=˛L��ٿ�;����@s>K+4@$7�6��!?q�ma��@=˛L��ٿ�;����@s>K+4@$7�6��!?q�ma��@=˛L��ٿ�;����@s>K+4@$7�6��!?q�ma��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@xxd��ٿK��܆��@��+��4@�À��!?�(/8��@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@� �,�~ٿ)o����@a5��4@,O_�ѐ!?¤�vJh�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@!`���ٿ��B'���@D&i��4@SAѐ!?dV�ז�@4W0�3�ٿ�@g!��@V�v�f4@�(y:��!?/�3'��@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@#�urQ�ٿ�'q���@Y|u� 4@�sf�!?�e�z�+�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@�4�@�ٿr���@Qe�|�4@v��!?P�mn�}�@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@DTS9�ٿEt�C5��@:��>�4@bi0P8�!?��F��@�����|ٿt�Bfu�@�*-R4@~4Ę�!?~�I�q�@�����|ٿt�Bfu�@�*-R4@~4Ę�!?~�I�q�@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@^�䧃ٿ�xP�͋�@d踹(4@���$��!?{�&��@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@��j��ٿx���-��@{���3@��N �!?У֊i:�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@�7t^�ٿ|�3�@ek�4@Z���!?�Q��-"�@[=Z�ٿ��%�3)�@qI<�4@ KŲ�!?V7�b�U�@[=Z�ٿ��%�3)�@qI<�4@ KŲ�!?V7�b�U�@[=Z�ٿ��%�3)�@qI<�4@ KŲ�!?V7�b�U�@[=Z�ٿ��%�3)�@qI<�4@ KŲ�!?V7�b�U�@���K�ٿ��u���@��?�4@�}nՐ!?�=����@���K�ٿ��u���@��?�4@�}nՐ!?�=����@���K�ٿ��u���@��?�4@�}nՐ!?�=����@���K�ٿ��u���@��?�4@�}nՐ!?�=����@���K�ٿ��u���@��?�4@�}nՐ!?�=����@(5{d�ٿ!6"5��@:��a�4@�����!?����D�@(5{d�ٿ!6"5��@:��a�4@�����!?����D�@(5{d�ٿ!6"5��@:��a�4@�����!?����D�@(5{d�ٿ!6"5��@:��a�4@�����!?����D�@(5{d�ٿ!6"5��@:��a�4@�����!?����D�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@��<I~ٿ���,�7�@v]�i	4@��Ԑ!?v���%�@�����~ٿ�_6���@]E��,	4@86<u�!?r��Z��@̼�ٿž4ӈM�@���8�4@��?�q�!?�TŦ��@N�.(�ٿ$Y���/�@P���4@8�@͐!?��j�7��@����'�ٿ��Ӆ��@�ȼJ�4@^t�~�!?��o@���@��CuL�ٿmq��>��@Ω>g�4@�؇XI�!?<'�Y��@�� čٿ���1���@MvF�M4@�?`�Ӑ!?q.)����@�� čٿ���1���@MvF�M4@�?`�Ӑ!?q.)����@_���:�ٿI"'	�@�F���4@λOi��!?�ƺ����@_���:�ٿI"'	�@�F���4@λOi��!?�ƺ����@_���:�ٿI"'	�@�F���4@λOi��!?�ƺ����@_���:�ٿI"'	�@�F���4@λOi��!?�ƺ����@��%���ٿ@�Ԑt��@z��� 4@�Ax�!?�r��SH�@��%���ٿ@�Ԑt��@z��� 4@�Ax�!?�r��SH�@T��}m�ٿ�X���	�@���4@�Ԍ�ؐ!?����Z��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@�e%s�ٿOs��N�@B��4@��g�Ր!?׎w�%��@2Yke�ٿ43lu��@��=�4@Ly�1�!?�:2M�@2Yke�ٿ43lu��@��=�4@Ly�1�!?�:2M�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@�9-�ٿ��&ݬx�@Z�\�_4@G)�!?�.���F�@5�b$�ٿ��B_��@�Ɇ���3@n�����!?��!<	�@5�b$�ٿ��B_��@�Ɇ���3@n�����!?��!<	�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@S�M��ٿ��-���@�GQ"K4@��<MC�!?���'�@�Lu��ٿ�-zSH�@��)�4@��;�!?������@�Lu��ٿ�-zSH�@��)�4@��;�!?������@�Lu��ٿ�-zSH�@��)�4@��;�!?������@�Lu��ٿ�-zSH�@��)�4@��;�!?������@�Lu��ٿ�-zSH�@��)�4@��;�!?������@#��2�ٿ��t��@�/��	4@�j�U!?�$�m���@#��2�ٿ��t��@�/��	4@�j�U!?�$�m���@#��2�ٿ��t��@�/��	4@�j�U!?�$�m���@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@B�S`�ٿ,z�7�:�@;� @\4@Z �x�!?�+D����@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@T����ٿ1�-y1��@�5�:4@M��Wא!?��7�.�@+i�ٿ<��%�L�@��CB4@��5�P�!?�pT�~2�@�P���ٿ�K��q��@˜�Eo4@'`�运!?�u��r�@�P���ٿ�K��q��@˜�Eo4@'`�运!?�u��r�@�P���ٿ�K��q��@˜�Eo4@'`�运!?�u��r�@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@'�H)�ٿ����V�@�8-�4@��sY��!?�1}����@&���F�ٿ��8wH�@�/;u$4@�m��!?�d����@&���F�ٿ��8wH�@�/;u$4@�m��!?�d����@�PR��ٿ�B��c�@����4@8�k��!?~0�hY�@�PR��ٿ�B��c�@����4@8�k��!?~0�hY�@��Q��ٿ��ʫs��@�N24@~�t"�!?�u9g��@��Q��ٿ��ʫs��@�N24@~�t"�!?�u9g��@��Q��ٿ��ʫs��@�N24@~�t"�!?�u9g��@z�R�N�ٿ�Tc�kI�@��A�4@TM�ِ!?� ���@z�R�N�ٿ�Tc�kI�@��A�4@TM�ِ!?� ���@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@�A�R�ٿ��3ӹ��@�Jv6/4@2;`�!?*�C�t�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@���)�ٿ �.p��@h)y��4@��C�P�!?�0���	�@O�0	�ٿ����N�@�$�U	4@���>e�!?r?E	w��@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@�Y$�ٿa�xr�@Ԉ!D�4@t�&�ڐ!?��F�	�@���yk�ٿ�6 ��@C��4@�s�Y��!?Jcy�
�@��%�ٿ(����@9Q'��4@�KŐ!?IV*\�@��%�ٿ(����@9Q'��4@�KŐ!?IV*\�@��%�ٿ(����@9Q'��4@�KŐ!?IV*\�@dx_Yٿ*
��\�@�?�<4@�ut�ې!?�W
�W��@dx_Yٿ*
��\�@�?�<4@�ut�ې!?�W
�W��@�M���ٿ�(w`�=�@��
�4@V����!?��h���@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@���ٿ\�i��g�@ݕ%b4@eR���!?	�����@J�U�ٿ�c���@�g4@@Z���!?"�6��@J�U�ٿ�c���@�g4@@Z���!?"�6��@�&��ٿ� Ԣ�5�@?�;�4@�Ǆ�ʐ!?��
���@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@��& V�ٿ���/���@`";t�4@�@Es��!?j?����@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@����ٿ��թ�@P�YAg4@�Q�	�!?�[��Mc�@���{�ٿ��u3Oe�@ʙ�߮4@տ�Ǻ�!?������@���{�ٿ��u3Oe�@ʙ�߮4@տ�Ǻ�!?������@���{�ٿ��u3Oe�@ʙ�߮4@տ�Ǻ�!?������@���{�ٿ��u3Oe�@ʙ�߮4@տ�Ǻ�!?������@hv�	�ٿS��@Aca�4@������!?|��#���@hv�	�ٿS��@Aca�4@������!?|��#���@�j�F�ٿfq�=���@���"�4@Tu:r�!?/�`S��@�j�F�ٿfq�=���@���"�4@Tu:r�!?/�`S��@�j�F�ٿfq�=���@���"�4@Tu:r�!?/�`S��@�j�F�ٿfq�=���@���"�4@Tu:r�!?/�`S��@��ٿ�Af���@����4@ �Ք�!?��m�c��@��ٿ�Af���@����4@ �Ք�!?��m�c��@^GE�ٿ�ُ�w�@"�'4@�RsQ
�!?�Y"0���@^GE�ٿ�ُ�w�@"�'4@�RsQ
�!?�Y"0���@^GE�ٿ�ُ�w�@"�'4@�RsQ
�!?�Y"0���@^GE�ٿ�ُ�w�@"�'4@�RsQ
�!?�Y"0���@W�Jߛ�ٿ�V6ئ �@����4@��R�!?!3�b��@W�Jߛ�ٿ�V6ئ �@����4@��R�!?!3�b��@W�Jߛ�ٿ�V6ئ �@����4@��R�!?!3�b��@W�Jߛ�ٿ�V6ئ �@����4@��R�!?!3�b��@W�Jߛ�ٿ�V6ئ �@����4@��R�!?!3�b��@����ٿ׬��e�@jVk��4@[(F/��!?����_&�@����ٿ׬��e�@jVk��4@[(F/��!?����_&�@����ٿ׬��e�@jVk��4@[(F/��!?����_&�@B����|ٿ^p����@Hqџ�4@.�X�\�!?�1�"�1�@���w�~ٿ���.���@#�4o4@a`�Ԑ!?Fh����@�T7]�ٿ�,d[��@�s��4@�L�Ai�!?+Z��9��@�T7]�ٿ�,d[��@�s��4@�L�Ai�!?+Z��9��@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@l)V�A�ٿ2��x��@T���4@�����!?��w�@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@�e�Ƀٿ�˻x��@.Wɡ4@�+)g��!?uPS��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@꽵r~ٿ��R"��@Z5��4@�hp5�!?y�{U}��@�P��Nٿ �>����@�Q5�4@+y��t�!?��Y���@�P��Nٿ �>����@�Q5�4@+y��t�!?��Y���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@�( ���ٿ_x����@A<vKw4@��q���!?���.���@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����%�ٿ����y��@#�W��4@	�*���!?��|�Q��@����W�ٿ��]H�@& ���4@>9���!?4����@#�	#��ٿS��/w��@=i>�4@��< �!?�.&#��@#�	#��ٿS��/w��@=i>�4@��< �!?�.&#��@#�	#��ٿS��/w��@=i>�4@��< �!?�.&#��@#�	#��ٿS��/w��@=i>�4@��< �!?�.&#��@#�	#��ٿS��/w��@=i>�4@��< �!?�.&#��@����~ٿ�Q�X���@��V4@�z�Đ!?��|��@?M�ٿ�E�@�I�S4@�ncܐ!?"�`�@?M�ٿ�E�@�I�S4@�ncܐ!?"�`�@?M�ٿ�E�@�I�S4@�ncܐ!?"�`�@?M�ٿ�E�@�I�S4@�ncܐ!?"�`�@?M�ٿ�E�@�I�S4@�ncܐ!?"�`�@�ԸkK{ٿ��+���@2@j�b4@�A7���!?- ޣ��@�ԸkK{ٿ��+���@2@j�b4@�A7���!?- ޣ��@�ԸkK{ٿ��+���@2@j�b4@�A7���!?- ޣ��@�*�6!}ٿCI��-�@j4�4i4@���~?�!?������@�*�6!}ٿCI��-�@j4�4i4@���~?�!?������@�*�6!}ٿCI��-�@j4�4i4@���~?�!?������@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@ ��\��ٿ+�.�-�@;�t�
4@��yC)�!?�^�O���@T���
zٿ��z����@�?�4@;�h��!?�=�
���@*
;�}ٿ ��xE�@�Q\�d4@3���!?���O�@*
;�}ٿ ��xE�@�Q\�d4@3���!?���O�@;u���ٿуTd�h�@O���4@�R_68�!?/0�]w�@;u���ٿуTd�h�@O���4@�R_68�!?/0�]w�@;u���ٿуTd�h�@O���4@�R_68�!?/0�]w�@;u���ٿуTd�h�@O���4@�R_68�!?/0�]w�@x�n���ٿ?VA����@���-4@RS�:�!?������@�Q���ٿO�P�ҟ�@�{�4@��7�!?�Q��Q,�@np��ٿ�6?�l��@ޗ"��4@��+��!?�4���@np��ٿ�6?�l��@ޗ"��4@��+��!?�4���@np��ٿ�6?�l��@ޗ"��4@��+��!?�4���@np��ٿ�6?�l��@ޗ"��4@��+��!?�4���@np��ٿ�6?�l��@ޗ"��4@��+��!?�4���@�qHl�ٿE�sŰ�@4S�?H4@+u�!?h�ޣZ�@�qHl�ٿE�sŰ�@4S�?H4@+u�!?h�ޣZ�@�qHl�ٿE�sŰ�@4S�?H4@+u�!?h�ޣZ�@XN���ٿXjѱ��@�k���4@����!?RA{��@XN���ٿXjѱ��@�k���4@����!?RA{��@XN���ٿXjѱ��@�k���4@����!?RA{��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@fp�N�ٿ�z'�UE�@��+4@�3ܐ!?tF��b��@4pɣ�ٿ�oH��@\4@Z���ϐ!?%�8�@4pɣ�ٿ�oH��@\4@Z���ϐ!?%�8�@4pɣ�ٿ�oH��@\4@Z���ϐ!?%�8�@�J:	�ٿ�?\Q���@d ��m4@�)��ސ!?5�vw���@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@l���ٿ�Zw8���@F��4@��)�Ӑ!?�*F�b��@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@��1�ٿ��H 0�@�P���4@4x����!?Yu���W�@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@e���P�ٿ8�wK���@�54��4@NL��Ð!?A�?G}��@S ��ٿu��qd9�@!x�A4@����!?}T����@S ��ٿu��qd9�@!x�A4@����!?}T����@S ��ٿu��qd9�@!x�A4@����!?}T����@S ��ٿu��qd9�@!x�A4@����!?}T����@S ��ٿu��qd9�@!x�A4@����!?}T����@��Xs�ٿixQW��@d
�4@���y�!?�ϯ�0�@��Xs�ٿixQW��@d
�4@���y�!?�ϯ�0�@��Xs�ٿixQW��@d
�4@���y�!?�ϯ�0�@���y�ٿ�;"���@?�o.� 4@~E5��!?X%����@�(�q��ٿu�sV��@;ӐH 4@�K	�K�!?#K�a��@�(�q��ٿu�sV��@;ӐH 4@�K	�K�!?#K�a��@w�s�ٿ�HAZ���@a���4@
�T��!?=�'l�@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@��=xN�ٿ� ��C�@�E�ϡ4@���׊�!?�RRD��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@�i =Z�ٿ���F���@Hz��4@t~�ի�!?Vyo��@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@*��X�ٿ�����@Аo�4@��J��!?"��I7�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@��r;ٿ�t9�)�@���^4@5���!?+)t�QL�@���H�ٿ��fMק�@	�:5?4@�4���!?5c���@���H�ٿ��fMק�@	�:5?4@�4���!?5c���@���H�ٿ��fMק�@	�:5?4@�4���!?5c���@���H�ٿ��fMק�@	�:5?4@�4���!?5c���@���H�ٿ��fMק�@	�:5?4@�4���!?5c���@���ٿ��A��@0iF��4@Śkʐ!?�1|��@���ٿ��A��@0iF��4@Śkʐ!?�1|��@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@g�b�ٿ�y���@w|��4@2<�=Ґ!?�� �%�@ԑ1�ٿ�u2��@XB]W�4@w��!?�
�,^��@ԑ1�ٿ�u2��@XB]W�4@w��!?�
�,^��@ԑ1�ٿ�u2��@XB]W�4@w��!?�
�,^��@ԑ1�ٿ�u2��@XB]W�4@w��!?�
�,^��@��A��ٿ��;9���@l l�& 4@�����!?��ْ��@��A��ٿ��;9���@l l�& 4@�����!?��ْ��@��A��ٿ��;9���@l l�& 4@�����!?��ْ��@��A��ٿ��;9���@l l�& 4@�����!?��ْ��@eF�V�ٿ&Sſ��@Z!6� 4@��3���!?�RY����@eF�V�ٿ&Sſ��@Z!6� 4@��3���!?�RY����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@�+�P�ٿ�� �١�@�Þ�4@8����!?a�a����@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@b��]{�ٿ�r؋s�@~��14@��Ђ��!?�[U���@�-8��ٿ��|�<u�@�t�4@q�GZ��!?��T���@�-8��ٿ��|�<u�@�t�4@q�GZ��!?��T���@]��qٿI��H�I�@xZ�2�4@٤�}�!?,PF����@�(�d�ٿ�cZ��y�@��[��4@G���q�!?��c�=��@�(�d�ٿ�cZ��y�@��[��4@G���q�!?��c�=��@�(�d�ٿ�cZ��y�@��[��4@G���q�!?��c�=��@�(�d�ٿ�cZ��y�@��[��4@G���q�!?��c�=��@T!��J�ٿހ�0d��@����4@�mB�ؐ!?�T�Y��@T!��J�ٿހ�0d��@����4@�mB�ؐ!?�T�Y��@T!��J�ٿހ�0d��@����4@�mB�ؐ!?�T�Y��@���ٿ��z��@�$�4@O)�!��!?��Sg���@���ٿ��z��@�$�4@O)�!��!?��Sg���@���ٿ��z��@�$�4@O)�!��!?��Sg���@���ٿ��z��@�$�4@O)�!��!?��Sg���@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@k��r]�ٿ4�ۙ���@t�0k4@�.���!?s0z�C�@m��Cg�ٿ�P�����@'_,�4@�3>�Ȑ!?sZ�ʨ��@m��Cg�ٿ�P�����@'_,�4@�3>�Ȑ!?sZ�ʨ��@m��Cg�ٿ�P�����@'_,�4@�3>�Ȑ!?sZ�ʨ��@~�pz�ٿOAv˯�@`���4@�S�!?��e K�@~�pz�ٿOAv˯�@`���4@�S�!?��e K�@~�pz�ٿOAv˯�@`���4@�S�!?��e K�@~�pz�ٿOAv˯�@`���4@�S�!?��e K�@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@�!�{�ٿ��KQ��@��R��4@��N?��!?��CL��@A���ٿ��g&i�@����W4@6SS���!?P�o�r�@�����ٿ�I����@SG�ٛ4@Ϧ�}�!?~�j=c�@���s�ٿ�l��42�@p)DZ4@N�R��!?��U�T�@��c�(�ٿֲ4��T�@�%�Q4@�='�X�!?�ޫ,�@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@3T����ٿޞ<U*�@/ӐLI4@Y�T�}�!?�G��>��@�~����ٿa�ώ��@���)4@��s��!?
>�f���@���c��ٿ��g;���@�m�8�4@6wAh��!?2��+_��@���c��ٿ��g;���@�m�8�4@6wAh��!?2��+_��@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�~@�ٿ=�r�i��@>x�74@�;⟐!?Q���D�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�y�ٿ������@�x�6�4@�/�ِ!?&�S-r�@�uC@�ٿ�((.�@;7^��4@�Q��!?��N\�)�@�uC@�ٿ�((.�@;7^��4@�Q��!?��N\�)�@�uC@�ٿ�((.�@;7^��4@�Q��!?��N\�)�@�uC@�ٿ�((.�@;7^��4@�Q��!?��N\�)�@�т���ٿ���:4�@ʯ(�D4@{�i��!?����z�@�т���ٿ���:4�@ʯ(�D4@{�i��!?����z�@�C�3t�ٿ^�D�Q�@OE�/n4@�Ȑ!?���醩�@�C�3t�ٿ^�D�Q�@OE�/n4@�Ȑ!?���醩�@�A=[�ٿ46��N�@b�_u4@gynX��!?�-~�4��@Wv�V�ٿ�:P�:��@+�X7Z4@��rؐ!?�Pk���@Wv�V�ٿ�:P�:��@+�X7Z4@��rؐ!?�Pk���@Wv�V�ٿ�:P�:��@+�X7Z4@��rؐ!?�Pk���@Wv�V�ٿ�:P�:��@+�X7Z4@��rؐ!?�Pk���@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@[q��)ٿ��!�g�@�g"� 4@<�*Ϣ�!?��kZ�@���~�ٿ;s��C�@���iQ4@<�9��!?�G�3	O�@���~�ٿ;s��C�@���iQ4@<�9��!?�G�3	O�@������ٿ�0���@��e�4@�9.̐!?��"���@ �U]�ٿ��iȠF�@2	4@��#⌐!?�u�2�
�@ �U]�ٿ��iȠF�@2	4@��#⌐!?�u�2�
�@ �U]�ٿ��iȠF�@2	4@��#⌐!?�u�2�
�@�XK�E�ٿ��8pK�@�qzs4@�湱��!?g��ϭ��@\�a�ٿ)F�9���@�{߀4@�u��!?��䭢U�@����}�ٿ��Wso��@���)74@�t!�U�!?yO*em�@/�#�ٿ�� �5��@�H=E�4@��-dh�!?�@��O�@/�#�ٿ�� �5��@�H=E�4@��-dh�!?�@��O�@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@��U�ٿ`܃8�@��7�4@���S|�!?.B�2���@ԍ��z�ٿ%l�F��@�7��4@�{�ސ!?J��q+s�@b���8�ٿe�>T~�@���?4@��G;�!?9�̣s��@b���8�ٿe�>T~�@���?4@��G;�!?9�̣s��@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@���2�ٿ��'q�^�@�@�4@4����!?��l�8�@�[H��ٿ��U{m�@"�HХ4@�E��!?�����d�@M�h�(�ٿ1r���@�}݅4@9�Y�!?�t���@-�Կ�ٿ��ت��@��<�4@��j�!?��L���@-�Կ�ٿ��ت��@��<�4@��j�!?��L���@-�Կ�ٿ��ت��@��<�4@��j�!?��L���@-�Կ�ٿ��ت��@��<�4@��j�!?��L���@-�Կ�ٿ��ت��@��<�4@��j�!?��L���@QZ;'��ٿ�GD)���@d+��4@���GI�!?D��3�@�B�ڒ�ٿk��sB��@)�΂�4@P�ah�!?aJ�jM��@���]�ٿ���(��@�
!34@]�Yk��!?����׻�@���]�ٿ���(��@�
!34@]�Yk��!?����׻�@�bU�^�ٿ�W�����@��4@��ė{�!?9 �Bf�@�bU�^�ٿ�W�����@��4@��ė{�!?9 �Bf�@y�v�ٿ�W�]���@:0��94@6�Z�`�!?�	�D@�@y�v�ٿ�W�]���@:0��94@6�Z�`�!?�	�D@�@y�v�ٿ�W�]���@:0��94@6�Z�`�!?�	�D@�@�?�ٿ�3m���@ߚ��A4@km�_�!?eyRvO[�@�?�ٿ�3m���@ߚ��A4@km�_�!?eyRvO[�@�?�ٿ�3m���@ߚ��A4@km�_�!?eyRvO[�@�?�ٿ�3m���@ߚ��A4@km�_�!?eyRvO[�@�?�ٿ�3m���@ߚ��A4@km�_�!?eyRvO[�@��~�~~ٿ(�w65�@._�F 4@H
;���!?����@��@��~�~~ٿ(�w65�@._�F 4@H
;���!?����@��@?�ӓ|ٿ���%���@�����4@�pW*Ȑ!?��}L���@?�ӓ|ٿ���%���@�����4@�pW*Ȑ!?��}L���@?�ӓ|ٿ���%���@�����4@�pW*Ȑ!?��}L���@��c눆ٿ�
�PEo�@��+`4@2�ِ!?_�ZF5j�@��c눆ٿ�
�PEo�@��+`4@2�ِ!?_�ZF5j�@��c눆ٿ�
�PEo�@��+`4@2�ِ!?_�ZF5j�@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@>b��L�ٿ�~�n0V�@����4@�V��!?WY�& ��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@�7��=�ٿ�\`��@<��[4@��Wm�!?;2l>M��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@��7�ٿ��_׷��@�(a�k4@OQؐ!?���[h��@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@c.�eӇٿ,&m��@ܙ���4@RC��!?�C�\�q�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@D�f렃ٿ�����@�p!]
4@�+E�!?D":�d�@ 8�V�ٿ��q��@��Ƚ�4@T�| ��!?�XI߿��@F���ٿ�P=����@��4�4@3�)o��!?]@���@F���ٿ�P=����@��4�4@3�)o��!?]@���@F���ٿ�P=����@��4�4@3�)o��!?]@���@�5A���ٿg8��n��@K ��4@�s�.�!?���R��@���=�ٿ�w����@�F5"D4@I�Ϙ�!?�v'=6�@���=�ٿ�w����@�F5"D4@I�Ϙ�!?�v'=6�@���=�ٿ�w����@�F5"D4@I�Ϙ�!?�v'=6�@D�l��ٿ��v&Ċ�@�g��4@��m��!?h��-��@D�l��ٿ��v&Ċ�@�g��4@��m��!?h��-��@� Ï�ٿаkBq��@ϩt^�4@;����!?�N�WV�@� Ï�ٿаkBq��@ϩt^�4@;����!?�N�WV�@� Ï�ٿаkBq��@ϩt^�4@;����!?�N�WV�@%�/��ٿƂ����@��@�4@Pcf�r�!?�Pƽ�k�@wǴS:�ٿf�;���@!�j4@�4�P^�!?�S�r��@wǴS:�ٿf�;���@!�j4@�4�P^�!?�S�r��@wǴS:�ٿf�;���@!�j4@�4�P^�!?�S�r��@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@�9�ٿ~��d6�@��x	I4@	�G䯐!?;�vz0�@i�ϕ�ٿwRղ�J�@rE#�4@B����!?�iɻy�@i�ϕ�ٿwRղ�J�@rE#�4@B����!?�iɻy�@�!����ٿ��KL���@��ne4@&��Ր!?�W���@��J��ٿM�R�O<�@�1��
4@G	�i�!?z�|��f�@��J��ٿM�R�O<�@�1��
4@G	�i�!?z�|��f�@٪L���ٿJ�6����@�rTa4@}I����!?\�
��@٪L���ٿJ�6����@�rTa4@}I����!?\�
��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@5�-I��ٿ�&O��p�@RN�/4@����!?[9X3��@��$�ٿ�H�bt�@�lL�2	4@݁���!?�IL��@�@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p��9�ٿ�ﶾ
��@�J�4@�p�`v�!?&s��@p1�ٿ
��r0��@�v$�4@�nP��!?�͐]6��@p1�ٿ
��r0��@�v$�4@�nP��!?�͐]6��@p1�ٿ
��r0��@�v$�4@�nP��!?�͐]6��@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@��QZ�ٿ@��m���@NN�`4@78�V��!?�@T�%�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@=��`C�ٿve��Q�@u���4@0ː!?��(�E�@��B���ٿ�Xbv*��@/���q4@AH�!?H���ݶ�@K�(�e�ٿ�)�T��@���� 4@�E��!?��+���@K�(�e�ٿ�)�T��@���� 4@�E��!?��+���@K�(�e�ٿ�)�T��@���� 4@�E��!?��+���@K�(�e�ٿ�)�T��@���� 4@�E��!?��+���@�a��ٿ�]*�:�@��R4@��$q�!?�K�,���@�a��ٿ�]*�:�@��R4@��$q�!?�K�,���@i��ˀٿ��i����@L�M��4@ԗ��!?�}�
��@i��ˀٿ��i����@L�M��4@ԗ��!?�}�
��@��C��ٿZEQ�g��@��I�4@�?.�!?չAu��@��Uڑٿ��j��@6�㠒4@͸��Ð!?�	E ���@�n�x��ٿ7&{!���@R��f4@@ܼ�Ӑ!?sO�k��@�n�x��ٿ7&{!���@R��f4@@ܼ�Ӑ!?sO�k��@�a7[��ٿ}�)�Al�@N�u4@���Ґ!?�C�p�P�@�a7[��ٿ}�)�Al�@N�u4@���Ґ!?�C�p�P�@�a7[��ٿ}�)�Al�@N�u4@���Ґ!?�C�p�P�@�a7[��ٿ}�)�Al�@N�u4@���Ґ!?�C�p�P�@���҇ٿ�O:K��@�J-�4@����!?�ƚyb�@���҇ٿ�O:K��@�J-�4@����!?�ƚyb�@���҇ٿ�O:K��@�J-�4@����!?�ƚyb�@���҇ٿ�O:K��@�J-�4@����!?�ƚyb�@+����ٿ �]����@����F4@�A|��!?Ya]�{��@+����ٿ �]����@����F4@�A|��!?Ya]�{��@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@��+��ٿ�Rh"q�@�9��j4@�Kf���!?Q���3_�@}b�{��ٿ�f�?���@Qګ�}4@�ڒ��!?�����@}b�{��ٿ�f�?���@Qګ�}4@�ڒ��!?�����@}b�{��ٿ�f�?���@Qګ�}4@�ڒ��!?�����@}b�{��ٿ�f�?���@Qګ�}4@�ڒ��!?�����@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@ϕ��q�ٿ�Y�*�@�;���4@r4C��!?���1��@��f�ʆٿ��GNk�@O��W
4@�F���!?}�kO�2�@��f�ʆٿ��GNk�@O��W
4@�F���!?}�kO�2�@��f�ʆٿ��GNk�@O��W
4@�F���!?}�kO�2�@$�og}ٿv�ā�9�@+� 4@����!?��,�/��@$�og}ٿv�ā�9�@+� 4@����!?��,�/��@<.�|ٿ��U�@.Y�4@Hv�Ð!?�(�����@<.�|ٿ��U�@.Y�4@Hv�Ð!?�(�����@-3�� �ٿ�E��@���P�	4@LX��!?��z�bg�@� �M�ٿLo�����@d�NZ4@�:F�!?ɉG&X_�@���ٿ��/�e�@��Ű�4@@� T�!?�N�!��@���ٿ��/�e�@��Ű�4@@� T�!?�N�!��@���ٿ��/�e�@��Ű�4@@� T�!?�N�!��@b.�[�ٿMl��0b�@"f�6�4@�*�'�!?�z�e#�@b.�[�ٿMl��0b�@"f�6�4@�*�'�!?�z�e#�@b.�[�ٿMl��0b�@"f�6�4@�*�'�!?�z�e#�@����ٿN?k�W�@�U�\�4@ި�.א!?j�#�j�@����ٿN?k�W�@�U�\�4@ި�.א!?j�#�j�@����ٿN?k�W�@�U�\�4@ި�.א!?j�#�j�@����ٿN?k�W�@�U�\�4@ި�.א!?j�#�j�@����ٿN?k�W�@�U�\�4@ި�.א!?j�#�j�@�Ke>�ٿ��]�N�@#�zS4@dX'�ː!?���/@��@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@F�-�-�ٿ�q����@�D�4@,\3Ň�!?7����@|���&�ٿ9�����@eC��4@*����!?(��t��@|���&�ٿ9�����@eC��4@*����!?(��t��@|���&�ٿ9�����@eC��4@*����!?(��t��@|���&�ٿ9�����@eC��4@*����!?(��t��@�8�~�ٿ��D"���@(�k4@5m,5j�!?�!
���@�8�~�ٿ��D"���@(�k4@5m,5j�!?�!
���@G�3��ٿ�r�K���@zr�כ4@�!�!?ɨ�O��@G�3��ٿ�r�K���@zr�כ4@�!�!?ɨ�O��@G�3��ٿ�r�K���@zr�כ4@�!�!?ɨ�O��@,wڄٿx+vP��@�G��4@
t��}�!?�"����@,wڄٿx+vP��@�G��4@
t��}�!?�"����@,wڄٿx+vP��@�G��4@
t��}�!?�"����@,wڄٿx+vP��@�G��4@
t��}�!?�"����@,wڄٿx+vP��@�G��4@
t��}�!?�"����@01P@�|ٿ�!6L�L�@�4DW4@n��H��!?U3�=�P�@01P@�|ٿ�!6L�L�@�4DW4@n��H��!?U3�=�P�@ŋ�Km�ٿ��~Aj�@�Nֆ4@�ѓ	��!?����'��@ŋ�Km�ٿ��~Aj�@�Nֆ4@�ѓ	��!?����'��@ŋ�Km�ٿ��~Aj�@�Nֆ4@�ѓ	��!?����'��@�ٿ�4��RG�@��|�4@�(�ހ�!?v��c=��@9I��ٿ]!��E�@%ޑ��	4@�{+q��!?��7��@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@Sk���ٿ�k���@��/UY4@0Ҕp��!?2`1 2�@���R��ٿ9��oT�@O�F�c4@���ې!?fV�~k'�@A�mY��ٿ��;$)��@��i�4@�}�Z��!?T�|\��@A�mY��ٿ��;$)��@��i�4@�}�Z��!?T�|\��@�ٿYA�1!��@���2�4@���ᦐ!? X�%��@�ٿYA�1!��@���2�4@���ᦐ!? X�%��@�ٿYA�1!��@���2�4@���ᦐ!? X�%��@�ٿYA�1!��@���2�4@���ᦐ!? X�%��@���i��ٿ��d$�@�z�4@�8X��!?߄�o���@���i��ٿ��d$�@�z�4@�8X��!?߄�o���@���i��ٿ��d$�@�z�4@�8X��!?߄�o���@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@2%���ٿg�]�[��@�$u�4@9�:��!?Y�!T�"�@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@���s�ٿH��u��@�X�%4@v����!?�� ���@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@����ٿZ(n�ڬ�@T�	�4@�I�탐!?Tu����@r��H��ٿ�����@6!	Y�4@�u�M��!?�ź����@r��H��ٿ�����@6!	Y�4@�u�M��!?�ź����@r��H��ٿ�����@6!	Y�4@�u�M��!?�ź����@r��H��ٿ�����@6!	Y�4@�u�M��!?�ź����@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@D����ٿ��A��@����4@�l��ߐ!?���B��@a�����ٿ���̌��@�_�Ð4@)v����!?E�9Hxh�@�V��m�ٿ�;����@ȗH�4@����!?�E�=���@�V��m�ٿ�;����@ȗH�4@����!?�E�=���@�V��m�ٿ�;����@ȗH�4@����!?�E�=���@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@~��M�ٿ�iQ����@����A4@FO�&֐!?;�3�@��(h�ٿ���]p��@+���=4@{�5��!?�q�6u�@��(h�ٿ���]p��@+���=4@{�5��!?�q�6u�@��(h�ٿ���]p��@+���=4@{�5��!?�q�6u�@��(h�ٿ���]p��@+���=4@{�5��!?�q�6u�@�S�D�ٿ�X����@w7�^4@��R8�!?٠i|���@&7�~ٿe嫩/�@z��Bs4@ģ���!?˷�ɝ�@G'�UE�ٿ<÷Y��@[��F4@�M5�S�!?��3w^,�@fX�ٿs'ܼ��@խ�>;4@���!?7,ҍI��@j�ȉшٿ��z6e��@UB��x4@\[gΐ!?�vs�.�@j�ȉшٿ��z6e��@UB��x4@\[gΐ!?�vs�.�@j�ȉшٿ��z6e��@UB��x4@\[gΐ!?�vs�.�@j�ȉшٿ��z6e��@UB��x4@\[gΐ!?�vs�.�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@t��#�ٿ���3���@ �O��4@D�Ƽ��!?�)��u�@Pⁿ�ٿ��y!c�@\Ou�4@T�]��!?�O��$�@Pⁿ�ٿ��y!c�@\Ou�4@T�]��!?�O��$�@.�lD��ٿ��<�d�@ȣ({4@u�� �!?���r��@.�lD��ٿ��<�d�@ȣ({4@u�� �!?���r��@.�lD��ٿ��<�d�@ȣ({4@u�� �!?���r��@�؄/��ٿ���&\��@<q{4@�v�H�!?�K����@�؄/��ٿ���&\��@<q{4@�v�H�!?�K����@�؄/��ٿ���&\��@<q{4@�v�H�!?�K����@�؄/��ٿ���&\��@<q{4@�v�H�!?�K����@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@K�E��ٿ��R���@ ,�<�4@:p�!?��pHZ�@CLc��ٿ��.��H�@�4@�@k��!?�/9����@CLc��ٿ��.��H�@�4@�@k��!?�/9����@CLc��ٿ��.��H�@�4@�@k��!?�/9����@CLc��ٿ��.��H�@�4@�@k��!?�/9����@CLc��ٿ��.��H�@�4@�@k��!?�/9����@CLc��ٿ��.��H�@�4@�@k��!?�/9����@Q� �ٿ�Ѻ�)�@_C���4@��n�!?��T�@Q� �ٿ�Ѻ�)�@_C���4@��n�!?��T�@����ٿ�M@q�<�@c1d�4@��x��!?��-�=�@~l�nk�ٿ�<���@�(�4@`�aԆ�!?6ndXr�@gܤŇٿOM�Q��@c���4@�&�t��!?h�|ilV�@-b$�1�ٿd�cw_��@X5���4@/�%ڂ�!?�[vCC��@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@.�cd�ٿ)�����@.-J�4@��腐!?l��z�@���(ܐٿc�l̩�@��G�4@�!-��!?�>����@���(��ٿ���.���@��^4@(0vw��!?�봴���@���(��ٿ���.���@��^4@(0vw��!?�봴���@��ٿ�������@��A�4@͂$Ĉ�!?s00�@��ٿ�������@��A�4@͂$Ĉ�!?s00�@��ٿ�������@��A�4@͂$Ĉ�!?s00�@��ٿ�������@��A�4@͂$Ĉ�!?s00�@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@:q9`��ٿ0�
����@�U�ղ4@d��!?���ך��@K���ٿ 7�v�@�?kc�4@��怐!?ܴ��@K���ٿ 7�v�@�?kc�4@��怐!?ܴ��@K���ٿ 7�v�@�?kc�4@��怐!?ܴ��@K���ٿ 7�v�@�?kc�4@��怐!?ܴ��@K���ٿ 7�v�@�?kc�4@��怐!?ܴ��@]E�~ٿ٧V���@���Ln4@I^kX��!?UP���@]E�~ٿ٧V���@���Ln4@I^kX��!?UP���@]E�~ٿ٧V���@���Ln4@I^kX��!?UP���@�R�nٿ�k���@��� �	4@��z���!?��e�w��@�R�nٿ�k���@��� �	4@��z���!?��e�w��@�R�nٿ�k���@��� �	4@��z���!?��e�w��@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@��Rښ�ٿ��i&��@v��I4@�s�ϐ!?�&�%y�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@O��G�ٿJ����@�@��0��4@�5�ݙ�!?�� �jr�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@��^$܅ٿ�}�S��@^d��4@!Y:�ِ!?�ܪ�;�@,ga��ٿ�X<�:�@�����4@��4s�!?r���q�@�����ٿ|�u�@Ŧ�S4@vEξ�!?�,���@�&G�P�ٿ��1hq��@����B4@����!?�8��@�&G�P�ٿ��1hq��@����B4@����!?�8��@��-c�ٿ���iq�@�6Jw{4@��Nޚ�!?s�֣(�@��b��ٿ���,��@�vH4@;���ː!?���.���@��b��ٿ���,��@�vH4@;���ː!?���.���@��b��ٿ���,��@�vH4@;���ː!?���.���@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@�f�B��ٿ|������@�XÔ4@�z�6{�!?��UhN��@^���J�ٿϑ)r��@ۇE4@�j��z�!?y�M�@��t/�ٿMn�`�@��/��4@���Ґ!?��	����@��t/�ٿMn�`�@��/��4@���Ґ!?��	����@��t/�ٿMn�`�@��/��4@���Ґ!?��	����@ ).��ٿƭ��@)ݺ�-4@t��w(�!?�F�(�@ ).��ٿƭ��@)ݺ�-4@t��w(�!?�F�(�@ ).��ٿƭ��@)ݺ�-4@t��w(�!?�F�(�@��Ì�ٿq��N�@���˖4@=oje̐!?�����@��Ì�ٿq��N�@���˖4@=oje̐!?�����@靝��ٿ�q�C�@�(x�:4@vHx(�!?���I���@靝��ٿ�q�C�@�(x�:4@vHx(�!?���I���@4L�R�ٿ ��h@�@��q� 4@Sł�Ր!?<��`�@�H���ٿ�lw���@��ވ� 4@C�آ>�!?V�'؉!�@����ٿ�����@���"4@2xwҐ!?��QW��@����ٿ�����@���"4@2xwҐ!?��QW��@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@t�)�~�ٿ~�p�I��@$�近 4@�(9��!?#ŇM�4�@~N	�ʋٿ
���dI�@E3�%4@_c+��!?@�{M/��@~N	�ʋٿ
���dI�@E3�%4@_c+��!?@�{M/��@~N	�ʋٿ
���dI�@E3�%4@_c+��!?@�{M/��@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@t��7�ٿ����E��@7ʞɭ4@f��ِ!?U}�_)�@ޒ�䏉ٿ��2��@�|�Q�4@{�V��!?���h��@ޒ�䏉ٿ��2��@�|�Q�4@{�V��!?���h��@ޒ�䏉ٿ��2��@�|�Q�4@{�V��!?���h��@ޒ�䏉ٿ��2��@�|�Q�4@{�V��!?���h��@ޒ�䏉ٿ��2��@�|�Q�4@{�V��!?���h��@��ԙ	�ٿ>I�
�@�s V�4@IG^y��!?#�����@��ԙ	�ٿ>I�
�@�s V�4@IG^y��!?#�����@��ԙ	�ٿ>I�
�@�s V�4@IG^y��!?#�����@�?���ٿ�4�!{��@���4@�(��Ȑ!?W�\��O�@�?���ٿ�4�!{��@���4@�(��Ȑ!?W�\��O�@�?���ٿ�4�!{��@���4@�(��Ȑ!?W�\��O�@KQ��g�ٿ?]�e<*�@�#�9E4@FH��ِ!?�K��L�@	�B�6�ٿ��g����@|%R�	4@7^Jj�!?~ⲱ�#�@	�B�6�ٿ��g����@|%R�	4@7^Jj�!?~ⲱ�#�@�p^�ƌٿ�#�z�r�@o��4@�~7�O�!?�Jŷ�@"���ٿHw���@�����4@��r�A�!?���y���@"���ٿHw���@�����4@��r�A�!?���y���@�P�ۍٿ4�A��@���$4@��3�Ð!?�>�g�<�@�P�ۍٿ4�A��@���$4@��3�Ð!?�>�g�<�@�P�ۍٿ4�A��@���$4@��3�Ð!?�>�g�<�@@���q�ٿ:P'�A��@�#/4@kr$ِ!?s�j��@�*:؛�ٿ����l��@�Z�R%4@b���!?W�	��D�@�*:؛�ٿ����l��@�Z�R%4@b���!?W�	��D�@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@G���ٿ�vTn�W�@3��^4@����!?�С:���@�f�Јٿ�Q�P��@���
4@�����!?�ʃ��@���沁ٿ%%�)f��@ۮ��	4@�V�Fא!?�IS��F�@���沁ٿ%%�)f��@ۮ��	4@�V�Fא!?�IS��F�@���沁ٿ%%�)f��@ۮ��	4@�V�Fא!?�IS��F�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@ո}
�ٿ�>��L�@r�˄�4@	q���!?�7�_v�@.i�g�ٿH"1y"��@���a�4@��/ː!?�s[����@.i�g�ٿH"1y"��@���a�4@��/ː!?�s[����@.i�g�ٿH"1y"��@���a�4@��/ː!?�s[����@.i�g�ٿH"1y"��@���a�4@��/ː!?�s[����@.i�g�ٿH"1y"��@���a�4@��/ː!?�s[����@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@�|}��~ٿV��'��@l{��4@3�J���!?r%p���@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@���$ٿ���`��@��(� 4@�[��͐!?c�D�N}�@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@$���E�ٿ
�<�p�@6�zf4@e� f��!?��H���@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@;�����ٿ����`�@�Av�4@�<ʮ�!?^� �CG�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@+��褁ٿJ*ظ���@�lCS4@�b���!?��Y�]�@�dVe>�ٿջ�%f��@�
�4@#_���!?���Õ��@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@��΀ٿ�j����@��84@Q�ѐ!?��D(6�@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@�E��ٿʒC����@�o���4@�N�QՐ!?�b� ���@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@��c�0�ٿ׮���	�@^ϕ84@Ca����!?�a��u�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@�>`�ٿ�s����@$^K}4@�}��!?-����@�@����ٿܓq����@X&�h+4@���K�!?Z�x�#��@����ٿܓq����@X&�h+4@���K�!?Z�x�#��@��t�
�ٿ��x���@nz��
4@��:��!?�xt��b�@#[<�g�ٿkڲ7�@��Q�'4@D�;}�!?PB�\��@��2?&�ٿ�)4���@&j$�	4@0#ҵ�!?���O,��@��2?&�ٿ�)4���@&j$�	4@0#ҵ�!?���O,��@Np1���ٿ�A��ko�@��y��4@�㆞Ґ!?Ø�?��@%B]�O�ٿyfD�g�@���U�4@υR\��!?�Ҋ8�^�@I�����ٿ��ܗ��@
��j4@���ߐ!?�������@I�����ٿ��ܗ��@
��j4@���ߐ!?�������@I�����ٿ��ܗ��@
��j4@���ߐ!?�������@I�����ٿ��ܗ��@
��j4@���ߐ!?�������@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@��5�τٿ�1�c��@����Y4@��d�!?<�?)��@~��o�ٿ(��|0��@_�&�4@�a����!?���ɖ�@~��o�ٿ(��|0��@_�&�4@�a����!?���ɖ�@�����ٿ�Z'�e��@�m���4@ΦE�!?a��kd�@~��݄ٿbS�-��@JV�x4@.rE��!?�;�a���@~��݄ٿbS�-��@JV�x4@.rE��!?�;�a���@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��B���ٿ�"��E
�@TQ���4@��E�ǐ!?���Z*�@��1삄ٿ�{`vE�@Եd(�	4@�ʐ!?M>O�@��1삄ٿ�{`vE�@Եd(�	4@�ʐ!?M>O�@���A��ٿ��qކ�@���	4@ƙ�Dv�!?iy�����@���A��ٿ��qކ�@���	4@ƙ�Dv�!?iy�����@���A��ٿ��qކ�@���	4@ƙ�Dv�!?iy�����@���A��ٿ��qކ�@���	4@ƙ�Dv�!?iy�����@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@j�C��ٿ ����@g��=4@}�7�[�!?y��R�%�@���]"�ٿ����5�@Ÿ4@	�$xp�!?跸5��@���]"�ٿ����5�@Ÿ4@	�$xp�!?跸5��@��j�g~ٿ�����@iw0v4@8���!?j�����@��j�g~ٿ�����@iw0v4@8���!?j�����@��j�g~ٿ�����@iw0v4@8���!?j�����@��j�g~ٿ�����@iw0v4@8���!?j�����@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@S؊�q�ٿ��9I,�@�梗I 4@=���͐!?N"�c���@�7i��}ٿ@�ߢv�@�_ʣ� 4@7EG���!?�R藕��@�7i��}ٿ@�ߢv�@�_ʣ� 4@7EG���!?�R藕��@�7i��}ٿ@�ߢv�@�_ʣ� 4@7EG���!?�R藕��@�7i��}ٿ@�ߢv�@�_ʣ� 4@7EG���!?�R藕��@�7i��}ٿ@�ߢv�@�_ʣ� 4@7EG���!?�R藕��@�
���ٿB��7a�@�ѳ5�4@�~��!?=�Vt�C�@�
���ٿB��7a�@�ѳ5�4@�~��!?=�Vt�C�@4�.k�ٿ��Ԁ	,�@l^��4@�{p޹�!?±5�=��@4�.k�ٿ��Ԁ	,�@l^��4@�{p޹�!?±5�=��@4�.k�ٿ��Ԁ	,�@l^��4@�{p޹�!?±5�=��@4�.k�ٿ��Ԁ	,�@l^��4@�{p޹�!?±5�=��@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�hA��ٿ y�@�E�@� ���4@��󀢐!?�[U�ϕ�@�|^���ٿ���g�\�@1�)i�4@sݧ�!?���V��@@���}�ٿ~E��\�@�NO
-4@����j�!? ����@@���}�ٿ~E��\�@�NO
-4@����j�!? ����@�6��:�ٿ�X��@V��#�4@?��n��!?���>��@ym�ٿ�RW���@�1c�4@d�����!?ؙ�g�O�@ym�ٿ�RW���@�1c�4@d�����!?ؙ�g�O�@ym�ٿ�RW���@�1c�4@d�����!?ؙ�g�O�@ym�ٿ�RW���@�1c�4@d�����!?ؙ�g�O�@ym�ٿ�RW���@�1c�4@d�����!?ؙ�g�O�@(�B��ٿS�\���@!��W4@)���̐!?������@(�B��ٿS�\���@!��W4@)���̐!?������@(�B��ٿS�\���@!��W4@)���̐!?������@(�B��ٿS�\���@!��W4@)���̐!?������@��&�ٿ5�6����@'�\ .4@9~���!?J�:�U��@��&�ٿ5�6����@'�\ .4@9~���!?J�:�U��@��&�ٿ5�6����@'�\ .4@9~���!?J�:�U��@��&�ٿ5�6����@'�\ .4@9~���!?J�:�U��@��`���ٿ�`(���@�8x�E4@�d����!?y@V���@��`���ٿ�`(���@�8x�E4@�d����!?y@V���@��`���ٿ�`(���@�8x�E4@�d����!?y@V���@��`���ٿ�`(���@�8x�E4@�d����!?y@V���@��`���ٿ�`(���@�8x�E4@�d����!?y@V���@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@&ؑI�ٿ�}���@,�� 4@��!x��!?μ����@���[��ٿ�{`����@�keX� 4@�(����!?9���V�@Ȏ��k�ٿ��eg(�@�>pk�4@�Mt���!?X	��д�@Ȏ��k�ٿ��eg(�@�>pk�4@�Mt���!?X	��д�@�}��ٿ �����@���4@S�Z��!?$����@�}��ٿ �����@���4@S�Z��!?$����@��TK��ٿ���4��@
ݺo4@"��ᗐ!?ы���@P�V��ٿ�<'1K�@�Wz#�4@_R�W�!?�d����@P�V��ٿ�<'1K�@�Wz#�4@_R�W�!?�d����@P�V��ٿ�<'1K�@�Wz#�4@_R�W�!?�d����@P�V��ٿ�<'1K�@�Wz#�4@_R�W�!?�d����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@�;v�|�ٿ�~����@�j��4@��^�!?�|�����@m+b�b�ٿ����R�@�V��4@<�<.\�!?�E���@m+b�b�ٿ����R�@�V��4@<�<.\�!?�E���@m+b�b�ٿ����R�@�V��4@<�<.\�!?�E���@m+b�b�ٿ����R�@�V��4@<�<.\�!?�E���@m+b�b�ٿ����R�@�V��4@<�<.\�!?�E���@`�7���ٿ�g�݆��@!���4@�����!?��:g_V�@`�7���ٿ�g�݆��@!���4@�����!?��:g_V�@`�7���ٿ�g�݆��@!���4@�����!?��:g_V�@`�7���ٿ�g�݆��@!���4@�����!?��:g_V�@�_+�D�ٿܷ��f�@JF�o�4@�͔�֐!?��ћ���@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@S��ٿ.���1_�@7l���4@��謢�!?��|/�@ݏvV|�ٿz�5�M��@��=w4@� �A��!?D%��t��@ݏvV|�ٿz�5�M��@��=w4@� �A��!?D%��t��@ݏvV|�ٿz�5�M��@��=w4@� �A��!?D%��t��@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@�^��m�ٿ��j=��@�X���4@M�dƐ!?R/To�@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@4�����ٿ����@I��4@L�*W�!?z֘���@瀌�ٿ�:�4�@!�C�4@���א!?�+�&F��@瀌�ٿ�:�4�@!�C�4@���א!?�+�&F��@瀌�ٿ�:�4�@!�C�4@���א!?�+�&F��@瀌�ٿ�:�4�@!�C�4@���א!?�+�&F��@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@aJwx�ٿBs�d���@�>Y4@8%��!?>."=�5�@-���ٿ	�k˂�@C$	L�4@n<�g7�!?qX�n�d�@-���ٿ	�k˂�@C$	L�4@n<�g7�!?qX�n�d�@-���ٿ	�k˂�@C$	L�4@n<�g7�!?qX�n�d�@�(;���ٿ�L�����@>�S�4@v&[2�!?DDV����@�ㆴs�ٿ �"��@iN04@F(���!?������@�ㆴs�ٿ �"��@iN04@F(���!?������@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�q�	�ٿ�tCf��@w�UV4@i�2��!?��Pɭ��@�����ٿV�a=�@���j�4@ZN�-��!?Hb�h��@�����ٿV�a=�@���j�4@ZN�-��!?Hb�h��@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@/O�>ʈٿ _J�1�@7g Y4@�����!?�#�c���@2��V �ٿ��)���@.���4@��Xг�!?��,��@2��V �ٿ��)���@.���4@��Xг�!?��,��@2��V �ٿ��)���@.���4@��Xг�!?��,��@:M��ٿ�I����@��\h4@+�K���!?�v� k�@:M��ٿ�I����@��\h4@+�K���!?�v� k�@:M��ٿ�I����@��\h4@+�K���!?�v� k�@:V�μ�ٿߴ�+��@f:$4@�?ȫ�!?�wD�qa�@:V�μ�ٿߴ�+��@f:$4@�?ȫ�!?�wD�qa�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@	��E�ٿ��$=��@]�˞�4@��ې!?@$��t�@r�Þ��ٿSK����@�r��4@�Lӎ�!?4��\=T�@r�Þ��ٿSK����@�r��4@�Lӎ�!?4��\=T�@���ٿ�۽v���@]vơ4@�$ꨐ!?�W+~���@���ٿ�۽v���@]vơ4@�$ꨐ!?�W+~���@���ٿ�۽v���@]vơ4@�$ꨐ!?�W+~���@o��8�ٿ�Y���@����B4@ouG��!?<l�Pyp�@d�E�ٿ������@�.U4@��Ö�!?���+�"�@d�E�ٿ������@�.U4@��Ö�!?���+�"�@�~��ٿ�L:�@o��@�4@.�ؐ!?D y5�!�@�~��ٿ�L:�@o��@�4@.�ؐ!?D y5�!�@�~��ٿ�L:�@o��@�4@.�ؐ!?D y5�!�@�`!	�ٿA�p���@h���4@_�M%�!?0�z���@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@<mݕ�ٿ4eǆ���@��>�34@��&�!?����o�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�Q嗲�ٿ�z�����@K�s4�4@O���!?�x/Q�<�@�<Xԉٿ��2uy�@�v�
�4@��Z���!?EJ���@�<Xԉٿ��2uy�@�v�
�4@��Z���!?EJ���@�<Xԉٿ��2uy�@�v�
�4@��Z���!?EJ���@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@SgvAY�ٿ��½��@Z�s��4@����!?�㏦x<�@���H��ٿ�]�Q7��@2�s]�4@�<��ʐ!?LH�[���@t�%�L�ٿ�l�Oz�@�a	Mm4@zN7��!?O1�	�W�@t�%�L�ٿ�l�Oz�@�a	Mm4@zN7��!?O1�	�W�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@�W�w�ٿ�v ��@:gK�4@e�\�!?���v3F�@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@瓡έ�ٿ�2���@{vʲ4@�"���!?��f����@�Cۈٿy`�0��@1O��>4@8�?}��!?s�M��@�Cۈٿy`�0��@1O��>4@8�?}��!?s�M��@�� m�ٿ�d�~j�@��m�14@$Ϭm�!?v�\V���@�.絋ٿ�PA�ŏ�@mб,�4@�k	✐!?_�g=��@�.絋ٿ�PA�ŏ�@mб,�4@�k	✐!?_�g=��@�.絋ٿ�PA�ŏ�@mб,�4@�k	✐!?_�g=��@�.絋ٿ�PA�ŏ�@mб,�4@�k	✐!?_�g=��@l���ٿwŴ���@ �+6�4@z��@ǐ!?`vG�0��@l���ٿwŴ���@ �+6�4@z��@ǐ!?`vG�0��@l���ٿwŴ���@ �+6�4@z��@ǐ!?`vG�0��@l���ٿwŴ���@ �+6�4@z��@ǐ!?`vG�0��@l���ٿwŴ���@ �+6�4@z��@ǐ!?`vG�0��@� S�ٿ�܍!���@~�*p�4@�(Z��!?�3H�<�@� S�ٿ�܍!���@~�*p�4@�(Z��!?�3H�<�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@���8��ٿ��\�� �@xCYy�4@,'�ϐ!?�[�&�@�1c?�ٿ�%Fח��@�ESE4@�Ӟ��!?�o߈��@�1c?�ٿ�%Fח��@�ESE4@�Ӟ��!?�o߈��@�1c?�ٿ�%Fח��@�ESE4@�Ӟ��!?�o߈��@�1c?�ٿ�%Fח��@�ESE4@�Ӟ��!?�o߈��@I�PY�ٿ�C�� ��@T3��:4@��@*�!?�p�Z��@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��	��ٿ���2��@ǟR4@@��o�!?��OoB�@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@��'ƣ�ٿ�����@bP�е4@��[א!?�)"���@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@Lw�K�ٿ.��.���@�zv�4@y�^㥐!?���8��@���;�ٿ��3�_g�@�!��Y4@�Ax-ϐ!?��JG��@=���A�ٿ�q�7%�@>�&�4@?]��ڐ!?�>����@AG����ٿ���,�@@�m��4@e��[�!?������@AG����ٿ���,�@@�m��4@e��[�!?������@���>�ٿ�X�\��@��q�4@7 ���!?�"�U�@���>�ٿ�X�\��@��q�4@7 ���!?�"�U�@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@�?z�ٿp�E0�i�@��ћ�4@�i���!?�G���@?�y7\�ٿ�N�My�@Ä���4@�_|�L�!?�+!g��@?�y7\�ٿ�N�My�@Ä���4@�_|�L�!?�+!g��@?�y7\�ٿ�N�My�@Ä���4@�_|�L�!?�+!g��@?�y7\�ٿ�N�My�@Ä���4@�_|�L�!?�+!g��@'?�8 �ٿ�lYYV�@�J��B4@V�X��!?�o��X�@'?�8 �ٿ�lYYV�@�J��B4@V�X��!?�o��X�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@ܹç@�ٿ��%s��@L ��4@���,ߐ!?�U�Jm�@��b~R�ٿ3�2&+X�@�sP4@
��Ʈ�!?F�R&���@>�Dh�ٿ{Ӝ��@�ts�[4@���Ŝ�!?{,���@�S�8S�ٿ-c�b<��@��ӧ(4@w��{��!?��G@�@�,!���ٿ�0�ly�@�+�o4@-2j(�!?�&����@�,!���ٿ�0�ly�@�+�o4@-2j(�!?�&����@�,!���ٿ�0�ly�@�+�o4@-2j(�!?�&����@�,!���ٿ�0�ly�@�+�o4@-2j(�!?�&����@�,!���ٿ�0�ly�@�+�o4@-2j(�!?�&����@��g�ٿ�:���@�=!!�4@^��Ր!?��?F�<�@��g�ٿ�:���@�=!!�4@^��Ր!?��?F�<�@��g�ٿ�:���@�=!!�4@^��Ր!?��?F�<�@��g�ٿ�:���@�=!!�4@^��Ր!?��?F�<�@��g�ٿ�:���@�=!!�4@^��Ր!?��?F�<�@��L�)�ٿ^��ّ�@���,�4@$���!?��>&�@��L�)�ٿ^��ّ�@���,�4@$���!?��>&�@��L�)�ٿ^��ّ�@���,�4@$���!?��>&�@��L�)�ٿ^��ّ�@���,�4@$���!?��>&�@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@�"*�ٿ��y���@�q�ќ4@��J�!?���f���@����ٿ���b���@�u>6�4@�DTА!?Ђެ���@����ٿ���b���@�u>6�4@�DTА!?Ђެ���@����ٿ���b���@�u>6�4@�DTА!?Ђެ���@����ٿ���b���@�u>6�4@�DTА!?Ђެ���@y��(��ٿ0�ҵ���@���NS4@\���ې!?�����@y��(��ٿ0�ҵ���@���NS4@\���ې!?�����@��"S��ٿo���''�@�w��q4@����֐!?�ILZc�@�N��ٿ>'S��@7�;S4@" �7Ԑ!?tFyI�@�N��ٿ>'S��@7�;S4@" �7Ԑ!?tFyI�@�N��ٿ>'S��@7�;S4@" �7Ԑ!?tFyI�@�N��ٿ>'S��@7�;S4@" �7Ԑ!?tFyI�@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@IU��D�ٿfp
_Zf�@'Xg�L4@�-�#�!?�ϓ�� �@�Y�a�ٿͷp8���@1��x�4@��֐!?&���@���^�ٿ=��O�h�@�n��4@�;{#ǐ!?mõ)ң�@���^�ٿ=��O�h�@�n��4@�;{#ǐ!?mõ)ң�@���^�ٿ=��O�h�@�n��4@�;{#ǐ!?mõ)ң�@���^�ٿ=��O�h�@�n��4@�;{#ǐ!?mõ)ң�@���^�ٿ=��O�h�@�n��4@�;{#ǐ!?mõ)ң�@�j�,��ٿu���@v4u�U4@�s�Ր!?j�Ф��@�j�,��ٿu���@v4u�U4@�s�Ր!?j�Ф��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@΅�>�ٿ�7�A��@~5�y�4@�y���!? �p�!��@��(��ٿ��*�7 �@�_��V4@@[��!?D�Kκ)�@��(��ٿ��*�7 �@�_��V4@@[��!?D�Kκ)�@c�F�0�ٿ�,	S1��@GS�b4@j�(P�!?�j�K�@c�F�0�ٿ�,	S1��@GS�b4@j�(P�!?�j�K�@c�F�0�ٿ�,	S1��@GS�b4@j�(P�!?�j�K�@c�F�0�ٿ�,	S1��@GS�b4@j�(P�!?�j�K�@c�F�0�ٿ�,	S1��@GS�b4@j�(P�!?�j�K�@.b�S�ٿ	-@d��@I�	/�4@���μ�!?鮪 �~�@.b�S�ٿ	-@d��@I�	/�4@���μ�!?鮪 �~�@.b�S�ٿ	-@d��@I�	/�4@���μ�!?鮪 �~�@t���>�ٿ_��$�@��qǀ4@�����!?֑�P���@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@F�%���ٿ�����@��/)�4@�{����!?��Af�~�@����o�ٿ֝+����@
V[4@�Bp�ܐ!?+�����@����o�ٿ֝+����@
V[4@�Bp�ܐ!?+�����@����o�ٿ֝+����@
V[4@�Bp�ܐ!?+�����@����o�ٿ֝+����@
V[4@�Bp�ܐ!?+�����@��U�ٿ"��7%�@�=!�.4@�R�I̐!?/�E \��@��U�ٿ"��7%�@�=!�.4@�R�I̐!?/�E \��@��U�ٿ"��7%�@�=!�.4@�R�I̐!?/�E \��@��U�ٿ"��7%�@�=!�.4@�R�I̐!?/�E \��@��U�ٿ"��7%�@�=!�.4@�R�I̐!?/�E \��@��ùֈٿ��BR�@���޸4@��2ΐ!?k�u��@��ùֈٿ��BR�@���޸4@��2ΐ!?k�u��@׺⣇ٿ���=�@|��084@D�'���!?�?�;J��@׺⣇ٿ���=�@|��084@D�'���!?�?�;J��@׺⣇ٿ���=�@|��084@D�'���!?�?�;J��@���	��ٿ������@\�G��4@���w��!?2I�����@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@�|��	�ٿ4�c'��@`r�+�4@<`���!??�S��V�@���+Ձٿ��ry���@��bj4@R���Ӑ!?w8��@�d��ٿhJ�(��@p��4@��8I�!?ć�A��@�d��ٿhJ�(��@p��4@��8I�!?ć�A��@!ս�ٿ]q'�E��@?S���4@D���B�!?�2���@�<��ٿ-����@%ub�$4@���]2�!?��]��@�<��ٿ-����@%ub�$4@���]2�!?��]��@ة㗷�ٿ�M��(��@U�˕��3@%6
2�!?�W�<U~�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@,B����ٿTj��(��@p��W4@3;m���!?�5��H�@SY���ٿ�Q��4�@PN��4@�1�ې!?���#�@SY���ٿ�Q��4�@PN��4@�1�ې!?���#�@SY���ٿ�Q��4�@PN��4@�1�ې!?���#�@SY���ٿ�Q��4�@PN��4@�1�ې!?���#�@SY���ٿ�Q��4�@PN��4@�1�ې!?���#�@���V4�ٿ�ۀ��@CY1��4@�!?Ua�M/�@���V4�ٿ�ۀ��@CY1��4@�!?Ua�M/�@�T��ٿL�����@�{��|4@�m��!?��[ ��@�d7W��ٿ#�Lf0{�@B��$��3@�0v�C�!?I,����@$E���ٿ���GR�@A�|�G4@U@c�!?�8����@$E���ٿ���GR�@A�|�G4@U@c�!?�8����@$E���ٿ���GR�@A�|�G4@U@c�!?�8����@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�UQ0�ٿY��R�@/y"[{4@ٌ�P�!?�y�*�A�@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�`a�K�ٿ3���8-�@d-�H74@u*jpn�!?�&�s���@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@�3o�X�ٿ��@R��@
h%W4@���ː!?�x��4��@��-���ٿpx�6��@�n5Á 4@�}����!?tL�O���@��-���ٿpx�6��@�n5Á 4@�}����!?tL�O���@��E�ٿ�z���@˯l_�4@v!(���!?�N����@��E�ٿ�z���@˯l_�4@v!(���!?�N����@��E�ٿ�z���@˯l_�4@v!(���!?�N����@�MyGщٿ3�C�#�@�թ�4@����!?�X���@�MyGщٿ3�C�#�@�թ�4@����!?�X���@�MyGщٿ3�C�#�@�թ�4@����!?�X���@�MyGщٿ3�C�#�@�թ�4@����!?�X���@�MyGщٿ3�C�#�@�թ�4@����!?�X���@�MyGщٿ3�C�#�@�թ�4@����!?�X���@������ٿPO;��@�ʉ�4@����!?
0����@o3���ٿk'����@7;G}�4@��o���!?��3�]3�@o3���ٿk'����@7;G}�4@��o���!?��3�]3�@o3���ٿk'����@7;G}�4@��o���!?��3�]3�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@]�i��ٿ��-����@cW�14@ϝ��)�!?��LZ�@ ��|C�ٿl8U�a��@��\�4@�[��!?*?q4���@ ��|C�ٿl8U�a��@��\�4@�[��!?*?q4���@ ��|C�ٿl8U�a��@��\�4@�[��!?*?q4���@An|�t�ٿ֙͑8'�@���#4@%���!?�8I���@An|�t�ٿ֙͑8'�@���#4@%���!?�8I���@ �Ob��ٿY��!�@q 5�H4@J��)��!?��I+}i�@�M~���ٿ�^/o���@[��4@�"���!?w���	E�@�M~���ٿ�^/o���@[��4@�"���!?w���	E�@1�E�n�ٿ���R
��@�]�t�4@خ� U�!?����X��@w��/�ٿ��9�W�@rI�q�4@i$�;Ґ!?���@w��/�ٿ��9�W�@rI�q�4@i$�;Ґ!?���@w��/�ٿ��9�W�@rI�q�4@i$�;Ґ!?���@ pZ�E�ٿ���L���@��.\�4@����Đ!?�^]���@ pZ�E�ٿ���L���@��.\�4@����Đ!?�^]���@68;�&�ٿ�M�}ҹ�@�P�4@�dB�L�!?���m��@68;�&�ٿ�M�}ҹ�@�P�4@�dB�L�!?���m��@68;�&�ٿ�M�}ҹ�@�P�4@�dB�L�!?���m��@68;�&�ٿ�M�}ҹ�@�P�4@�dB�L�!?���m��@��x��ٿs�� �F�@��p?4@��(da�!?�y���5�@��x��ٿs�� �F�@��p?4@��(da�!?�y���5�@
v��ǋٿc�;���@$�B4@�(i�[�!?�j�߶��@��&���ٿ�np��@A��)
4@�G��P�!?��K���@_7g�D�ٿ8�].�@P�}Dc4@A��؛�!?�y�SF��@_7g�D�ٿ8�].�@P�}Dc4@A��؛�!?�y�SF��@_7g�D�ٿ8�].�@P�}Dc4@A��؛�!?�y�SF��@_7g�D�ٿ8�].�@P�}Dc4@A��؛�!?�y�SF��@_7g�D�ٿ8�].�@P�}Dc4@A��؛�!?�y�SF��@66�!ٿ�� �)�@.��2�4@�ȝ�!?�h��>"�@}a�݄�ٿ50h���@�^7y�4@?����!?����O�@}a�݄�ٿ50h���@�^7y�4@?����!?����O�@��ᎋٿ�/��|�@�X6y�4@���n��!?A���7	�@��ᎋٿ�/��|�@�X6y�4@���n��!?A���7	�@��ᎋٿ�/��|�@�X6y�4@���n��!?A���7	�@��ᎋٿ�/��|�@�X6y�4@���n��!?A���7	�@��\:E�ٿ댛���@R�Dy�4@�2AT�!?p��.���@LΦ�|�ٿ������@�K�{	4@{�\��!?}�� D��@�A�Tyٿ�N����@/o��A4@�|�R1�!?�0lB�@�A�Tyٿ�N����@/o��A4@�|�R1�!?�0lB�@�p�Q��ٿ}�#W�@͂ܲ4@���V��!?�sS�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@�h�#~ٿ�Q�2��@�ֿT4@#p��Ґ!?�j��I�@��\׃ٿFD��@�&�f4@[o�Ӑ!?oF�<.�@��\׃ٿFD��@�&�f4@[o�Ӑ!?oF�<.�@��\׃ٿFD��@�&�f4@[o�Ӑ!?oF�<.�@��\׃ٿFD��@�&�f4@[o�Ӑ!?oF�<.�@H���܅ٿ��g�S�@Z-.�1	4@��b.��!?X�Njn��@W����ٿ8f�8�	�@�w��4@]�?i�!?���aY��@}O/��ٿ *�XЃ�@��4@]T��2�!?���w�@}O/��ٿ *�XЃ�@��4@]T��2�!?���w�@}O/��ٿ *�XЃ�@��4@]T��2�!?���w�@}O/��ٿ *�XЃ�@��4@]T��2�!?���w�@}O/��ٿ *�XЃ�@��4@]T��2�!?���w�@���Y�ٿ���&�s�@����4@��!?}�>�@���Y�ٿ���&�s�@����4@��!?}�>�@�6.�6�ٿ��nJ�l�@	�{"H4@��� ��!?��@ʂ��@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@<��>ԃٿ���)�[�@5m́4@������!?��,R���@P��n�ٿƝ�w���@���4@
`�\�!?�]�`(]�@P��n�ٿƝ�w���@���4@
`�\�!?�]�`(]�@�>BŅٿ��]��@�r��3@Tw�Ґ�!?	��;+s�@�>BŅٿ��]��@�r��3@Tw�Ґ�!?	��;+s�@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@����Ãٿ˗ja<�@�cY��4@ܧ�n�!?�{p��@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@��,�ٿ���vl�@{�E<C4@��Mg��!?�M�F�@Px�q�ٿE�QV�z�@�A#Y�4@	H�!?����@Px�q�ٿE�QV�z�@�A#Y�4@	H�!?����@Px�q�ٿE�QV�z�@�A#Y�4@	H�!?����@Px�q�ٿE�QV�z�@�A#Y�4@	H�!?����@�*!�2�ٿu�7,��@��;_4@G��9�!?ܺ�R�U�@�*!�2�ٿu�7,��@��;_4@G��9�!?ܺ�R�U�@�*!�2�ٿu�7,��@��;_4@G��9�!?ܺ�R�U�@�*!�2�ٿu�7,��@��;_4@G��9�!?ܺ�R�U�@�*!�2�ٿu�7,��@��;_4@G��9�!?ܺ�R�U�@��ok̃ٿ�\_Q8�@s�$4@�&"Ő!?%N�єJ�@��ok̃ٿ�\_Q8�@s�$4@�&"Ő!?%N�єJ�@��ok̃ٿ�\_Q8�@s�$4@�&"Ő!?%N�єJ�@��ok̃ٿ�\_Q8�@s�$4@�&"Ő!?%N�єJ�@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@�y[f<�ٿ�f}g���@sa���4@��Gܞ�!?�����@���vʅٿQ�lm���@�*#/4@`��!��!?]Kɟ��@���vʅٿQ�lm���@�*#/4@`��!��!?]Kɟ��@���vʅٿQ�lm���@�*#/4@`��!��!?]Kɟ��@���vʅٿQ�lm���@�*#/4@`��!��!?]Kɟ��@���vʅٿQ�lm���@�*#/4@`��!��!?]Kɟ��@A�P��ٿ��ff;��@?^:�;4@ys�Ȑ!?���3��@A�P��ٿ��ff;��@?^:�;4@ys�Ȑ!?���3��@A�P��ٿ��ff;��@?^:�;4@ys�Ȑ!?���3��@A�P��ٿ��ff;��@?^:�;4@ys�Ȑ!?���3��@�[0��ٿ"�L7N4�@�O0�4@!	�m�!?L�Grƶ�@�[0��ٿ"�L7N4�@�O0�4@!	�m�!?L�Grƶ�@�[0��ٿ"�L7N4�@�O0�4@!	�m�!?L�Grƶ�@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�Ns�ٿN<UA�K�@�6��4@�*!0��!?��t����@�����ٿ��QM2�@�}-�94@�>~cՐ!?�C��4	�@�����ٿ��QM2�@�}-�94@�>~cՐ!?�C��4	�@�����ٿ��QM2�@�}-�94@�>~cՐ!?�C��4	�@�&��R}ٿ'���@QS�4@H��ռ�!?��5��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@,�Eq�ٿ�@
T��@�7�j4@zس�!?��X�\��@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@���v�ٿ*�3V��@O���D4@P����!??q�����@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�J�;5�ٿ��4���@E�v�[4@�Ffx��!?%�qk�@�gA�ٿr����@���#4@hKː!?���+�@��{��~ٿO@��@�P�~4@ߒg{�!?�����@��{��~ٿO@��@�P�~4@ߒg{�!?�����@��{��~ٿO@��@�P�~4@ߒg{�!?�����@��{��~ٿO@��@�P�~4@ߒg{�!?�����@��{��~ٿO@��@�P�~4@ߒg{�!?�����@J z��ٿ�;3m8�@�5 4@��ٴ�!?/��,`�@J z��ٿ�;3m8�@�5 4@��ٴ�!?/��,`�@J z��ٿ�;3m8�@�5 4@��ٴ�!?/��,`�@J z��ٿ�;3m8�@�5 4@��ٴ�!?/��,`�@J z��ٿ�;3m8�@�5 4@��ٴ�!?/��,`�@�C���ٿ&����@���VV4@{�'�v�!?��G���@�C���ٿ&����@���VV4@{�'�v�!?��G���@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@�5aB�ٿ��K-���@���@4@��e���!?����_ �@S�@|�ٿ�#J@��@�y��" 4@��ِ!?�2�"��@S�@|�ٿ�#J@��@�y��" 4@��ِ!?�2�"��@S�@|�ٿ�#J@��@�y��" 4@��ِ!?�2�"��@S�@|�ٿ�#J@��@�y��" 4@��ِ!?�2�"��@�[]�=�ٿ���G9��@g�E4@�f��!?�j6Ӄ��@�[]�=�ٿ���G9��@g�E4@�f��!?�j6Ӄ��@�[]�=�ٿ���G9��@g�E4@�f��!?�j6Ӄ��@���8��ٿ�X4����@S����4@�%�`��!?w�REX�@���8��ٿ�X4����@S����4@�%�`��!?w�REX�@���8��ٿ�X4����@S����4@�%�`��!?w�REX�@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���^^�ٿ�ll2���@w��CU4@�PCpw�!?��1e}��@���6�ٿ�)m[�
�@�<���4@�O�zސ!?�W��2�@U�#���ٿi�Vd���@��Kj4@�#�J̐!?W:S@�2�@3�{�ٿ�rӴ-�@o/�׬4@�G�x��!?�p�k1��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@����A�ٿ"�:�=�@=�Li4@��r�j�!?�!n	��@Z�Z|ٿ����@��<4@���Q��!?(큂�@Z�Z|ٿ����@��<4@���Q��!?(큂�@+?#��ٿ�����@C��4@���!?�.����@,=��ٿ���W��@z�iv4@�#P���!?��8)���@,=��ٿ���W��@z�iv4@�#P���!?��8)���@,=��ٿ���W��@z�iv4@�#P���!?��8)���@,=��ٿ���W��@z�iv4@�#P���!?��8)���@,=��ٿ���W��@z�iv4@�#P���!?��8)���@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@��jt�ٿ��R)�@��S\�4@�XDd��!?���m'�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@����G�ٿX��}c�@�� ��4@�<��!?�u�o�@�W*m҅ٿ���w��@BF4@�0̌ΐ!?���n��@�W*m҅ٿ���w��@BF4@�0̌ΐ!?���n��@�W*m҅ٿ���w��@BF4@�0̌ΐ!?���n��@�W*m҅ٿ���w��@BF4@�0̌ΐ!?���n��@�W*m҅ٿ���w��@BF4@�0̌ΐ!?���n��@fo͈ٿ-U����@sf��4@ngz͐!?�M�1�h�@fo͈ٿ-U����@sf��4@ngz͐!?�M�1�h�@fo͈ٿ-U����@sf��4@ngz͐!?�M�1�h�@fo͈ٿ-U����@sf��4@ngz͐!?�M�1�h�@V-"��ٿ,!�bc�@��d�4@x.@���!?�պ��<�@V-"��ٿ,!�bc�@��d�4@x.@���!?�պ��<�@V-"��ٿ,!�bc�@��d�4@x.@���!?�պ��<�@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@��hʊٿ����@'K�g'4@��]���!?���m���@����B�ٿc���Q��@9O3�4@D,���!?e^�NmT�@��H���ٿ��7�I��@��:4@w%�h��!?�<�x�P�@k_N�j�ٿDK���@ͬ=�4@NU�m�!?�E�aLF�@k_N�j�ٿDK���@ͬ=�4@NU�m�!?�E�aLF�@k_N�j�ٿDK���@ͬ=�4@NU�m�!?�E�aLF�@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@�S��Äٿq�@��@��Y*�4@��x��!?��D֦��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@$q�嘇ٿ^��w�@'%Vް4@M$f���!?)|-��@0�8���ٿ�w����@���g�4@,�����!?��H��(�@0�8���ٿ�w����@���g�4@,�����!?��H��(�@�'LT��ٿlk����@f�Ye�4@�H���!?�Ǽ�w�@�'LT��ٿlk����@f�Ye�4@�H���!?�Ǽ�w�@�'LT��ٿlk����@f�Ye�4@�H���!?�Ǽ�w�@�'LT��ٿlk����@f�Ye�4@�H���!?�Ǽ�w�@K�	Ԁٿʪ<^�R�@�KT��4@����!?��U�8�@K�	Ԁٿʪ<^�R�@�KT��4@����!?��U�8�@K�	Ԁٿʪ<^�R�@�KT��4@����!?��U�8�@K�	Ԁٿʪ<^�R�@�KT��4@����!?��U�8�@6;0���ٿ��s��}�@ʋ��4@(R����!?�#�O��@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@����z�ٿ�t�r�a�@B���4@�y�+�!?S�����@G�!���ٿ7�/��u�@�h��4@Y���͐!?��^��@G�!���ٿ7�/��u�@�h��4@Y���͐!?��^��@G�!���ٿ7�/��u�@�h��4@Y���͐!?��^��@G�!���ٿ7�/��u�@�h��4@Y���͐!?��^��@GFf�ٿ�_*��@��o�4@�`8
��!?�M�A/��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@/�o��ٿ�m�����@����4@��u���!?��e��@��h)��ٿ,��5��@����4@0��
�!?j����v�@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@~��ٿc<�v�r�@zr�v~4@|ƭ��!?�5�n���@W�}f�ٿ	�)Z��@,�D�4@����*�!?!�wJ���@W�}f�ٿ	�)Z��@,�D�4@����*�!?!�wJ���@W�}f�ٿ	�)Z��@,�D�4@����*�!?!�wJ���@W�}f�ٿ	�)Z��@,�D�4@����*�!?!�wJ���@i�=�ۈٿݰ��!�@g'�4@ᙑp9�!?�6��_�@i�=�ۈٿݰ��!�@g'�4@ᙑp9�!?�6��_�@i�=�ۈٿݰ��!�@g'�4@ᙑp9�!?�6��_�@i�=�ۈٿݰ��!�@g'�4@ᙑp9�!?�6��_�@9S ~�ٿ�x�x���@ ���_4@�!ǐ!?�`�ŵ�@l1'{�ٿPHOW��@�V�4@%NgpĐ!?Z�N�xe�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@�-���ٿe>��׼�@b�ĭ4@0�)�!?��Q<�@U����~ٿ��8��@	sE�04@�a6B��!?��6�]�@U����~ٿ��8��@	sE�04@�a6B��!?��6�]�@t�[��~ٿ�ư�#�@a$���4@�,,��!?
�=�5�@t�[��~ٿ�ư�#�@a$���4@�,,��!?
�=�5�@t�[��~ٿ�ư�#�@a$���4@�,,��!?
�=�5�@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@PsꕀٿE�Ű���@p��`
4@�CH�!?+|��[��@Or�t��ٿr��c�q�@	��ީ4@�ʩdĐ!?�����@U�S}�ٿT�@�d�@E���	4@m1��!?��I�'F�@i�����ٿ*RU# +�@��N0I4@�MO`��!?j�$
�l�@i�����ٿ*RU# +�@��N0I4@�MO`��!?j�$
�l�@i�����ٿ*RU# +�@��N0I4@�MO`��!?j�$
�l�@S�E�
�ٿ�r�r���@]�͘k4@�pOG��!?��z~���@S�E�
�ٿ�r�r���@]�͘k4@�pOG��!?��z~���@�"[r�ٿ,���n�@X�d4@�Nb˻�!?�����-�@�"[r�ٿ,���n�@X�d4@�Nb˻�!?�����-�@�"[r�ٿ,���n�@X�d4@�Nb˻�!?�����-�@��व~ٿ�~�#��@;���U4@� ?�!?�rG��3�@��व~ٿ�~�#��@;���U4@� ?�!?�rG��3�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@y��,�ٿ
0�W�@P$�4@Pe7��!?F�u��1�@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@6�,�ٿ\��:�5�@"]Ƙ� 4@e�:�ѐ!?( �=\��@�ȮV�ٿ�2�,��@���4@�^c��!?a�6�w�@�ȮV�ٿ�2�,��@���4@�^c��!?a�6�w�@�ȮV�ٿ�2�,��@���4@�^c��!?a�6�w�@�ȮV�ٿ�2�,��@���4@�^c��!?a�6�w�@�ȮV�ٿ�2�,��@���4@�^c��!?a�6�w�@i%)��ٿ����G<�@�!�5s4@�����!?��W���@i%)��ٿ����G<�@�!�5s4@�����!?��W���@i%)��ٿ����G<�@�!�5s4@�����!?��W���@i%)��ٿ����G<�@�!�5s4@�����!?��W���@i%)��ٿ����G<�@�!�5s4@�����!?��W���@�Lǝ��ٿ=��6���@�"�4@���r�!?�R;&{�@�Lǝ��ٿ=��6���@�"�4@���r�!?�R;&{�@�Lǝ��ٿ=��6���@�"�4@���r�!?�R;&{�@E�/4�ٿQu�Ϻ�@C�-�=4@���P%�!?O���P�@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@𙴟�ٿ��W\�@�}l�;4@o?R2!?OBE���@�<�نٿ��Q?�p�@`���I4@���(��!?��q7���@�<�نٿ��Q?�p�@`���I4@���(��!?��q7���@�<�نٿ��Q?�p�@`���I4@���(��!?��q7���@�<�نٿ��Q?�p�@`���I4@���(��!?��q7���@����ٿ�?�I7��@�jy�E4@N�&��!?~�ԅK�@R�U��ٿ��[��@���8�4@U%�{�!?v�Vw?�@R�U��ٿ��[��@���8�4@U%�{�!?v�Vw?�@R�U��ٿ��[��@���8�4@U%�{�!?v�Vw?�@T1W�ٿu$�)��@�	��4@���x�!?�!�k^{�@T1W�ٿu$�)��@�	��4@���x�!?�!�k^{�@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@�xȆٿ����@��V��4@ S��ސ!?�"�H���@;��n�}ٿ��~ń)�@�а�4@�z`��!?��l=zl�@�27��ٿKJ���@%��yk4@[���w�!?��R����@�27��ٿKJ���@%��yk4@[���w�!?��R����@�27��ٿKJ���@%��yk4@[���w�!?��R����@�H�'��ٿ��m���@^��4@񒍋�!?���s؆�@�H�'��ٿ��m���@^��4@񒍋�!?���s؆�@��:�ٿԥ>]f�@)}�U!4@���}�!?�d�w|�@Pt�{�ٿO��u�@��M��4@@��!?D�@l�Y�@Pt�{�ٿO��u�@��M��4@@��!?D�@l�Y�@Pt�{�ٿO��u�@��M��4@@��!?D�@l�Y�@`7z͈ٿa�D����@R���4@�qA��!? ���ȓ�@G���ٿx&����@��_�c4@���K�!?�j��
�@G���ٿx&����@��_�c4@���K�!?�j��
�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�T�gǋٿ�{�;��@�d��4@*���!?� ��>�@�Y���ٿ��[��@[�C�4@���Ґ!?4���[v�@�Y���ٿ��[��@[�C�4@���Ґ!?4���[v�@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@��!��ٿ�8��a�@�i�N�4@>/S���!?爭`���@t��P-�ٿ7���7��@�$��4@��Y%�!?��x�7��@%�*��ٿYd���@NM�4@#�'jt�!?��d�%�@���8�ٿe�����@��X�	4@@✟�!?Uv'�V�@�y�>��ٿ����|��@��[~4@�]܍��!?��>6��@�y�>��ٿ����|��@��[~4@�]܍��!?��>6��@�y�>��ٿ����|��@��[~4@�]܍��!?��>6��@�y�>��ٿ����|��@��[~4@�]܍��!?��>6��@�$c�c�ٿ�ٷDn��@�n�6�4@�c�Ր!?V~d��;�@�$c�c�ٿ�ٷDn��@�n�6�4@�c�Ր!?V~d��;�@���a�ٿ�'����@S|W��4@-����!?V���.�@�O�'}�ٿ�;u�t�@ECu�4@�j�%��!?��x�u�@��{H�ٿ,�u51�@��JL4@~��p��!?�ũj�a�@��{H�ٿ,�u51�@��JL4@~��p��!?�ũj�a�@A�ß��ٿ*#��@�b#��4@a�b߲�!?ңS��@A�ß��ٿ*#��@�b#��4@a�b߲�!?ңS��@A�ß��ٿ*#��@�b#��4@a�b߲�!?ңS��@A�ß��ٿ*#��@�b#��4@a�b߲�!?ңS��@��Z#G�ٿ6����@/H�(W4@A���W�!?�a� x �@��Z#G�ٿ6����@/H�(W4@A���W�!?�a� x �@��Z#G�ٿ6����@/H�(W4@A���W�!?�a� x �@��7��ٿ#<����@�k][Q 4@��Q�Ð!?��T�H�@��7��ٿ#<����@�k][Q 4@��Q�Ð!?��T�H�@��7��ٿ#<����@�k][Q 4@��Q�Ð!?��T�H�@��7��ٿ#<����@�k][Q 4@��Q�Ð!?��T�H�@��7��ٿ#<����@�k][Q 4@��Q�Ð!?��T�H�@||l̊ٿ̏ R���@&�vms4@v��鮐!?z�-���@||l̊ٿ̏ R���@&�vms4@v��鮐!?z�-���@||l̊ٿ̏ R���@&�vms4@v��鮐!?z�-���@����ٿo�As���@��>�4@-+a���!?��;,�@����ٿo�As���@��>�4@-+a���!?��;,�@����ٿo�As���@��>�4@-+a���!?��;,�@����ٿo�As���@��>�4@-+a���!?��;,�@����ٿo�As���@��>�4@-+a���!?��;,�@�F�ٿ�o(};�@� ̬Y4@�&57��!?ԏ�����@KG<؂ٿ�G�� ��@:	�+�4@�~8b��!?VB����@Bt���ٿ�'�� ��@d��4@��f[9�!?�p����@Bt���ٿ�'�� ��@d��4@��f[9�!?�p����@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@c��݊ٿI'ԴG��@��4@b(U�6�!?Ā�3Y��@�|�x�ٿǄ]��:�@��u�>4@+c��!?��r^
��@�|�x�ٿǄ]��:�@��u�>4@+c��!?��r^
��@�|�x�ٿǄ]��:�@��u�>4@+c��!?��r^
��@<����ٿ�ӜՀ�@�%0�t4@�W��T�!?b���w�@<����ٿ�ӜՀ�@�%0�t4@�W��T�!?b���w�@<����ٿ�ӜՀ�@�%0�t4@�W��T�!?b���w�@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@��X"�ٿ~,��RV�@���)�4@�k���!?��,���@ k�x�ٿF���@��a�y4@CFTE	�!?So	�@(�$3�ٿ�a�����@�7ĉc4@�_��Z�!?ҔG�@(�$3�ٿ�a�����@�7ĉc4@�_��Z�!?ҔG�@(�$3�ٿ�a�����@�7ĉc4@�_��Z�!?ҔG�@���P��ٿŽ}��@���Q4@Up�l�!?�U��@���P��ٿŽ}��@���Q4@Up�l�!?�U��@͉'h��ٿ�z�7<��@���94@�ݴ&�!?���r�@�o�F�ٿ%��>��@����4@�%S��!?Ͼ�;���@�o�F�ٿ%��>��@����4@�%S��!?Ͼ�;���@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@���x�ٿJ������@��O=4@i�2��!?��W*�@+�1�ٿ�P�
P�@���Fs4@ȟR�V�!?/�Զ~f�@+�1�ٿ�P�
P�@���Fs4@ȟR�V�!?/�Զ~f�@_l�U��ٿ�e���
�@�y�'�4@Y�� ��!?�\�X"�@_l�U��ٿ�e���
�@�y�'�4@Y�� ��!?�\�X"�@��;όٿ�G�6��@?fҺ4@k�ti�!?�e@��`�@>Ϊh>�ٿwӓs��@�t> �4@���(ɐ!?GA���@>Ϊh>�ٿwӓs��@�t> �4@���(ɐ!?GA���@>Ϊh>�ٿwӓs��@�t> �4@���(ɐ!?GA���@>Ϊh>�ٿwӓs��@�t> �4@���(ɐ!?GA���@S���ٿ*؇����@��1��4@L1��!?#z�)���@S���ٿ*؇����@��1��4@L1��!?#z�)���@S���ٿ*؇����@��1��4@L1��!?#z�)���@fj�m|�ٿO��mȹ�@#D�		4@���e�!?�	H1��@�C9�j�ٿb�!���@�����4@(�y	�!?�-݂0G�@�C9�j�ٿb�!���@�����4@(�y	�!?�-݂0G�@�C9�j�ٿb�!���@�����4@(�y	�!?�-݂0G�@�� *�ٿSe��+�@)s
^	4@}���ڐ!?�2z���@%WaO�ٿl�/ٔ��@�Z�?4@�M���!?sQ'>��@�𬺪�ٿ�v��@�t�*�4@O�胐!?C���Ϳ�@�𬺪�ٿ�v��@�t�*�4@O�胐!?C���Ϳ�@�𬺪�ٿ�v��@�t�*�4@O�胐!?C���Ϳ�@�𬺪�ٿ�v��@�t�*�4@O�胐!?C���Ϳ�@�\_��ٿm�"���@ȟ��4@P3�ri�!?8�`����@�\_��ٿm�"���@ȟ��4@P3�ri�!?8�`����@�\_��ٿm�"���@ȟ��4@P3�ri�!?8�`����@�\_��ٿm�"���@ȟ��4@P3�ri�!?8�`����@�\_��ٿm�"���@ȟ��4@P3�ri�!?8�`����@�E���ٿ�֞(���@᷻�/4@��x#I�!?RZ��_��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@$7��D�ٿ�w��3�@S��c4@�D�Qr�!?�:�ۋ��@�|��ٿb���z�@�39��4@������!?��C�l��@�|��ٿb���z�@�39��4@������!?��C�l��@����ٿ��wC�*�@� ��4@0�Ґ!?������@T��I�ٿ��9�2�@�I�` 4@�<M6�!?���C��@T��I�ٿ��9�2�@�I�` 4@�<M6�!?���C��@�h|ٿ�^N��@��t�4@����!?[�q�W�@�h|ٿ�^N��@��t�4@����!?[�q�W�@f4t���ٿ��$��p�@L���D	4@�R$��!?(��G���@f4t���ٿ��$��p�@L���D	4@�R$��!?(��G���@b;._��ٿ��9�@Xq�n4@\Qb�!?�S0���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�)�i̓ٿ�"�_Z�@��pp�4@�b{���!?�H���@�;b�{�ٿ%����@q�P4@g�����!?��.4��@�;b�{�ٿ%����@q�P4@g�����!?��.4��@���9�ٿ8��-�"�@�l2>4@6-�ؒ�!?���.BY�@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@;�r؇ٿ%�s���@^�c<q4@�Euxb�!?�Yr���@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@���c�ٿ���h�@S4w4@wZb��!?�r��_�@ڹ!���ٿBY, gf�@v��74@���"��!?����|�@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@_����ٿ	��yk��@	_>�@4@�ᴗ��!?�<��@�ވ���ٿZ]�ϴ�@6Ζ�4@��M@א!?iy���7�@�ވ���ٿZ]�ϴ�@6Ζ�4@��M@א!?iy���7�@�ވ���ٿZ]�ϴ�@6Ζ�4@��M@א!?iy���7�@�ވ���ٿZ]�ϴ�@6Ζ�4@��M@א!?iy���7�@�d�k�ٿ���
��@p��@4@4%���!?keu���@�d�k�ٿ���
��@p��@4@4%���!?keu���@�d�k�ٿ���
��@p��@4@4%���!?keu���@�QY}�ٿ�F��oF�@��x��4@��W4�!?'=,�d��@�QY}�ٿ�F��oF�@��x��4@��W4�!?'=,�d��@�QY}�ٿ�F��oF�@��x��4@��W4�!?'=,�d��@�'��ٿ���"%J�@���X�4@�.�q��!?yߦk�@�Ш �ٿ�8��/G�@Uߎ]d4@\6�!?\o>Y��@�Ш �ٿ�8��/G�@Uߎ]d4@\6�!?\o>Y��@Q��Bۆٿ2 �Ʒ�@a�1	4@�~`Y��!?=�|*���@Q��Bۆٿ2 �Ʒ�@a�1	4@�~`Y��!?=�|*���@Q��Bۆٿ2 �Ʒ�@a�1	4@�~`Y��!?=�|*���@Q��Bۆٿ2 �Ʒ�@a�1	4@�~`Y��!?=�|*���@Q��Bۆٿ2 �Ʒ�@a�1	4@�~`Y��!?=�|*���@A��'N�ٿ���?�@o8O�"4@��MF��!?�GCq�Z�@A��'N�ٿ���?�@o8O�"4@��MF��!?�GCq�Z�@�Q&e�ٿ���aM�@�wS�4@��-5��!?��t4�J�@�Q&e�ٿ���aM�@�wS�4@��-5��!?��t4�J�@�Q&e�ٿ���aM�@�wS�4@��-5��!?��t4�J�@�Q&e�ٿ���aM�@�wS�4@��-5��!?��t4�J�@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@ɸ�g�{ٿ���!:��@t??ֵ4@$�B饐!?�˕����@��ٿ1M��I�@=�r�/�3@��Yu��!?�b^N�	�@��ٿ1M��I�@=�r�/�3@��Yu��!?�b^N�	�@ܒ�ٿ�2/�b��@�ގ
N 4@)�;��!?�Tr���@���@ʁٿf�(�>��@��勃4@I!�j��!?�g[����@���@ʁٿf�(�>��@��勃4@I!�j��!?�g[����@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��G�/�ٿﾚB���@̙Z�4@*�N�$�!?�I�j��@��&�}ٿ�o�虌�@|��a4@`J��א!?�D�ܠ��@��&�}ٿ�o�虌�@|��a4@`J��א!?�D�ܠ��@��&�}ٿ�o�虌�@|��a4@`J��א!?�D�ܠ��@;Y�r�ٿ	P&ia��@y��E�4@��(
�!?� cF��@;Y�r�ٿ	P&ia��@y��E�4@��(
�!?� cF��@�Y��/�ٿʪ�M��@ʉ��4@�@�:1�!?�ײ�y�@�Y��/�ٿʪ�M��@ʉ��4@�@�:1�!?�ײ�y�@�Y��/�ٿʪ�M��@ʉ��4@�@�:1�!?�ײ�y�@�Y��/�ٿʪ�M��@ʉ��4@�@�:1�!?�ײ�y�@���ځٿB�.���@,��k4@�W�'ǐ!?�u���@���ځٿB�.���@,��k4@�W�'ǐ!?�u���@Ts����ٿS3�,��@mpcl04@6b��̐!?��u����@Ts����ٿS3�,��@mpcl04@6b��̐!?��u����@Ts����ٿS3�,��@mpcl04@6b��̐!?��u����@Ts����ٿS3�,��@mpcl04@6b��̐!?��u����@VS��ٿ���|�@�*��4@a�CRɐ!?�:���@VS��ٿ���|�@�*��4@a�CRɐ!?�:���@VS��ٿ���|�@�*��4@a�CRɐ!?�:���@VS��ٿ���|�@�*��4@a�CRɐ!?�:���@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�V��=�ٿ��&�t�@��qp4@q#޾�!?;��:�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@�z��u�ٿ�Z�C���@]��4@�|TӐ!?��J�@4��T~�ٿҔ:H�2�@�ܺF4@�ZV4�!?� ,���@4��T~�ٿҔ:H�2�@�ܺF4@�ZV4�!?� ,���@4��T~�ٿҔ:H�2�@�ܺF4@�ZV4�!?� ,���@�5��Ǐٿ:W-����@�@��4@�m��H�!?68��w@�@�5��Ǐٿ:W-����@�@��4@�m��H�!?68��w@�@��{/�ٿiJ����@׬J�4@����$�!?1��@���@��{/�ٿiJ����@׬J�4@����$�!?1��@���@��{/�ٿiJ����@׬J�4@����$�!?1��@���@��{/�ٿiJ����@׬J�4@����$�!?1��@���@��{/�ٿiJ����@׬J�4@����$�!?1��@���@��{/�ٿiJ����@׬J�4@����$�!?1��@���@���ٿ�3��@/xM�4@VH���!?B��K��@��֓�|ٿ���@FX�U'4@����|�!?��A(c�@�¢$�ٿ&�[k*�@�1�	!4@�f;��!?v!��p�@�¢$�ٿ&�[k*�@�1�	!4@�f;��!?v!��p�@�"��އٿ�kp��]�@j���H4@\r�}o�!?ƽ����@�"��އٿ�kp��]�@j���H4@\r�}o�!?ƽ����@�"��އٿ�kp��]�@j���H4@\r�}o�!?ƽ����@�"��އٿ�kp��]�@j���H4@\r�}o�!?ƽ����@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@���S��ٿԐd����@f/tG>4@h����!?Gb	�m�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@� �1)�ٿ��=N��@�W�F4@��{ѐ!?0�,`h�@����ٿ7���&�@`�̶��3@D�Ϙ��!?�&F5���@����ٿ7���&�@`�̶��3@D�Ϙ��!?�&F5���@����ٿ7���&�@`�̶��3@D�Ϙ��!?�&F5���@1t4Z�ٿ�LǛ�@iCLJ�3@v\s��!?�]��2�@1�{ΐ�ٿ'$��@�)y�n 4@�?-��!?��㔑��@1�{ΐ�ٿ'$��@�)y�n 4@�?-��!?��㔑��@W�)�W�ٿ�#=/�@ַ�n4@�hg�!?����|�@W�)�W�ٿ�#=/�@ַ�n4@�hg�!?����|�@����ٿ��70N��@��u�m4@����!?q��Hm��@����ٿ��70N��@��u�m4@����!?q��Hm��@����ٿ��70N��@��u�m4@����!?q��Hm��@����ٿ��70N��@��u�m4@����!?q��Hm��@����ٿ��70N��@��u�m4@����!?q��Hm��@����ٿ��70N��@��u�m4@����!?q��Hm��@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@Q�����ٿ�%_��@�@�u��4@�d"�c�!?$ٟ�G�@�	T�'�ٿ����C��@�J��4@���M�!?���4��@�	T�'�ٿ����C��@�J��4@���M�!?���4��@�	T�'�ٿ����C��@�J��4@���M�!?���4��@�	T�'�ٿ����C��@�J��4@���M�!?���4��@�	T�'�ٿ����C��@�J��4@���M�!?���4��@��Q6�ٿz��ԏ�@~g�4@�ʆü�!?�8l��@��Q6�ٿz��ԏ�@~g�4@�ʆü�!?�8l��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@bT�6|ٿ����1s�@D�0��4@3�r��!?-�֙��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@�L�Z�ٿ��T)B�@�j�ӣ4@�5��!?d��Xg��@���@�ٿ����@̾��4@{��Z�!?P!�c[��@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@���ˁٿ�W	���@gG�64@g%^�!?��\����@��:ٿ
�-��@E	s�4@����Q�!?�a� @�@��:ٿ
�-��@E	s�4@����Q�!?�a� @�@��:ٿ
�-��@E	s�4@����Q�!?�a� @�@��:ٿ
�-��@E	s�4@����Q�!?�a� @�@�:6m�ٿ�^�C���@��T�t4@W2�|g�!?;�	�T\�@�:6m�ٿ�^�C���@��T�t4@W2�|g�!?;�	�T\�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@?C��zٿ:����@t���	4@'�J��!?�^�ZV/�@`8Ⱦzٿ'���?�@#��.4@��;z�!?O�JD�@`8Ⱦzٿ'���?�@#��.4@��;z�!?O�JD�@`8Ⱦzٿ'���?�@#��.4@��;z�!?O�JD�@����ٿ��ߏ?3�@�n<I�4@��E�!?�R��M��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@Y�>�ٿ ,����@]u�:�4@t����!?�%X[��@zQL�0�ٿ
B��'}�@5v["
4@;p)��!?�KD����@zQL�0�ٿ
B��'}�@5v["
4@;p)��!?�KD����@zQL�0�ٿ
B��'}�@5v["
4@;p)��!?�KD����@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@"$[�ٿ?$��Z��@4+���4@�� )t�!?{,�G��@�9�t�ٿ.Įm���@�֏w4@{�n���!?&���G�@7�Nƙ�ٿ�L�^��@�/6RC4@6$?|	�!?�1A0y�@7�Nƙ�ٿ�L�^��@�/6RC4@6$?|	�!?�1A0y�@7�Nƙ�ٿ�L�^��@�/6RC4@6$?|	�!?�1A0y�@7�Nƙ�ٿ�L�^��@�/6RC4@6$?|	�!?�1A0y�@{Ќ��ٿTY@�`e�@��H4@/�]"ΐ!?Fc˅���@�$��ٿ"j�g��@��ґ4@O��I�!?~j)K���@�$��ٿ"j�g��@��ґ4@O��I�!?~j)K���@f�R:��ٿl*�n��@�]��_4@�S�#ؐ!?�.��P��@f�R:��ٿl*�n��@�]��_4@�S�#ؐ!?�.��P��@f�R:��ٿl*�n��@�]��_4@�S�#ؐ!?�.��P��@��d�a�ٿOo�����@�+_9�3@?n>א!?o��@���@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Y_�$�ٿ{�����@0t���4@��h���!?[�.3�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�Z�n�ٿT�3���@����4@�Bm���!?����q-�@�95[��ٿoam����@O�R.4@{�i���!?����ǖ�@��T���ٿc�ʭK�@�E� 4@G9=}ې!?=�|���@��T���ٿc�ʭK�@�E� 4@G9=}ې!?=�|���@�x�p)�ٿ �.΀��@ ��4�3@%�C2��!?��zT��@�x�p)�ٿ �.΀��@ ��4�3@%�C2��!?��zT��@�x�p)�ٿ �.΀��@ ��4�3@%�C2��!?��zT��@	�U���ٿ�ҘU��@D0�4@>�D��!?�MF�%f�@	�U���ٿ�ҘU��@D0�4@>�D��!?�MF�%f�@����ٿ�����@�6��4@_۬��!?=X���(�@����ǅٿ+��}���@yLD��4@u3|��!?��{�~�@����ǅٿ+��}���@yLD��4@u3|��!?��{�~�@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@n��.u�ٿ/Q�@�(�M�4@������!?j�\_��@x?�
��ٿ}YG&'��@:�� e4@[-ƈ�!?��XH��@x?�
��ٿ}YG&'��@:�� e4@[-ƈ�!?��XH��@K�CK�ٿ@�-�9�@�a��4@iIOzϐ!?�_�i�m�@�}���ٿ` Z<���@�A�ۚ	4@�]�ڐ!?��QE�y�@�}���ٿ` Z<���@�A�ۚ	4@�]�ڐ!?��QE�y�@&��{��ٿ�"�WPh�@>N�. 4@ bS���!?p_�?0�@&��{��ٿ�"�WPh�@>N�. 4@ bS���!?p_�?0�@&��{��ٿ�"�WPh�@>N�. 4@ bS���!?p_�?0�@&��{��ٿ�"�WPh�@>N�. 4@ bS���!?p_�?0�@&��{��ٿ�"�WPh�@>N�. 4@ bS���!?p_�?0�@�ߺ0�ٿ5�Ֆ���@XZ�4@�*=��!?�u�[���@�ߺ0�ٿ5�Ֆ���@XZ�4@�*=��!?�u�[���@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@4G^hM�ٿ����t�@�UO4@m�>���!?P�/e`!�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@l0,ߊٿG��n��@�;�W�4@fX���!?��t�.=�@.Ӷ���ٿ�B÷b�@?��#4@�kf���!?��8���@.Ӷ���ٿ�B÷b�@?��#4@�kf���!?��8���@.Ӷ���ٿ�B÷b�@?��#4@�kf���!?��8���@H��"��ٿm6�錋�@fw��t4@��̐!?s�._��@H��"��ٿm6�錋�@fw��t4@��̐!?s�._��@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@U^�Y��ٿ� ?;x��@2��g�4@��-�ߐ!?�0���@�5���ٿ|�&h@8�@�Q"l�4@ H��ǐ!?�\����@�5���ٿ|�&h@8�@�Q"l�4@ H��ǐ!?�\����@�5���ٿ|�&h@8�@�Q"l�4@ H��ǐ!?�\����@���XQ~ٿ�=��@E�[L	4@��;��!?�0����@���XQ~ٿ�=��@E�[L	4@��;��!?�0����@���XQ~ٿ�=��@E�[L	4@��;��!?�0����@���XQ~ٿ�=��@E�[L	4@��;��!?�0����@���XQ~ٿ�=��@E�[L	4@��;��!?�0����@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@E�w�-�ٿK~<�@��J�4@7���!?R�Z3:p�@�}ӨK}ٿw�*%���@�����4@UZ��!?��]¹<�@�<���}ٿ��2�@殨*34@4����!?�s����@�<���}ٿ��2�@殨*34@4����!?�s����@�<���}ٿ��2�@殨*34@4����!?�s����@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@W]��}ٿ�QMv5��@�T!�4@��m�~�!?��6b>C�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@N�O��ٿ苘j�@�#y�4@R tQr�!?L��@�@_)D��ٿ�����Y�@Uk�4@2S*C�!?�%f����@_)D��ٿ�����Y�@Uk�4@2S*C�!?�%f����@_)D��ٿ�����Y�@Uk�4@2S*C�!?�%f����@_>���ٿrPa���@�[�4@2�1�!?µ6�i�@>V��"�ٿ����w�@�q��4@Waշ��!?�B�czj�@>V��"�ٿ����w�@�q��4@Waշ��!?�B�czj�@>V��"�ٿ����w�@�q��4@Waշ��!?�B�czj�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@kS,���ٿ�A�v �@ihPRH4@1����!?Z��X1�@�(c���ٿ�#����@İ��4@ �k�Ր!?�ag��i�@]rr*H�ٿ�/��4�@�u�4@�w�Đ!?�HcHc��@'�$�C�ٿ�?Uܗ'�@��U�e4@;je�!?���`]�@���ٿ���B��@�@��}4@ă�#r�!?۫�� �@���ٿ���B��@�@��}4@ă�#r�!?۫�� �@���ٿ���B��@�@��}4@ă�#r�!?۫�� �@&�C�A�ٿ���@�P���4@iTO��!?�˲�8�@&�C�A�ٿ���@�P���4@iTO��!?�˲�8�@&�C�A�ٿ���@�P���4@iTO��!?�˲�8�@&�C�A�ٿ���@�P���4@iTO��!?�˲�8�@&�C�A�ٿ���@�P���4@iTO��!?�˲�8�@����Ջٿ�ja�%k�@&�(� 4@��%!?�s�1��@����Ջٿ�ja�%k�@&�(� 4@��%!?�s�1��@����Ջٿ�ja�%k�@&�(� 4@��%!?�s�1��@����Ջٿ�ja�%k�@&�(� 4@��%!?�s�1��@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@$xG(�ٿV8P���@�^� "4@U�:��!?G���a�@����ٿ��&�e�@�K��'4@
=P��!?S��k��@����ٿ��&�e�@�K��'4@
=P��!?S��k��@����ٿ��&�e�@�K��'4@
=P��!?S��k��@�2��/�ٿ������@j�Ȏ�4@K��F�!?���6���@�2��/�ٿ������@j�Ȏ�4@K��F�!?���6���@�2��/�ٿ������@j�Ȏ�4@K��F�!?���6���@�p,*��ٿ|��]��@PN��4@���_�!?ҳ���@�p,*��ٿ|��]��@PN��4@���_�!?ҳ���@9����ٿO����3�@�ҽ��4@���*�!?ySN���@9����ٿO����3�@�ҽ��4@���*�!?ySN���@9����ٿO����3�@�ҽ��4@���*�!?ySN���@9����ٿO����3�@�ҽ��4@���*�!?ySN���@�@N���ٿ��� �E�@-����4@P�X1�!?����'��@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@~"v���ٿ i�=�@C�о 4@}��!z�!?�2�%�{�@Sd�)�ٿ%������@6�{� 4@k�i�ؐ!?�aC�V��@Sd�)�ٿ%������@6�{� 4@k�i�ؐ!?�aC�V��@Sd�)�ٿ%������@6�{� 4@k�i�ؐ!?�aC�V��@Sd�)�ٿ%������@6�{� 4@k�i�ؐ!?�aC�V��@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@��d���ٿ'؆ ��@Yd�[�4@�˲�ǐ!?�����@���g��ٿ��ǔ,d�@���(4@����!?�OD��P�@���g��ٿ��ǔ,d�@���(4@����!?�OD��P�@���g��ٿ��ǔ,d�@���(4@����!?�OD��P�@ !��ٿ��.�Y��@�$P�4@���9s�!?��>�R�@ !��ٿ��.�Y��@�$P�4@���9s�!?��>�R�@ !��ٿ��.�Y��@�$P�4@���9s�!?��>�R�@ !��ٿ��.�Y��@�$P�4@���9s�!?��>�R�@��{���ٿ�
G�@��@Hp\�4@{Qg�!?��r��@��{���ٿ�
G�@��@Hp\�4@{Qg�!?��r��@��{���ٿ�
G�@��@Hp\�4@{Qg�!?��r��@o�`��ٿȌ �[��@j�9��4@�C����!?fwn����@o�`��ٿȌ �[��@j�9��4@�C����!?fwn����@o�`��ٿȌ �[��@j�9��4@�C����!?fwn����@o�`��ٿȌ �[��@j�9��4@�C����!?fwn����@���&ٿ6�HЧ�@��E��4@T��ʓ�!?��O|N�@K��V�ٿ{��c��@x��t4@̹�!?=�D�w�@S�Qo��ٿ��͐��@��J�4@h�Y�Ր!?fn��&��@S�Qo��ٿ��͐��@��J�4@h�Y�Ր!?fn��&��@S�Qo��ٿ��͐��@��J�4@h�Y�Ր!?fn��&��@S�Qo��ٿ��͐��@��J�4@h�Y�Ր!?fn��&��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@��*�ٿ�P9[ �@���Zz4@���#��!?'�m|��@%�ٿ.� ���@p�3�4@}�7��!?��>��@%�ٿ.� ���@p�3�4@}�7��!?��>��@<=I[�ٿ�d���@$�uK4@&Ȼ��!?��ژi�@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��r�!�ٿ�S�W���@���H4@]��*��!?��R���@��z�ٿ�u�y��@v�|h4@;��?�!?��t���@��z�ٿ�u�y��@v�|h4@;��?�!?��t���@��z�ٿ�u�y��@v�|h4@;��?�!?��t���@�D&��ٿ�ci���@_�1\�4@�?����!?� ��h�@�g����ٿ1t��DW�@��N�P4@�搶�!? w�tp�@�g����ٿ1t��DW�@��N�P4@�搶�!? w�tp�@�g����ٿ1t��DW�@��N�P4@�搶�!? w�tp�@�g����ٿ1t��DW�@��N�P4@�搶�!? w�tp�@�+�t�ٿ����!��@�L?4@_&R���!?�V�# �@����ٿ?ϵ�N��@b�U��4@Y�"�'�!?�Cx���@�{�p�}ٿ�>����@"�и�4@ԍ�=�!?m���>�@�{�p�}ٿ�>����@"�и�4@ԍ�=�!?m���>�@k�����ٿX���S��@�	j��4@iߗ��!?1C��!�@k�����ٿX���S��@�	j��4@iߗ��!?1C��!�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�e�";�ٿM@!�/��@���T�4@ʜ:��!?(�]�Hc�@�.o���ٿ�*���@=�c�e4@�Zyk�!?Qo=�9�@�.o���ٿ�*���@=�c�e4@�Zyk�!?Qo=�9�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@^m���ٿ��mF��@qp��4@��(��!?���@�k�@��hďٿ��&���@Ex1� 4@
Y�Ȑ!?��٠��@��hďٿ��&���@Ex1� 4@
Y�Ȑ!?��٠��@��hďٿ��&���@Ex1� 4@
Y�Ȑ!?��٠��@��hďٿ��&���@Ex1� 4@
Y�Ȑ!?��٠��@��JP�ٿ5E��� �@@��"64@��y���!?��@�Bn�@��JP�ٿ5E��� �@@��"64@��y���!?��@�Bn�@��JP�ٿ5E��� �@@��"64@��y���!?��@�Bn�@X
z&>�ٿ-N}���@s$�4@��_А!?��N��r�@N;���ٿ}nh��e�@�X�4@�|��֐!?_�y�hZ�@N;���ٿ}nh��e�@�X�4@�|��֐!?_�y�hZ�@N;���ٿ}nh��e�@�X�4@�|��֐!?_�y�hZ�@N;���ٿ}nh��e�@�X�4@�|��֐!?_�y�hZ�@N;���ٿ}nh��e�@�X�4@�|��֐!?_�y�hZ�@H:��ٿ��2��@�^��v4@Y��f+�!?V�eA���@H:��ٿ��2��@�^��v4@Y��f+�!?V�eA���@zו��ٿ�O��?��@b�pd� 4@{�̐!?���`a�@zו��ٿ�O��?��@b�pd� 4@{�̐!?���`a�@zו��ٿ�O��?��@b�pd� 4@{�̐!?���`a�@��♌ٿ��i9(�@p���� 4@�%6g��!?�E:���@��♌ٿ��i9(�@p���� 4@�%6g��!?�E:���@��♌ٿ��i9(�@p���� 4@�%6g��!?�E:���@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@2S��ٿ"H}4c�@���-�4@��bD�!?���;�@�i���ٿI�U=�@j,��4@��@��!?��?W��@\��kޅٿӱ�݅�@j�U��4@E�`�!?_������@\��kޅٿӱ�݅�@j�U��4@E�`�!?_������@\��kޅٿӱ�݅�@j�U��4@E�`�!?_������@\��kޅٿӱ�݅�@j�U��4@E�`�!?_������@��}�ۈٿv�c�/�@��	�;4@g�֜5�!?������@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@�r�[��ٿ����g�@���V4@d�L�!?QJA���@GI�D�ٿ��Z*{�@�^	�H4@�N��!?Ue/"s��@GI�D�ٿ��Z*{�@�^	�H4@�N��!?Ue/"s��@GI�D�ٿ��Z*{�@�^	�H4@�N��!?Ue/"s��@*~ʐȒٿ��`�E�@��W�4@���ې!?{�Ea[��@�g��ϔٿ4ܗ@/(�@G-d�s4@b;gb�!?�h�6��@�g��ϔٿ4ܗ@/(�@G-d�s4@b;gb�!?�h�6��@�g��ϔٿ4ܗ@/(�@G-d�s4@b;gb�!?�h�6��@�g��ϔٿ4ܗ@/(�@G-d�s4@b;gb�!?�h�6��@�Ф��ٿ�����k�@-�^a�4@�>�!?.�K�[�@�Ф��ٿ�����k�@-�^a�4@�>�!?.�K�[�@K	�-ـٿn����@��4@� BQ�!?�j����@K	�-ـٿn����@��4@� BQ�!?�j����@��V�~ٿ�� (�@����0 4@���~�!?�,��<�@��V�~ٿ�� (�@����0 4@���~�!?�,��<�@��V�~ٿ�� (�@����0 4@���~�!?�,��<�@��V�~ٿ�� (�@����0 4@���~�!?�,��<�@͵�G��ٿx���1o�@�>Cl4@#1H��!?��'@	:�@͵�G��ٿx���1o�@�>Cl4@#1H��!?��'@	:�@͵�G��ٿx���1o�@�>Cl4@#1H��!?��'@	:�@͵�G��ٿx���1o�@�>Cl4@#1H��!?��'@	:�@͵�G��ٿx���1o�@�>Cl4@#1H��!?��'@	:�@G	bh�ٿ)sq����@k�+��4@q#� }�!?�e����@G	bh�ٿ)sq����@k�+��4@q#� }�!?�e����@G	bh�ٿ)sq����@k�+��4@q#� }�!?�e����@G	bh�ٿ)sq����@k�+��4@q#� }�!?�e����@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@mk�O�ٿR^���@�O�|4@�E�U��!?��8ҩ�@}�܀C�ٿ��J���@d"B4@�>�X��!?���W�9�@}�܀C�ٿ��J���@d"B4@�>�X��!?���W�9�@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��z0��ٿ��|��^�@���4@)�����!?��aY��@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@��g♋ٿ��%'+�@f�ApM4@D���m�!?4��%���@�"���ٿ�u���@��<ψ4@�51w�!?�P�b�@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@�V,V�ٿN�?��@�"Z8�4@�9��b�!?^�����@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@Z�� ��ٿ�Ā�?��@�D��w4@���4��!?�Г�S�@{���ٿO_�ThC�@�.@��4@��l��!?�b)��@{���ٿO_�ThC�@�.@��4@��l��!?�b)��@{���ٿO_�ThC�@�.@��4@��l��!?�b)��@(��^�ٿ��X���@�Ŏ��4@�m�֐!?�x�
4��@��5��ٿ~��=��@<��4@��=�Ő!?�St���@��'��ٿp�kT���@̾���4@� ɢ�!?� ����@��'��ٿp�kT���@̾���4@� ɢ�!?� ����@��'��ٿp�kT���@̾���4@� ɢ�!?� ����@��'��ٿp�kT���@̾���4@� ɢ�!?� ����@��'��ٿp�kT���@̾���4@� ɢ�!?� ����@xh��ٿ|�u��u�@\��b4@��ԣ�!?������@xh��ٿ|�u��u�@\��b4@��ԣ�!?������@o����ٿL��th��@�o��j 4@���͐!?�*9YM�@o����ٿL��th��@�o��j 4@���͐!?�*9YM�@o����ٿL��th��@�o��j 4@���͐!?�*9YM�@o����ٿL��th��@�o��j 4@���͐!?�*9YM�@o����ٿL��th��@�o��j 4@���͐!?�*9YM�@0\�]��ٿ�_G.؊�@�!��4@�oh��!?��x	\�@0\�]��ٿ�_G.؊�@�!��4@�oh��!?��x	\�@x���ٿ����p��@�$��j4@�/�r�!?��6l�C�@x���ٿ����p��@�$��j4@�/�r�!?��6l�C�@��;h�ٿ%9�D�5�@)E�P4@�Y)p�!?���&�@��;h�ٿ%9�D�5�@)E�P4@�Y)p�!?���&�@��;h�ٿ%9�D�5�@)E�P4@�Y)p�!?���&�@��Ԕp�ٿ�HH�I�@��y~�4@H�&���!?�������@��Ԕp�ٿ�HH�I�@��y~�4@H�&���!?�������@���كٿ#� P�@+���,4@�
�F��!?Ӏ`�{��@���كٿ#� P�@+���,4@�
�F��!?Ӏ`�{��@���كٿ#� P�@+���,4@�
�F��!?Ӏ`�{��@��وٿ���p��@���4@����Ԑ!? �O���@��وٿ���p��@���4@����Ԑ!? �O���@D�!�ٿ�s�Q��@:���4@�|E7��!?�c9{N8�@D�!�ٿ�s�Q��@:���4@�|E7��!?�c9{N8�@D�!�ٿ�s�Q��@:���4@�|E7��!?�c9{N8�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@��/)�ٿj�Ы�J�@�OI-r4@R qI��!?!4�ͮ�@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@(� ��ٿ_+�c���@m��ek4@@�\�!?%1"0���@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@��_��ٿI-i�7��@B��͠4@�-�~K�!?�>+̑�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@X�BX�ٿ�Og���@ܰ+M+4@�N�I�!?��9�F�@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@Hv���ٿc=�0���@���4@�2��{�!?f+��v��@�>Y}�ٿ�g��8�@@��z4@�#��s�!?3/�-�@���Ƀٿ_�;|�@�����4@䌞���!?~�s>���@���Ƀٿ_�;|�@�����4@䌞���!?~�s>���@�^ ��|ٿ�����@B�S��4@3�^��!?.ݧ�/�@�^ ��|ٿ�����@B�S��4@3�^��!?.ݧ�/�@����ٿ5.�����@ѩ�	4@���^��!?�2�����@����ٿ5.�����@ѩ�	4@���^��!?�2�����@i��b*�ٿ>���?�@ZT���4@(��c�!?`u��}�@i��b*�ٿ>���?�@ZT���4@(��c�!?`u��}�@i��b*�ٿ>���?�@ZT���4@(��c�!?`u��}�@i��b*�ٿ>���?�@ZT���4@(��c�!?`u��}�@i��b*�ٿ>���?�@ZT���4@(��c�!?`u��}�@IBW#�ٿ]##����@�z���4@����>�!?����B�@IBW#�ٿ]##����@�z���4@����>�!?����B�@IBW#�ٿ]##����@�z���4@����>�!?����B�@IBW#�ٿ]##����@�z���4@����>�!?����B�@�<���ٿ+�@0��@_o�X4@�ͧ��!?���&��@�<���ٿ+�@0��@_o�X4@�ͧ��!?���&��@�<���ٿ+�@0��@_o�X4@�ͧ��!?���&��@�<���ٿ+�@0��@_o�X4@�ͧ��!?���&��@���x^�ٿ�a�>VF�@w��6J4@-C,ِ!?w����|�@���x^�ٿ�a�>VF�@w��6J4@-C,ِ!?w����|�@��t�ٿ4q4��@:'5�4@ǡF֐!?�1�۞�@��t�ٿ4q4��@:'5�4@ǡF֐!?�1�۞�@��t�ٿ4q4��@:'5�4@ǡF֐!?�1�۞�@ӃNY$�ٿ8�+o$��@��R��4@d+���!?@�+���@ӃNY$�ٿ8�+o$��@��R��4@d+���!?@�+���@ӃNY$�ٿ8�+o$��@��R��4@d+���!?@�+���@ӃNY$�ٿ8�+o$��@��R��4@d+���!?@�+���@ӃNY$�ٿ8�+o$��@��R��4@d+���!?@�+���@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@t�x�ٿ��4��@z~�u4@�fZ��!?�.�b2�@�j�m��ٿ�_�����@#�7*��3@_�j��!?�
�� �@�j�m��ٿ�_�����@#�7*��3@_�j��!?�
�� �@�j�m��ٿ�_�����@#�7*��3@_�j��!?�
�� �@Ԛ Q�ٿ��)]�@����4@J3�1.�!?�ɾ���@�<�R;�ٿ��oy�^�@A��T�4@�\�c�!?+u �D�@�<�R;�ٿ��oy�^�@A��T�4@�\�c�!?+u �D�@�<�R;�ٿ��oy�^�@A��T�4@�\�c�!?+u �D�@w��&D�ٿ�6͌��@Qk=4@}�`�!?���'��@w��&D�ٿ�6͌��@Qk=4@}�`�!?���'��@w��&D�ٿ�6͌��@Qk=4@}�`�!?���'��@w��&D�ٿ�6͌��@Qk=4@}�`�!?���'��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@ݵsٿ3���B��@1fȒ4@������!?���P��@����4�ٿp]����@0�ƫ�4@0E:�А!?Rj��~��@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@氓r��ٿ^�N,�@�
��4@�M��!?F��2[�@|�o΅�ٿ��#�
P�@J}��[4@T!-��!?趦ɺ��@|�o΅�ٿ��#�
P�@J}��[4@T!-��!?趦ɺ��@|�o΅�ٿ��#�
P�@J}��[4@T!-��!?趦ɺ��@|�o΅�ٿ��#�
P�@J}��[4@T!-��!?趦ɺ��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@����ٿ��Hy�@��c$14@��F*}�!?�C<?Y��@{KR<P�ٿM�F�v�@:�OYc4@�ìwڐ!?C����1�@{KR<P�ٿM�F�v�@:�OYc4@�ìwڐ!?C����1�@{KR<P�ٿM�F�v�@:�OYc4@�ìwڐ!?C����1�@{KR<P�ٿM�F�v�@:�OYc4@�ìwڐ!?C����1�@{KR<P�ٿM�F�v�@:�OYc4@�ìwڐ!?C����1�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@���h�ٿ��誎��@�/�A=4@Y3�̸�!?hG�;�F�@-���_�ٿSLKg�@��yΕ4@�z>Ͷ�!?D*�Br��@�^��ŉٿB�ky���@��.��4@Z�O��!?��%y0��@�oʳ�ٿm������@�T�VR4@m��Ā�!?c�i�}��@�oʳ�ٿm������@�T�VR4@m��Ā�!?c�i�}��@�oʳ�ٿm������@�T�VR4@m��Ā�!?c�i�}��@w����ٿYi�f�q�@�(uw�4@���j��!?!q���|�@w����ٿYi�f�q�@�(uw�4@���j��!?!q���|�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@
Ŏ�Z�ٿ����m�@�o5l4@D01�Đ!?ඩܗ�@���m��ٿ�H�J��@\Pc(|4@���ϐ!?l�6sC��@���m��ٿ�H�J��@\Pc(|4@���ϐ!?l�6sC��@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@����{ٿ�:ۙ��@jhI+�4@-�}��!?�������@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��g��ٿ+��t��@�G��4@UJ�7��!?�4�ja��@��W�S�ٿ�d�T2�@��Z�4@?�d��!?�Z9��8�@��W�S�ٿ�d�T2�@��Z�4@?�d��!?�Z9��8�@��W�S�ٿ�d�T2�@��Z�4@?�d��!?�Z9��8�@��W�S�ٿ�d�T2�@��Z�4@?�d��!?�Z9��8�@��W�S�ٿ�d�T2�@��Z�4@?�d��!?�Z9��8�@ꍵ�?�ٿ�2dZB��@ ���4@�҈��!?'Q��*�@ꍵ�?�ٿ�2dZB��@ ���4@�҈��!?'Q��*�@ꍵ�?�ٿ�2dZB��@ ���4@�҈��!?'Q��*�@ꍵ�?�ٿ�2dZB��@ ���4@�҈��!?'Q��*�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@1J�/�ٿŻ\�*�@T`Q4@V�_l��!?Lj\)�D�@8A|��ٿls9��@����4@�G�!?]�^��@8A|��ٿls9��@����4@�G�!?]�^��@8A|��ٿls9��@����4@�G�!?]�^��@_��HшٿoZ� :Q�@�Ct4@i�+,�!?��!WJW�@_��HшٿoZ� :Q�@�Ct4@i�+,�!?��!WJW�@_��HшٿoZ� :Q�@�Ct4@i�+,�!?��!WJW�@��_�ٿ���'�C�@V���94@�Zr��!?(�۷N��@��_�ٿ���'�C�@V���94@�Zr��!?(�۷N��@$���ٿt�ղI�@��G�	4@j�d��!?1*�Pcc�@eԈ��ٿ UG�@�(�� 4@ַ� �!?H�Վ!�@eԈ��ٿ UG�@�(�� 4@ַ� �!?H�Վ!�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@~�L���ٿ�1*\��@fxYR4@��t�+�!?Oa��I�@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@���,�ٿ��*�	�@�%8�C4@* �Đ!?�� ��@$O1�ٿ��K4�7�@�8�Հ4@��|���!?S���א�@$O1�ٿ��K4�7�@�8�Հ4@��|���!?S���א�@�Hi��ٿ�	G���@�:�L�4@�u.癐!?�U*�c�@`u�}�ٿ��~����@���,Z4@��
�!?��SY�@`u�}�ٿ��~����@���,Z4@��
�!?��SY�@`u�}�ٿ��~����@���,Z4@��
�!?��SY�@`u�}�ٿ��~����@���,Z4@��
�!?��SY�@`u�}�ٿ��~����@���,Z4@��
�!?��SY�@]�.�ٿ�3�
P��@i'IZ�4@�8���!?bpu%&��@]�.�ٿ�3�
P��@i'IZ�4@�8���!?bpu%&��@]�.�ٿ�3�
P��@i'IZ�4@�8���!?bpu%&��@�ٿ�E�����@�@�#4@1��u�!?D��Ӽ�@�ٿ�E�����@�@�#4@1��u�!?D��Ӽ�@�ٿ�E�����@�@�#4@1��u�!?D��Ӽ�@�ٿ�E�����@�@�#4@1��u�!?D��Ӽ�@�ٿ�E�����@�@�#4@1��u�!?D��Ӽ�@@CΠ��ٿj6�g���@F�x�4@��.�!?�(��8�@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@o��I0�ٿ�Bx���@��N7
4@6H����!?�r�%��@���@,�ٿf����I�@t4؍4@�uж�!?��wa��@�r�oq�ٿh���^�@6�e4@|7�i�!?�>0�0�@�r�oq�ٿh���^�@6�e4@|7�i�!?�>0�0�@y��	��ٿ4�K�W�@�Oȱ`4@�s�!?2�J����@y��	��ٿ4�K�W�@�Oȱ`4@�s�!?2�J����@y��	��ٿ4�K�W�@�Oȱ`4@�s�!?2�J����@y��	��ٿ4�K�W�@�Oȱ`4@�s�!?2�J����@y��	��ٿ4�K�W�@�Oȱ`4@�s�!?2�J����@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@\ ��l�ٿP��R^��@��iYh4@Vv����!?!�Eg��@�:�^�ٿ�%�*Q�@2<��w4@_�}��!?��E�G�@��O��ٿ����A�@u&��94@�<1ox�!?J���@��O��ٿ����A�@u&��94@�<1ox�!?J���@��O��ٿ����A�@u&��94@�<1ox�!?J���@��O��ٿ����A�@u&��94@�<1ox�!?J���@��O��ٿ����A�@u&��94@�<1ox�!?J���@��O��ٿ����A�@u&��94@�<1ox�!?J���@���(.�ٿ@>XÊ�@K'`�o4@^`/縷!?���1��@���(.�ٿ@>XÊ�@K'`�o4@^`/縷!?���1��@���(.�ٿ@>XÊ�@K'`�o4@^`/縷!?���1��@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@�g��]�ٿڴ8��@�3���4@ח��א!?��9ǯ@�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@x"�q�ٿ��:�Q�@��tk
4@�9z���!?d�=�%K�@>��@��ٿ�S�9��@Ü�l%4@9���!?�N���d�@>��@��ٿ�S�9��@Ü�l%4@9���!?�N���d�@>��@��ٿ�S�9��@Ü�l%4@9���!?�N���d�@>��@��ٿ�S�9��@Ü�l%4@9���!?�N���d�@,��ܨ�ٿR�p���@qe�|�4@"�p�!?���3o�@,��ܨ�ٿR�p���@qe�|�4@"�p�!?���3o�@,��ܨ�ٿR�p���@qe�|�4@"�p�!?���3o�@,��ܨ�ٿR�p���@qe�|�4@"�p�!?���3o�@,��ܨ�ٿR�p���@qe�|�4@"�p�!?���3o�@�myLc�ٿMwP���@�N���4@3��轐!?��wA%H�@�myLc�ٿMwP���@�N���4@3��轐!?��wA%H�@�myLc�ٿMwP���@�N���4@3��轐!?��wA%H�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@"y�O�ٿ��}b�@e͟��4@e�g��!?0�f�0f�@E%�ٿ%<����@4�C`f4@���_��!?�Ǐ����@E%�ٿ%<����@4�C`f4@���_��!?�Ǐ����@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@PO�W�ٿ+��R�@W���,4@-�'Ѭ�!?Sx[�Z�@9����ٿHB��+�@pߋ��4@_� i�!?7bf��$�@9����ٿHB��+�@pߋ��4@_� i�!?7bf��$�@9����ٿHB��+�@pߋ��4@_� i�!?7bf��$�@9����ٿHB��+�@pߋ��4@_� i�!?7bf��$�@��t��ٿ�L�Y���@�8�7�4@zz6LG�!?��Vt`�@z�F���ٿ�6P3w�@Z�2I4@��Jm�!?J��|��@z�F���ٿ�6P3w�@Z�2I4@��Jm�!?J��|��@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@�|{
�ٿ~�]���@0�w�4@I@�T��!?7�k�T�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@���ݏٿ>b����@ߎ�� 4@���Eʐ!?<�Ϙ�^�@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@����ٿ��z�	��@��/4@7$�ͪ�!?kd\2��@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@�~�l�ٿ�\|h��@&�:�E4@��R�l�!?Ic��q�@`wI|a�ٿ�	�v��@p	��4@i���Ð!?0	]�@��0A��ٿ�i���@�n��4@O7)��!?�(��Ҭ�@��0A��ٿ�i���@�n��4@O7)��!?�(��Ҭ�@��0A��ٿ�i���@�n��4@O7)��!?�(��Ҭ�@	rS�3�ٿ|fW���@S�c�4@�8��̐!?���=T�@	rS�3�ٿ|fW���@S�c�4@�8��̐!?���=T�@	rS�3�ٿ|fW���@S�c�4@�8��̐!?���=T�@	rS�3�ٿ|fW���@S�c�4@�8��̐!?���=T�@	rS�3�ٿ|fW���@S�c�4@�8��̐!?���=T�@.̠	�ٿ990��,�@�'�+�4@&޸��!?��c	�@.̠	�ٿ990��,�@�'�+�4@&޸��!?��c	�@.̠	�ٿ990��,�@�'�+�4@&޸��!?��c	�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@G/~� �ٿY`�r���@�-� 4@NJq�ː!?~��=�@E�Z&%�ٿJF�8���@�'j�)4@���А!?��:aH#�@�!WD��ٿ��z�?��@(�{�4@W�q�ݐ!?�,1R�@�!WD��ٿ��z�?��@(�{�4@W�q�ݐ!?�,1R�@�!WD��ٿ��z�?��@(�{�4@W�q�ݐ!?�,1R�@�!WD��ٿ��z�?��@(�{�4@W�q�ݐ!?�,1R�@�!WD��ٿ��z�?��@(�{�4@W�q�ݐ!?�,1R�@�ȍ
R�ٿ�,��\��@�5^34@*#4��!?�ڡ�}�@�ȍ
R�ٿ�,��\��@�5^34@*#4��!?�ڡ�}�@�ȍ
R�ٿ�,��\��@�5^34@*#4��!?�ڡ�}�@�ȍ
R�ٿ�,��\��@�5^34@*#4��!?�ڡ�}�@w��77�ٿ�Nl���@�Y���4@+1���!?l��$��@�?}�(�ٿ]b�i���@y��I4@i��t*�!?�<*���@�?}�(�ٿ]b�i���@y��I4@i��t*�!?�<*���@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@&<�ƍٿ\C����@����4@�ؐ!?:����@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@�H�ٿ\��s+��@�͈e-4@y�k�!?��!<���@-�<�ٿ��P��c�@�?>� 4@��[�!??��F���@-�<�ٿ��P��c�@�?>� 4@��[�!??��F���@u��}ٿ�,��O�@�Rn��4@�]R��!?��b��@l��.��ٿ��'��@���4@������!?�����@l��.��ٿ��'��@���4@������!?�����@6���W}ٿ��oK@��@��Ѡ�4@G�̽�!?�5z��t�@6���W}ٿ��oK@��@��Ѡ�4@G�̽�!?�5z��t�@6���W}ٿ��oK@��@��Ѡ�4@G�̽�!?�5z��t�@6���W}ٿ��oK@��@��Ѡ�4@G�̽�!?�5z��t�@6���W}ٿ��oK@��@��Ѡ�4@G�̽�!?�5z��t�@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@��|,�~ٿ��Cx@8�@�#���4@�Q�1v�!?������@�O��9�ٿ.��=�@R )�4@�2v�!?*븭���@�O��9�ٿ.��=�@R )�4@�2v�!?*븭���@�7�yٿ�2�̹�@���54@&��͐!?�������@�7�yٿ�2�̹�@���54@&��͐!?�������@ۙRif�ٿ�I�5��@�6��4@��Gެ�!?�2/$��@ۙRif�ٿ�I�5��@�6��4@��Gެ�!?�2/$��@ۙRif�ٿ�I�5��@�6��4@��Gެ�!?�2/$��@W1bf�ٿ�2��v��@ȭ�4@�a�֎�!?�ޛm�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@��C�/�ٿ�+y�S�@%���4@�t�	��!?كef�V�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@K
1چٿ�	A�o�@Ƌ�״4@O�)�l�!?,0x�m,�@��.�ٿo�O"{j�@����4@.�n�q�!?�O��"}�@��.�ٿo�O"{j�@����4@.�n�q�!?�O��"}�@�g�)Z�ٿ��M���@g�eME4@4��{�!?��@��@~3^�ٿ������@a���4@l1y-͐!?��
�a�@~3^�ٿ������@a���4@l1y-͐!?��
�a�@T��R�ٿXp|���@r�CDi4@r����!?����@�@k�����ٿ�M#����@uIqx4@��V7'�!?�:%�qn�@k�����ٿ�M#����@uIqx4@��V7'�!?�:%�qn�@3�8ٿ�)����@�S��M4@
��z'�!?��?L��@3�8ٿ�)����@�S��M4@
��z'�!?��?L��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@Yi�˄ٿ�;�����@�.�J.4@��`c	�!?v��9��@��7�Q�ٿ��ڕ�{�@1?zg�	4@�^W���!?q�nX��@8"��ٿ��0�q�@k�G<4@��ґ��!?�Vc��@8"��ٿ��0�q�@k�G<4@��ґ��!?�Vc��@8"��ٿ��0�q�@k�G<4@��ґ��!?�Vc��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@;�$(��ٿ������@C�@�4@�NN��!?Ŝ��-��@�wF��ٿY�$��@�#��v4@#공�!?jض����@z�w�ٿX^����@<����4@AU�!?�^���@z�w�ٿX^����@<����4@AU�!?�^���@z�w�ٿX^����@<����4@AU�!?�^���@z�w�ٿX^����@<����4@AU�!?�^���@z�w�ٿX^����@<����4@AU�!?�^���@z�w�ٿX^����@<����4@AU�!?�^���@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@1��E8�ٿ^n�ص��@0���n4@o��~Ґ!?&j��N�@��)u�ٿ��`o8�@��i4@N��h�!??=-�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@�F�Oυٿ�@c	��@��04@���VT�!?�XۜI�@��I�B�ٿ�,Х�+�@߀���4@���C��!? �J%�N�@��I�B�ٿ�,Х�+�@߀���4@���C��!? �J%�N�@��I�B�ٿ�,Х�+�@߀���4@���C��!? �J%�N�@��I�B�ٿ�,Х�+�@߀���4@���C��!? �J%�N�@�^���ٿ��շY��@��f�4@��@�!?�e=��@�^���ٿ��շY��@��f�4@��@�!?�e=��@3�ه�ٿ5w(����@�~��{4@����L�!?�/o \�@3�ه�ٿ5w(����@�~��{4@����L�!?�/o \�@��5R��ٿ��9r��@�
8ۈ4@6�A��!?�&"��@��z| �ٿ���V���@_(�94@������!?a
$���@��z| �ٿ���V���@_(�94@������!?a
$���@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@_�]e�ٿ[��& �@S���
4@�Y���!?"F3O��@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@�|ez��ٿdB�[�@u�h�4@v2����!?�BWFP�@��-�ٿÕ���f�@(*��	4@�����!?�r�@+��@��-�ٿÕ���f�@(*��	4@�����!?�r�@+��@�@Ȇٿ�a	��@��F��4@����!?N���E�@�@Ȇٿ�a	��@��F��4@����!?N���E�@�@Ȇٿ�a	��@��F��4@����!?N���E�@�@Ȇٿ�a	��@��F��4@����!?N���E�@�@Ȇٿ�a	��@��F��4@����!?N���E�@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@�C?+��ٿ�O&G��@�jG�{4@�����!?��<N���@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@%�`��ٿ�`�H��@ݭ�G�4@._ �Ր!?o!�Ά7�@��VLȁٿ�$�@^�*�K4@`�U ��!?Ng�ʨ�@��VLȁٿ�$�@^�*�K4@`�U ��!?Ng�ʨ�@
�GvЂٿ���,��@ij���4@	B���!?�bRF���@
�GvЂٿ���,��@ij���4@	B���!?�bRF���@
�GvЂٿ���,��@ij���4@	B���!?�bRF���@
�GvЂٿ���,��@ij���4@	B���!?�bRF���@
�GvЂٿ���,��@ij���4@	B���!?�bRF���@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@�"�[I�ٿ������@0�=�>4@�r-Ր!?x6�YIO�@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@+<7�T�ٿ~U^e�@��`�4@|.���!?�͇v��@���ԍٿ5N����@�m��h4@6-�Ð!?hN��S�@���ԍٿ5N����@�m��h4@6-�Ð!?hN��S�@���ԍٿ5N����@�m��h4@6-�Ð!?hN��S�@���ԍٿ5N����@�m��h4@6-�Ð!?hN��S�@���ԍٿ5N����@�m��h4@6-�Ð!?hN��S�@Х�ٿ����t�@;ݦk4@�kЎ�!?��LF���@Х�ٿ����t�@;ݦk4@�kЎ�!?��LF���@Х�ٿ����t�@;ݦk4@�kЎ�!?��LF���@<I���ٿ�W|��^�@��h��4@z����!?rOO��@<I���ٿ�W|��^�@��h��4@z����!?rOO��@<I���ٿ�W|��^�@��h��4@z����!?rOO��@<I���ٿ�W|��^�@��h��4@z����!?rOO��@c�"o؄ٿ6����@](�D4@2� ��!?��U����@c�"o؄ٿ6����@](�D4@2� ��!?��U����@c�"o؄ٿ6����@](�D4@2� ��!?��U����@c�"o؄ٿ6����@](�D4@2� ��!?��U����@nJR�ٿ�$���@���^4@���V��!?���S�F�@nJR�ٿ�$���@���^4@���V��!?���S�F�@nJR�ٿ�$���@���^4@���V��!?���S�F�@nJR�ٿ�$���@���^4@���V��!?���S�F�@nJR�ٿ�$���@���^4@���V��!?���S�F�@i53iٿ2�龞��@I�G��4@V� ���!?�m<���@i53iٿ2�龞��@I�G��4@V� ���!?�m<���@�C.4�{ٿ�@ѯ�@6%y^C4@�.Z��!?dBu;���@�C.4�{ٿ�@ѯ�@6%y^C4@�.Z��!?dBu;���@�C.4�{ٿ�@ѯ�@6%y^C4@�.Z��!?dBu;���@�C.4�{ٿ�@ѯ�@6%y^C4@�.Z��!?dBu;���@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@�܊)�~ٿiK��	l�@��r �4@m�,)��!?�j]B=)�@jo�_�ٿ�ʚ����@��b��4@�����!?�v�c��@jo�_�ٿ�ʚ����@��b��4@�����!?�v�c��@jo�_�ٿ�ʚ����@��b��4@�����!?�v�c��@)�ZM�ٿ�3q%�x�@�/AyP4@�����!?��\%�C�@)�ZM�ٿ�3q%�x�@�/AyP4@�����!?��\%�C�@c��_�ٿJm�����@�	Q��4@�(���!?�u
BM�@��G��ٿ��3ˁ�@�;��4@����w�!?փka���@PRy�/�ٿn���E�@-��R�4@��O�1�!?w"�๤�@+��d	�ٿ�P ����@�@��4@���̐!?b�x��p�@+��d	�ٿ�P ����@�@��4@���̐!?b�x��p�@+��d	�ٿ�P ����@�@��4@���̐!?b�x��p�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@�j灅ٿI:xi?�@+�z��4@� ���!?B���(T�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@S�P�@�ٿ;��9���@�~�H�4@Q���!?q���[�@x_PtF�ٿ�-�D]!�@�4��4@����!?:q����@x_PtF�ٿ�-�D]!�@�4��4@����!?:q����@x_PtF�ٿ�-�D]!�@�4��4@����!?:q����@x_PtF�ٿ�-�D]!�@�4��4@����!?:q����@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@q� �}ٿ��$���@NѠA�4@K7�H��!?za4M��@�9���ٿ(�}^]�@E?�Uf4@�鿮o�!?��q����@�9���ٿ(�}^]�@E?�Uf4@�鿮o�!?��q����@�9���ٿ(�}^]�@E?�Uf4@�鿮o�!?��q����@�9���ٿ(�}^]�@E?�Uf4@�鿮o�!?��q����@�9���ٿ(�}^]�@E?�Uf4@�鿮o�!?��q����@�]��}ٿ�yս��@A�*O�4@]���!?A�z�@�]��}ٿ�yս��@A�*O�4@]���!?A�z�@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@��G��~ٿ�V�@����4@)�/�ڐ!?8S��+��@VK�$�ٿ��|����@��<�4@I^e	�!?S�a�\f�@VK�$�ٿ��|����@��<�4@I^e	�!?S�a�\f�@VK�$�ٿ��|����@��<�4@I^e	�!?S�a�\f�@����	�ٿ,�9���@h��94@,c�0͐!?
u��V�@����	�ٿ,�9���@h��94@,c�0͐!?
u��V�@����	�ٿ,�9���@h��94@,c�0͐!?
u��V�@����	�ٿ,�9���@h��94@,c�0͐!?
u��V�@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���+�ٿ�HJc�|�@ˢ��4@�ktא!?Э`��@���ٿ}p�z6V�@�&����3@�����!?�ŇX+�@���ٿ}p�z6V�@�&����3@�����!?�ŇX+�@���ٿ}p�z6V�@�&����3@�����!?�ŇX+�@���ٿ}p�z6V�@�&����3@�����!?�ŇX+�@���e�ٿ���?�@�0Id4@����!?��BJo�@���e�ٿ���?�@�0Id4@����!?��BJo�@���e�ٿ���?�@�0Id4@����!?��BJo�@���e�ٿ���?�@�0Id4@����!?��BJo�@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@�᎜�ٿ�f���7�@�ѩn4@SB�j��!?gŦ���@���_Z�ٿ0bg�8�@%i8��4@5� '��!?�"��P��@�<d뗈ٿ�p�t��@ZQ4@�n�R�!?��J���@�Y�~ٿ����}��@�P�U4@F~4;��!?��9YC
�@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@cVp�^�ٿ�9����@4X4@�:z�!?�L��n��@�L:7�|ٿ���[�	�@H�}1�4@F��7�!?4�ij���@�L:7�|ٿ���[�	�@H�}1�4@F��7�!?4�ij���@�L:7�|ٿ���[�	�@H�}1�4@F��7�!?4�ij���@�sT�}ٿNJ�c���@�=��4@cLgI�!?韧���@��)4�ٿ�	M���@�����4@Է��!?��B����@��)4�ٿ�	M���@�����4@Է��!?��B����@��)4�ٿ�	M���@�����4@Է��!?��B����@��)4�ٿ�	M���@�����4@Է��!?��B����@��)4�ٿ�	M���@�����4@Է��!?��B����@��)4�ٿ�	M���@�����4@Է��!?��B����@�}�ٿ ������@Πic4@���`ِ!?�?ի���@�}�ٿ ������@Πic4@���`ِ!?�?ի���@�}�ٿ ������@Πic4@���`ِ!?�?ի���@�}�ٿ ������@Πic4@���`ِ!?�?ի���@�}�ٿ ������@Πic4@���`ِ!?�?ի���@�}�ٿ ������@Πic4@���`ِ!?�?ի���@Qw'��ٿŻwم��@|I�<?4@n�C*��!?������@Qw'��ٿŻwم��@|I�<?4@n�C*��!?������@�b4|ٿ����~�@`�N��4@FJ4���!?��vZ�B�@�b4|ٿ����~�@`�N��4@FJ4���!?��vZ�B�@�,�R|ٿ�JF*n2�@�24@�o��,�!?��g"�@�,�R|ٿ�JF*n2�@�24@�o��,�!?��g"�@�,�R|ٿ�JF*n2�@�24@�o��,�!?��g"�@�,�R|ٿ�JF*n2�@�24@�o��,�!?��g"�@�,�R|ٿ�JF*n2�@�24@�o��,�!?��g"�@���d4�ٿ���~��@���]4@�����!?��C��s�@���d4�ٿ���~��@���]4@�����!?��C��s�@���d4�ٿ���~��@���]4@�����!?��C��s�@��x�4�ٿ�#�����@^�ם4@�#z�!?t1%���@��x�4�ٿ�#�����@^�ם4@�#z�!?t1%���@�k�&�ٿ���زz�@��5.&4@0�L �!?	s��@�k�&�ٿ���زz�@��5.&4@0�L �!?	s��@�k�&�ٿ���زz�@��5.&4@0�L �!?	s��@k9�5�ٿ����k�@E"v^4@�ؔ(��!?*����@k9�5�ٿ����k�@E"v^4@�ؔ(��!?*����@�,�Ƅٿ`�<@�$�@]�	�4@�z��!?+�߾���@���H$zٿ�oW,�@���4@��_-��!?�V�\u�@1��V̂ٿґH!%�@�X^N4@
u�}�!?�PG �@1��V̂ٿґH!%�@�X^N4@
u�}�!?�PG �@9L����ٿ���@�"��4@e�f��!?֊�	@�@9L����ٿ���@�"��4@e�f��!?֊�	@�@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@J� �7�ٿ�1����@�d��&4@�����!?�yt e��@]��G�ٿ^1v���@�2̔�4@X�z���!?��2r$�@]��G�ٿ^1v���@�2̔�4@X�z���!?��2r$�@]��G�ٿ^1v���@�2̔�4@X�z���!?��2r$�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@����ٿ#k�&�@H�ڂ�4@�S���!?�0���}�@'���ƅٿBe2{��@�H���4@��,Dk�!?���I8H�@'���ƅٿBe2{��@�H���4@��,Dk�!?���I8H�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��&��ٿ��^1��@	����4@�)%�=�!?���r%�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@��V���ٿ�o�L�@n�1ɼ4@�pٌ�!?0%4f�&�@�L�Ԓٿ��S����@YQ	t�4@�=��!?sL-��2�@�L�Ԓٿ��S����@YQ	t�4@�=��!?sL-��2�@�L�Ԓٿ��S����@YQ	t�4@�=��!?sL-��2�@�,�e�ٿ�D�����@��C�4@r0�!?%ғ��@��ږ��ٿط�#�@�ud�	4@�7O�V�!?�^���@��ږ��ٿط�#�@�ud�	4@�7O�V�!?�^���@��ږ��ٿط�#�@�ud�	4@�7O�V�!?�^���@g=���ٿ '���y�@��tw4@�ԁM�!?Ta�*�q�@g=���ٿ '���y�@��tw4@�ԁM�!?Ta�*�q�@g=���ٿ '���y�@��tw4@�ԁM�!?Ta�*�q�@%ǫ��ٿM2���z�@�۟��4@�ns�7�!?H.묤�@gX[�<�ٿ�x�2y��@l%��4@#�1�&�!?WϢO��@gX[�<�ٿ�x�2y��@l%��4@#�1�&�!?WϢO��@gX[�<�ٿ�x�2y��@l%��4@#�1�&�!?WϢO��@\���ٿ��h<ɕ�@	�-2�3@�����!?��z�ó�@�ph�x�ٿ��w�^+�@�I�3@\&!��!?T��GE�@�ph�x�ٿ��w�^+�@�I�3@\&!��!?T��GE�@�ph�x�ٿ��w�^+�@�I�3@\&!��!?T��GE�@�ph�x�ٿ��w�^+�@�I�3@\&!��!?T��GE�@�ph�x�ٿ��w�^+�@�I�3@\&!��!?T��GE�@g�e�ٿTF:wth�@���'P4@��*���!?�|j�W(�@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@kn4<�ٿ��C���@rԎN4@�xG�ؐ!?�������@��Q�ƃٿ˘P-���@[a ��4@ϸ�A�!?B�[YN��@��l�Ղٿ�	�9q�@;/P�L4@�;���!?b��C/H�@��l�Ղٿ�	�9q�@;/P�L4@�;���!?b��C/H�@��l�Ղٿ�	�9q�@;/P�L4@�;���!?b��C/H�@��l�Ղٿ�	�9q�@;/P�L4@�;���!?b��C/H�@l�T�ٿ��A���@X�� A4@\ᜫ�!?���M�w�@�{l�փٿ�-�c5�@�E�4@���b��!?MS�-�8�@�{l�փٿ�-�c5�@�E�4@���b��!?MS�-�8�@�{l�փٿ�-�c5�@�E�4@���b��!?MS�-�8�@�{l�փٿ�-�c5�@�E�4@���b��!?MS�-�8�@�{l�փٿ�-�c5�@�E�4@���b��!?MS�-�8�@��ٿك���i�@�[�4@9qW���!?�Ь��@�T�E~ٿ�{(��@cG2�54@���}�!?�v�%8��@�T�E~ٿ�{(��@cG2�54@���}�!?�v�%8��@�T�E~ٿ�{(��@cG2�54@���}�!?�v�%8��@�f.�ٿܭ���P�@Y���4@��S��!?�^�c��@�f.�ٿܭ���P�@Y���4@��S��!?�^�c��@�f.�ٿܭ���P�@Y���4@��S��!?�^�c��@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@���t��ٿ���NZr�@1�ݴ�4@ٜ����!?�%y���@�=�H�ٿ�Ԧ��@=�b	4@οM	��!?���i�-�@�=�H�ٿ�Ԧ��@=�b	4@οM	��!?���i�-�@�=�H�ٿ�Ԧ��@=�b	4@οM	��!?���i�-�@�=�H�ٿ�Ԧ��@=�b	4@οM	��!?���i�-�@�=�H�ٿ�Ԧ��@=�b	4@οM	��!?���i�-�@�V,���ٿG���@�u?4@\�E`��!?t�}Ph��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@vl6��ٿ�/	P��@�D�m�4@I*ۜ�!?�!��@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@�$Q���ٿ�Fb$���@y�$�4@�;f�!?Ӏ>z�@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@5K0���ٿ\�K[h�@��y��4@hE���!?��Ue��@KX�]��ٿE��w���@��e�4@���א!?�=�2�@����ٿ�MiF �@��v�84@�]�ǌ�!?����c��@y��U�ٿ?|E�2�@�.jٱ 4@�[��w�!?�Cd���@y��U�ٿ?|E�2�@�.jٱ 4@�[��w�!?�Cd���@cԆl�ٿ4\�j7��@\�w 4@B�V��!?6��孾�@cԆl�ٿ4\�j7��@\�w 4@B�V��!?6��孾�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@���ٿ�G���@�B��4@2g�Ŷ�!?�rWUT�@C��ٿX��P��@\9*��4@P�m��!?ޤ���	�@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@����A�ٿ�^�^���@�l�4@�q�&ߐ!?F��r��@׫�ٿ�So���@\c�4@s�p��!?�4�w��@�gO���ٿ��^��@5�[4@~$o�"�!?vp�?�@�gO���ٿ��^��@5�[4@~$o�"�!?vp�?�@�gO���ٿ��^��@5�[4@~$o�"�!?vp�?�@��à�ٿ���kd=�@D<���4@��U�!?y�w�@��/ִ�ٿ����%��@sz�I%4@BT��!?���o��@��ع�ٿ�N��0�@�[�W74@_	R�!?H`>��s�@��ع�ٿ�N��0�@�[�W74@_	R�!?H`>��s�@���`��ٿ
�[5M8�@�NI>4@�T|���!?#
#;p�@���`��ٿ
�[5M8�@�NI>4@�T|���!?#
#;p�@�?O�Ѕٿ���=�@�r� 4@y�ϻ�!?�p�e+�@�?O�Ѕٿ���=�@�r� 4@y�ϻ�!?�p�e+�@�?O�Ѕٿ���=�@�r� 4@y�ϻ�!?�p�e+�@E�WY��ٿ�u[E��@>�,�� 4@��!?��i��@E�WY��ٿ�u[E��@>�,�� 4@��!?��i��@E�WY��ٿ�u[E��@>�,�� 4@��!?��i��@E�WY��ٿ�u[E��@>�,�� 4@��!?��i��@�8P
yٿ�J�����@j���M4@����!?9���YB�@�8P
yٿ�J�����@j���M4@����!?9���YB�@߿-{ٿ�ѐ���@;*�84@�"�
�!?h̯�)�@߿-{ٿ�ѐ���@;*�84@�"�
�!?h̯�)�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@�|��ǀٿM�Ƕ��@���o�4@��Rd�!?�Q�	~]�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@;����ٿ�]�K���@���1�4@.�A�$�!?�BUs�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@�Y����ٿ�6�iG��@�js� 4@R���֐!?xK_"�a�@7�r�U�ٿ=�YDz��@�h���4@���ǐ!?1�6E
�@7�r�U�ٿ=�YDz��@�h���4@���ǐ!?1�6E
�@7�r�U�ٿ=�YDz��@�h���4@���ǐ!?1�6E
�@_�&O�ٿ?�V=9��@�bV.4@y/�!?<g���@��F�	�ٿ"!���e�@M��L4@�U ��!?�Q�u	��@��F�	�ٿ"!���e�@M��L4@�U ��!?�Q�u	��@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@_j ۉ�ٿ�&^�}�@ت�4@�~s�!?călzR�@�h�b�ٿӿ�ǎ��@�~Xt 4@�5է�!?ܱdU_�@��>T�ٿ�WDA�@��y��3@s�ᘐ!?�dxDL �@Ҡ7���ٿU�pw%��@ӄ�C4@�����!?�`�0Qi�@Ҡ7���ٿU�pw%��@ӄ�C4@�����!?�`�0Qi�@Ҡ7���ٿU�pw%��@ӄ�C4@�����!?�`�0Qi�@co�q�ٿ�˅�Y��@�rw;�4@"&c��!?޻;��@co�q�ٿ�˅�Y��@�rw;�4@"&c��!?޻;��@co�q�ٿ�˅�Y��@�rw;�4@"&c��!?޻;��@co�q�ٿ�˅�Y��@�rw;�4@"&c��!?޻;��@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@0tI}3�ٿ0�B��@�����4@g�݋�!?�̒o���@���ٿ�7���M�@'��g4@����d�!?�&=6���@���ٿ�7���M�@'��g4@����d�!?�&=6���@���ٿ�7���M�@'��g4@����d�!?�&=6���@���ٿ�7���M�@'��g4@����d�!?�&=6���@���ٿ�7���M�@'��g4@����d�!?�&=6���@���ٿ�7���M�@'��g4@����d�!?�&=6���@�b��ٿY�ͬ�@^��ԟ4@~Zeh��!?y�.�@�b��ٿY�ͬ�@^��ԟ4@~Zeh��!?y�.�@�b��ٿY�ͬ�@^��ԟ4@~Zeh��!?y�.�@�|r_/�ٿf\����@K��P4@���!?�_ ��T�@�|r_/�ٿf\����@K��P4@���!?�_ ��T�@�|r_/�ٿf\����@K��P4@���!?�_ ��T�@�|r_/�ٿf\����@K��P4@���!?�_ ��T�@�|r_/�ٿf\����@K��P4@���!?�_ ��T�@`A���~ٿ���ֻ��@S/L,4@��1��!?���ɛ�@`A���~ٿ���ֻ��@S/L,4@��1��!?���ɛ�@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@?L1�ٿ��8Pf��@�(����3@�ے��!?M�����@BG��ٿ��MbL$�@�wŕ4@�@��v�!?�<�!E�@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@C#�/X�ٿs�AI��@э���4@� ݄��!?�i?���@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@]�G|ǎٿ#ގ���@�ps�4@b/W�u�!?��z=�C�@�YM�a�ٿ6<a���@{k[4@Kv�	�!?�����@�ζH�ٿYT��܋�@�jU�34@�TM���!?��T���@�ζH�ٿYT��܋�@�jU�34@�TM���!?��T���@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@$:-�ٿ��j>u�@�nb4@X}3���!?a[��T�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�d�[��ٿU������@@
\4@�iy��!?૜�n~�@�#y7�ٿ���E��@9�W*�4@�m��!?8i�Zf��@�#y7�ٿ���E��@9�W*�4@�m��!?8i�Zf��@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@LSƅٿ'� ����@xzX�4@Έ��?�!?E���K�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@U�q/�ٿE���@6��4@6�/��!?ya;�47�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@�����ٿ�>�.ͷ�@��z��4@��㳐!?%C;�&�@[lT��ٿl:�A��@o���4@�XVt�!?Lvz[�@[lT��ٿl:�A��@o���4@�XVt�!?Lvz[�@[lT��ٿl:�A��@o���4@�XVt�!?Lvz[�@�p��j�ٿK��\ޮ�@L���4@&��!��!?�mN��@�p��j�ٿK��\ޮ�@L���4@&��!��!?�mN��@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@�u��ٿ,��M��@T�%ls4@ߏ9�!?w*{
���@[�uG�ٿ0���D��@Cw��y4@0�����!?�����@[�uG�ٿ0���D��@Cw��y4@0�����!?�����@��%iՇٿ�;��@�u���4@GI�>�!?^��}�{�@��%iՇٿ�;��@�u���4@GI�>�!?^��}�{�@��%iՇٿ�;��@�u���4@GI�>�!?^��}�{�@bT���ٿ�<�!��@
�Y�B4@�u�ɐ!?�T�m�@bT���ٿ�<�!��@
�Y�B4@�u�ɐ!?�T�m�@bT���ٿ�<�!��@
�Y�B4@�u�ɐ!?�T�m�@vx�
�ٿu�$*/��@6%oj4@�蹃��!?{N��M[�@vx�
�ٿu�$*/��@6%oj4@�蹃��!?{N��M[�@vx�
�ٿu�$*/��@6%oj4@�蹃��!?{N��M[�@vx�
�ٿu�$*/��@6%oj4@�蹃��!?{N��M[�@V�gJ2�ٿ?܇=���@���M�4@H`4�!?8=�����@V�gJ2�ٿ?܇=���@���M�4@H`4�!?8=�����@5���ٿwu�i?��@�0���3@����!?����8��@5���ٿwu�i?��@�0���3@����!?����8��@5���ٿwu�i?��@�0���3@����!?����8��@5���ٿwu�i?��@�0���3@����!?����8��@5���ٿwu�i?��@�0���3@����!?����8��@WmF�I�ٿ�bȉ��@��a+��3@��I�d�!?`P��i��@WmF�I�ٿ�bȉ��@��a+��3@��I�d�!?`P��i��@WmF�I�ٿ�bȉ��@��a+��3@��I�d�!?`P��i��@WmF�I�ٿ�bȉ��@��a+��3@��I�d�!?`P��i��@WmF�I�ٿ�bȉ��@��a+��3@��I�d�!?`P��i��@�D[pu�ٿ���7Ȣ�@��6��3@*��ʐ!?Vl�AYf�@�����ٿ�3�@�@�{��B�3@���!?9ضGD4�@��VD}�ٿ�bj}��@��ֹ��3@���&5�!?�s�����@��VD}�ٿ�bj}��@��ֹ��3@���&5�!?�s�����@��VD}�ٿ�bj}��@��ֹ��3@���&5�!?�s�����@��VD}�ٿ�bj}��@��ֹ��3@���&5�!?�s�����@��VD}�ٿ�bj}��@��ֹ��3@���&5�!?�s�����@����ŕٿ���m��@�}P5H4@��{O%�!?{ժ9��@����ŕٿ���m��@�}P5H4@��{O%�!?{ժ9��@����ŕٿ���m��@�}P5H4@��{O%�!?{ժ9��@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�(HR͖ٿv��X5�@�Z��4@��:��!?J
�0�@�%4�ٿF�3�1\�@1ʑ4@�r]⽐!?���>E��@�%4�ٿF�3�1\�@1ʑ4@�r]⽐!?���>E��@�%4�ٿF�3�1\�@1ʑ4@�r]⽐!?���>E��@��i��ٿ�:��xI�@�	H#�3@`u�o�!?ݰ�Ӭ�@��i��ٿ�:��xI�@�	H#�3@`u�o�!?ݰ�Ӭ�@��i��ٿ�:��xI�@�	H#�3@`u�o�!?ݰ�Ӭ�@��i��ٿ�:��xI�@�	H#�3@`u�o�!?ݰ�Ӭ�@��i��ٿ�:��xI�@�	H#�3@`u�o�!?ݰ�Ӭ�@91���ٿ�|��@)�cw� 4@�$�<��!??J�V���@91���ٿ�|��@)�cw� 4@�$�<��!??J�V���@91���ٿ�|��@)�cw� 4@�$�<��!??J�V���@�Xѷ��ٿI�K��4�@Iβ8� 4@�����!?v�Q��a�@�Xѷ��ٿI�K��4�@Iβ8� 4@�����!?v�Q��a�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@xtQI�ٿ���@^W�ɺ4@�H����!?�|P��R�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@=O�"�ٿ�x��f��@��H2�4@9�q�!?$]x9�@W4�y��ٿ�Mz��s�@$G�4@�8����!?�,N�>�@W4�y��ٿ�Mz��s�@$G�4@�8����!?�,N�>�@W4�y��ٿ�Mz��s�@$G�4@�8����!?�,N�>�@W4�y��ٿ�Mz��s�@$G�4@�8����!?�,N�>�@W.�!(�ٿ	��ZD�@�a3X4@�%�'��!?ԲX�u�@W.�!(�ٿ	��ZD�@�a3X4@�%�'��!?ԲX�u�@W.�!(�ٿ	��ZD�@�a3X4@�%�'��!?ԲX�u�@�4(�ۆٿ6�9��@@�,��4@r�G���!?S�����@p�l�|�ٿ��n	9�@z�d�D4@��$��!?=�JH��@p�l�|�ٿ��n	9�@z�d�D4@��$��!?=�JH��@p�l�|�ٿ��n	9�@z�d�D4@��$��!?=�JH��@p�l�|�ٿ��n	9�@z�d�D4@��$��!?=�JH��@p�l�|�ٿ��n	9�@z�d�D4@��$��!?=�JH��@��Ք��ٿÿ=�S�@b	�$Z4@��8���!?���Ӏ�@��Ք��ٿÿ=�S�@b	�$Z4@��8���!?���Ӏ�@��Ք��ٿÿ=�S�@b	�$Z4@��8���!?���Ӏ�@��Ք��ٿÿ=�S�@b	�$Z4@��8���!?���Ӏ�@��Ք��ٿÿ=�S�@b	�$Z4@��8���!?���Ӏ�@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@�<1L�ٿE.D��@��!��3@��`�ސ!?�'�b���@��^	�ٿ�{��`��@��@�4@Ͳ����!?�gr��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@yT���ٿ�3��@��7؍4@����!?�+�؍��@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@������ٿ�Iߎ+�@��	4@�7u~y�!?����U"�@]��� �ٿ�֏���@�œ��4@D�P�!?)Oc5��@]��� �ٿ�֏���@�œ��4@D�P�!?)Oc5��@]��� �ٿ�֏���@�œ��4@D�P�!?)Oc5��@]��� �ٿ�֏���@�œ��4@D�P�!?)Oc5��@]��� �ٿ�֏���@�œ��4@D�P�!?)Oc5��@Tͭ���ٿn�����@�d^�4@��n�!?H�h���@Tͭ���ٿn�����@�d^�4@��n�!?H�h���@�ǘK��ٿ�n�k��@�Ȓ�4@9T���!?���˃��@�ǘK��ٿ�n�k��@�Ȓ�4@9T���!?���˃��@r�'�ٿqP�9��@&�X��4@�Ng^Ӑ!?�/ĕ�m�@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@���W��ٿ9-�-D�@��[�4@M�L�!?h�z��@3�|���ٿҵ����@Bl���4@7�<O@�!?	�ƟmY�@3�|���ٿҵ����@Bl���4@7�<O@�!?	�ƟmY�@3�|���ٿҵ����@Bl���4@7�<O@�!?	�ƟmY�@3�|���ٿҵ����@Bl���4@7�<O@�!?	�ƟmY�@3�|���ٿҵ����@Bl���4@7�<O@�!?	�ƟmY�@��O��ٿ�\�Th�@�O��?4@i�ş�!?�z)r;�@�Ҫ���ٿZ��e�H�@��ʻ�3@�Q��y�!?�%>����@��]�w�ٿ�lڳC�@�u0b�4@Vᎅ^�!?�.YH�@]3˷��ٿ�mC��@ܜ�64@�GL�!?j��[0��@]3˷��ٿ�mC��@ܜ�64@�GL�!?j��[0��@���ٿ���@EPNY�4@~���!?vx���@���ٿ���@EPNY�4@~���!?vx���@���ٿ���@EPNY�4@~���!?vx���@���ٿ���@EPNY�4@~���!?vx���@WV��ٿ��d6��@˿���4@	C]�M�!??.~���@�=V�}ٿ~Gf�g��@��f��4@���	�!?9!e���@�=V�}ٿ~Gf�g��@��f��4@���	�!?9!e���@�=V�}ٿ~Gf�g��@��f��4@���	�!?9!e���@�=V�}ٿ~Gf�g��@��f��4@���	�!?9!e���@�=V�}ٿ~Gf�g��@��f��4@���	�!?9!e���@ �ߠ$�ٿ�G��~b�@��UB�4@

���!?�ʗ^���@J,��ٿ��^�c�@0�d��4@��A��!? ~�+�@J,��ٿ��^�c�@0�d��4@��A��!? ~�+�@J,��ٿ��^�c�@0�d��4@��A��!? ~�+�@J,��ٿ��^�c�@0�d��4@��A��!? ~�+�@J,��ٿ��^�c�@0�d��4@��A��!? ~�+�@s�ۉ	�ٿ��Q}���@P�uz�4@)k0�ѐ!?-�X�M��@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@��x��ٿ��EwD�@�;��4@�
��ː!?mU`e
�@,�AJ�ٿL9Β �@���ŀ4@[��2��!?���O��@�>�)�~ٿ�ŪB���@J6| P4@G����!?/���Z]�@1��~ٿ�.+%��@QȘ��4@\ ���!?���S��@1��~ٿ�.+%��@QȘ��4@\ ���!?���S��@��濆ٿ��\!��@]��4@>����!?dl��U�@��濆ٿ��\!��@]��4@>����!?dl��U�@��濆ٿ��\!��@]��4@>����!?dl��U�@��濆ٿ��\!��@]��4@>����!?dl��U�@��濆ٿ��\!��@]��4@>����!?dl��U�@��濆ٿ��\!��@]��4@>����!?dl��U�@�s:�ٿ�Yk_���@`��4@Ex�!?=Y��H�@�s:�ٿ�Yk_���@`��4@Ex�!?=Y��H�@�s:�ٿ�Yk_���@`��4@Ex�!?=Y��H�@�&�1o�ٿvw�`���@$P$�p4@���ܐ!?J?q7��@�&�1o�ٿvw�`���@$P$�p4@���ܐ!?J?q7��@�}�#{ٿ�s�
	��@rc�Q4@9)}��!?�9Z�K�@�}�#{ٿ�s�
	��@rc�Q4@9)}��!?�9Z�K�@�}�#{ٿ�s�
	��@rc�Q4@9)}��!?�9Z�K�@�q>+�}ٿk��圙�@�w�b�4@��E���!?<\+F��@�q>+�}ٿk��圙�@�w�b�4@��E���!?<\+F��@�q>+�}ٿk��圙�@�w�b�4@��E���!?<\+F��@��&z{ٿq�w��f�@L�L�4@}�-��!?�:ܾ���@��ۖ�{ٿ*�ǚ,�@A�T�	4@ho�ŗ�!?:���@��ۖ�{ٿ*�ǚ,�@A�T�	4@ho�ŗ�!?:���@��ۖ�{ٿ*�ǚ,�@A�T�	4@ho�ŗ�!?:���@��ۖ�{ٿ*�ǚ,�@A�T�	4@ho�ŗ�!?:���@���;k{ٿ/�z9��@��ɏ4@��Mʦ�!?��
a$��@���;k{ٿ/�z9��@��ɏ4@��Mʦ�!?��
a$��@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@��\�~ٿ�̪#���@��-|Z4@�DU��!?�^�����@Wҙ�ٿ�9wh:�@�B�'; 4@Rcw0��!?9��J�<�@Wҙ�ٿ�9wh:�@�B�'; 4@Rcw0��!?9��J�<�@Wҙ�ٿ�9wh:�@�B�'; 4@Rcw0��!?9��J�<�@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@��旈ٿ�0縣�@�)��4@ܮ���!?�c����@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@l�	�ׇٿ�b>%΋�@�YB�4@A0'^ʐ!?�?1R�@���᪀ٿQi�q��@�C$
4@��er�!?4S`��@���᪀ٿQi�q��@�C$
4@��er�!?4S`��@���᪀ٿQi�q��@�C$
4@��er�!?4S`��@���᪀ٿQi�q��@�C$
4@��er�!?4S`��@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@ �f�ٿK2��E�@e�|�4@�.ތ��!?��K�@����ٿ^
�{)��@�lT�s4@T�:��!?p�BЇ�@��~�V�ٿ>�]���@�C7A�4@��W=�!?������@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@ӧ��[�ٿl�A�@���ؒ4@^�ʇ�!?l�?����@r=�,e�ٿC�נ��@�[�44@g���!?nz�|o��@r=�,e�ٿC�נ��@�[�44@g���!?nz�|o��@r=�,e�ٿC�נ��@�[�44@g���!?nz�|o��@r=�,e�ٿC�נ��@�[�44@g���!?nz�|o��@.��IՇٿ]������@��A�q4@/��R�!?gE�B��@.��IՇٿ]������@��A�q4@/��R�!?gE�B��@.��IՇٿ]������@��A�q4@/��R�!?gE�B��@.��IՇٿ]������@��A�q4@/��R�!?gE�B��@.��IՇٿ]������@��A�q4@/��R�!?gE�B��@��Cy)�ٿ�LO0���@�+6p�4@�0�a��!?�W�p��@��Cy)�ٿ�LO0���@�+6p�4@�0�a��!?�W�p��@��Cy)�ٿ�LO0���@�+6p�4@�0�a��!?�W�p��@P�"AI�ٿl�/��@��/��4@�M���!?Wep��/�@P�"AI�ٿl�/��@��/��4@�M���!?Wep��/�@t#1aT�ٿ���P�t�@��1�4@P�fy�!?ԫ��0�@�25��ٿ��O����@��M�a�3@?�?�l�!?>@����@�25��ٿ��O����@��M�a�3@?�?�l�!?>@����@��u�ٿ����@t�H�4@�����!?�O̘X�@��u�ٿ����@t�H�4@�����!?�O̘X�@��u�ٿ����@t�H�4@�����!?�O̘X�@��u�ٿ����@t�H�4@�����!?�O̘X�@<a�,ӈٿ��$����@v�s�4@"8ܠ�!?���c���@<a�,ӈٿ��$����@v�s�4@"8ܠ�!?���c���@<a�,ӈٿ��$����@v�s�4@"8ܠ�!?���c���@<a�,ӈٿ��$����@v�s�4@"8ܠ�!?���c���@<a�,ӈٿ��$����@v�s�4@"8ܠ�!?���c���@�Ұ�ֈٿ��-��@�]��4@'0їh�!?�(�2�%�@�Ұ�ֈٿ��-��@�]��4@'0їh�!?�(�2�%�@�$}ڇٿ6OQ��U�@��\�4@͏�N|�!?�>S�\�@�$}ڇٿ6OQ��U�@��\�4@͏�N|�!?�>S�\�@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@r2W$ҋٿ2M�����@�k�u4@�V�ߐ!?Z��=��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@c1#S��ٿ���C ��@���4@0�3��!?/XB{��@�R�s��ٿ]���s�@ę��4@\!7��!?��)��@�R�s��ٿ]���s�@ę��4@\!7��!?��)��@\�r�ٿ\�����@�^q�`4@6�$��!?�������@=�ꨂٿ� d\���@?�pz34@?Oz�ې!?O�O1��@�w	��}ٿ�Άl��@��aK4@�f�cא!?0Īw��@&�)�ٿ����%�@(���� 4@ M�!?�%�٪��@&�)�ٿ����%�@(���� 4@ M�!?�%�٪��@_E1�ٿiC�Qj��@�@6#4@��v�!?�
 ��z�@���Ìٿ���F���@�!�� 4@�a�m��!?�y�ۀJ�@���Ìٿ���F���@�!�� 4@�a�m��!?�y�ۀJ�@�Q�ٿ�Wr��@��9���3@0g�TȐ!??z�����@�}fڐٿu:���@����Q4@��a箐!?�z'w�a�@�}fڐٿu:���@����Q4@��a箐!?�z'w�a�@�}fڐٿu:���@����Q4@��a箐!?�z'w�a�@{Z'l�ٿ�O�2?�@�y�-K4@�{���!?�T�\Ǟ�@{Z'l�ٿ�O�2?�@�y�-K4@�{���!?�T�\Ǟ�@{Z'l�ٿ�O�2?�@�y�-K4@�{���!?�T�\Ǟ�@n��،ٿ��_�K+�@a���$4@�|��A�!?�M�$h��@.��B��ٿ.�=���@�QABx4@�/q)V�!?�qŶ��@.��B��ٿ.�=���@�QABx4@�/q)V�!?�qŶ��@.��B��ٿ.�=���@�QABx4@�/q)V�!?�qŶ��@.��B��ٿ.�=���@�QABx4@�/q)V�!?�qŶ��@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@��0T"�ٿ�c[s��@�F��4@廉ws�!?rId�Pl�@�̒$�ٿ�S'X5��@B5��4@^�$��!?��ϋ���@P����ٿ�Ջ��T�@:���4@��ҭ*�!?s�����@P����ٿ�Ջ��T�@:���4@��ҭ*�!?s�����@P����ٿ�Ջ��T�@:���4@��ҭ*�!?s�����@P����ٿ�Ջ��T�@:���4@��ҭ*�!?s�����@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@����ٿc'����@]'��4@3��#ߐ!?Y0���k�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@^����ٿ����W�@�M�7�4@�~ ��!?�@ ��^�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@M����ٿ0���O�@���p4@Pq�s�!?Z�X�l�@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@�%�<�ٿ��kd,�@�GP��4@h&TJ!?�������@/ѥ`�ٿ%���@3S�R�4@| �!?�c�X��@B9����ٿ��|�"��@�C~��4@.9؆ڐ!?�R����@B9����ٿ��|�"��@�C~��4@.9؆ڐ!?�R����@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@LD
��ٿ���@�'�@3G:bq4@Q�>��!?Í7TQ��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@Mź��ٿp��T� �@Fڄ4@� ���!?���6��@��V�ٿ�������@���1�4@c��@�!?eД<�U�@��V�ٿ�������@���1�4@c��@�!?eД<�U�@w5�5ňٿ%�	���@ƕۀ4@�0&2�!?�P�E�@w5�5ňٿ%�	���@ƕۀ4@�0&2�!?�P�E�@w5�5ňٿ%�	���@ƕۀ4@�0&2�!?�P�E�@w5�5ňٿ%�	���@ƕۀ4@�0&2�!?�P�E�@��a0�ٿ��~�g�@nd5'E 4@���9��!?���߰4�@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@��*��ٿ��*��t�@&oL�� 4@�e�
ؐ!? �k�M��@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ff;{e�ٿ�ІT�5�@φ�-4@��WА!?��^4N�@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@Ӡ���}ٿ�|����@�YL�4@��L���!?P&|���@[h��|�ٿ�$(ĐL�@L��T4@0N�Ȩ�!?���N��@�� ��ٿ���F �@�ʐz4@m��͐!?s	�K�@�� ��ٿ���F �@�ʐz4@m��͐!?s	�K�@�� ��ٿ���F �@�ʐz4@m��͐!?s	�K�@J���ٿ	t��'��@cts��4@��0���!?4.k�@J���ٿ	t��'��@cts��4@��0���!?4.k�@J���ٿ	t��'��@cts��4@��0���!?4.k�@J���ٿ	t��'��@cts��4@��0���!?4.k�@J���ٿ	t��'��@cts��4@��0���!?4.k�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@7�<Z�ٿ&��>6�@1|V��4@r��lڐ!?��iAp�@b��ԡ�ٿ�����J�@/GZ=�4@��]��!?Q6ʲ�@�,�O�ٿUqg�A�@��d��4@�Y�!?	qi �@�,�O�ٿUqg�A�@��d��4@�Y�!?	qi �@N"˙��ٿO�ב�2�@�DV^4@�:xΈ�!?I�D�r��@N"˙��ٿO�ב�2�@�DV^4@�:xΈ�!?I�D�r��@N"˙��ٿO�ב�2�@�DV^4@�:xΈ�!?I�D�r��@6֤� �ٿ�C2��@J{J4@V!6Ɛ!?d����@6֤� �ٿ�C2��@J{J4@V!6Ɛ!?d����@6֤� �ٿ�C2��@J{J4@V!6Ɛ!?d����@��c�A�ٿ^�'f��@!�.24@�����!?�o���@��c�A�ٿ^�'f��@!�.24@�����!?�o���@��c�A�ٿ^�'f��@!�.24@�����!?�o���@��c�A�ٿ^�'f��@!�.24@�����!?�o���@��c�A�ٿ^�'f��@!�.24@�����!?�o���@��c�A�ٿ^�'f��@!�.24@�����!?�o���@�/�oN�ٿ�H-�[�@`��4@P����!?u�;���@�/�oN�ٿ�H-�[�@`��4@P����!?u�;���@�/�oN�ٿ�H-�[�@`��4@P����!?u�;���@���j�ٿB �`E%�@���4@�e��!?�֙�6|�@��<�-~ٿsE�ת�@��BJ4@������!?X�	Ɔ�@��<�-~ٿsE�ת�@��BJ4@������!?X�	Ɔ�@��<�-~ٿsE�ת�@��BJ4@������!?X�	Ɔ�@��<�-~ٿsE�ת�@��BJ4@������!?X�	Ɔ�@��<�-~ٿsE�ת�@��BJ4@������!?X�	Ɔ�@���ٿ|!�Fy1�@��%��4@��k�!?e�T���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@;�žK�ٿ:���X�@��U��4@��K��!?��"m���@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@�vܿ~ٿ�x�h���@C��	4@��a4ѐ!?l(�{�@���-~ٿ_��\Q��@.�p�
4@��Y���!?t��	�d�@���N�ٿ�\]2�@5S{�T4@��H��!?lCE�c�@���N�ٿ�\]2�@5S{�T4@��H��!?lCE�c�@,|>�ٿ�&����@��뒢4@�	y��!?Qj��:m�@f�1��ٿ��YU���@9�.b�	4@�67�!?��?��0�@f�1��ٿ��YU���@9�.b�	4@�67�!?��?��0�@f�1��ٿ��YU���@9�.b�	4@�67�!?��?��0�@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�qpZ1�ٿ�I�K0�@���X�4@(j�hǐ!?��

���@�to	�ٿ(���	6�@�?�Ȧ4@Ce;&��!?�s||�H�@�to	�ٿ(���	6�@�?�Ȧ4@Ce;&��!?�s||�H�@���ˏٿ��X��@�?���4@TO ���!?�%G���@���ˏٿ��X��@�?���4@TO ���!?�%G���@���ˏٿ��X��@�?���4@TO ���!?�%G���@��>�ٿ��(���@���%4@l�͐!?]��I6��@��ĉٿ�	6/ߵ�@���\�4@>�?�!?~�����@��ĉٿ�	6/ߵ�@���\�4@>�?�!?~�����@��ĉٿ�	6/ߵ�@���\�4@>�?�!?~�����@q�Q3k�ٿ\TB�,�@Ϡ4@�����!?�M-��@q�Q3k�ٿ\TB�,�@Ϡ4@�����!?�M-��@q�Q3k�ٿ\TB�,�@Ϡ4@�����!?�M-��@q�Q3k�ٿ\TB�,�@Ϡ4@�����!?�M-��@q�Q3k�ٿ\TB�,�@Ϡ4@�����!?�M-��@E��~ٿ̪�0�@��E�4@{�
�!?�� '��@E��~ٿ̪�0�@��E�4@{�
�!?�� '��@E��~ٿ̪�0�@��E�4@{�
�!?�� '��@EQ+��ٿ�����@s�
� 4@�Q�ː!?�?9�@EQ+��ٿ�����@s�
� 4@�Q�ː!?�?9�@EQ+��ٿ�����@s�
� 4@�Q�ː!?�?9�@EQ+��ٿ�����@s�
� 4@�Q�ː!?�?9�@EQ+��ٿ�����@s�
� 4@�Q�ː!?�?9�@�m��*�ٿ����"�@Fn��Z 4@��o��!?�X���j�@�m��*�ٿ����"�@Fn��Z 4@��o��!?�X���j�@�m��*�ٿ����"�@Fn��Z 4@��o��!?�X���j�@�N|1Txٿ��B��@�pxQ
4@�˲��!?�t'��@�N|1Txٿ��B��@�pxQ
4@�˲��!?�t'��@�N|1Txٿ��B��@�pxQ
4@�˲��!?�t'��@x¡<ւٿ��ǔi[�@���)�3@H�~Z�!?#B1C��@x¡<ւٿ��ǔi[�@���)�3@H�~Z�!?#B1C��@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�{�ٿ�}ǳ�m�@�;@Hy4@�v�!?JBA�h�@�N��ٿH�w�]!�@X�l�4@	�]!�!?G8�&=�@��:|�ٿ�a=U��@�8��4@gn򢲐!?[Լ�NG�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@	��y�ٿǏ	eK�@��� 4@�rϜ�!?̫��b�@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�岓E�ٿǘ0V���@&��
^4@�.�E�!?��;���@�6	��ٿ?;�%��@Յ=�� 4@��� �!?�UDV��@�6	��ٿ?;�%��@Յ=�� 4@��� �!?�UDV��@�6	��ٿ?;�%��@Յ=�� 4@��� �!?�UDV��@��>� �ٿ��qKl}�@�2k@4@�;���!?Ko�"s}�@��>� �ٿ��qKl}�@�2k@4@�;���!?Ko�"s}�@��>� �ٿ��qKl}�@�2k@4@�;���!?Ko�"s}�@��>� �ٿ��qKl}�@�2k@4@�;���!?Ko�"s}�@�u����ٿ��6���@~�떔4@QbA[��!?";߳���@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@���bцٿ��
SD�@�� l44@q�I���!?p3I��|�@M���ٿM��
��@�bq��4@R�,��!?R:x��L�@M���ٿM��
��@�bq��4@R�,��!?R:x��L�@�~ٿ�֗R�@��R�4@ Cݺ�!?��͕5��@�~ٿ�֗R�@��R�4@ Cݺ�!?��͕5��@JG�'��ٿ{%�2��@w�=L�4@>�.Ő!?9��d��@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@,�t!)�ٿ
S��D��@
�� 
4@��l��!?z[x���@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@��cSq�ٿ��0=8��@�]Q��4@�<ZQ��!?�7I"/�@9�ٿ#�<m~��@�$e?�4@O�૾�!?���72i�@�f��8ٿ�A���@^��4@Պ�o�!?��	,�@�f��8ٿ�A���@^��4@Պ�o�!?��	,�@�f��8ٿ�A���@^��4@Պ�o�!?��	,�@�f��8ٿ�A���@^��4@Պ�o�!?��	,�@��V0~ٿIY�#��@���NC4@����~�!?b��_��@��V0~ٿIY�#��@���NC4@����~�!?b��_��@��V0~ٿIY�#��@���NC4@����~�!?b��_��@L����ٿ�X~���@*�X�e4@F�K���!?^�g9�a�@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@�}p�"�ٿ5��at�@��~�)4@$�&�א!?0�д��@pc�{ٿ�>냬��@�!?�4@P�c��!? �i/���@Y����ٿ��wK�@�ҩ�;4@#;BlҐ!?�&o�G��@Y����ٿ��wK�@�ҩ�;4@#;BlҐ!?�&o�G��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@�{��)�ٿ �6C��@��k�=4@�,f拐!?��}��@���_�ٿb���f/�@�V$��4@<]]4��!?�[��@���_�ٿb���f/�@�V$��4@<]]4��!?�[��@���_�ٿb���f/�@�V$��4@<]]4��!?�[��@���0�ٿ���F66�@!���4@��T��!?����':�@���0�ٿ���F66�@!���4@��T��!?����':�@���0�ٿ���F66�@!���4@��T��!?����':�@���3�ٿ���4	��@.�A�4@Hٹ�!?�Y�B��@�L$�~�ٿQ�F���@EYti@4@�6ejא!?�HuQ6��@w[MKٿLM��Q�@�[�n�4@s�C��!?:�PqS�@w[MKٿLM��Q�@�[�n�4@s�C��!?:�PqS�@w[MKٿLM��Q�@�[�n�4@s�C��!?:�PqS�@w[MKٿLM��Q�@�[�n�4@s�C��!?:�PqS�@w[MKٿLM��Q�@�[�n�4@s�C��!?:�PqS�@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@�i"�ٿ��9���@t�|{}4@�t�Ȑ!?��}q��@���m�ٿTA?Ѭ�@��I4@U��̐!?8L�;N��@���m�ٿTA?Ѭ�@��I4@U��̐!?8L�;N��@���m�ٿTA?Ѭ�@��I4@U��̐!?8L�;N��@���m�ٿTA?Ѭ�@��I4@U��̐!?8L�;N��@���m�ٿTA?Ѭ�@��I4@U��̐!?8L�;N��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@�;���ٿES]���@��� 4@�x/�ː!?�IÂ��@2aX�&�ٿ�ze���@{��<4@@Xi��!?K�x�@2aX�&�ٿ�ze���@{��<4@@Xi��!?K�x�@2aX�&�ٿ�ze���@{��<4@@Xi��!?K�x�@2aX�&�ٿ�ze���@{��<4@@Xi��!?K�x�@���iS�ٿ�^���@�zt�4@�3�u��!?�dv�]E�@���iS�ٿ�^���@�zt�4@�3�u��!?�dv�]E�@�K`��ٿYA�=5r�@�s� 4@�bP��!?�,F�X�@�K`��ٿYA�=5r�@�s� 4@�bP��!?�,F�X�@�&����ٿ�*c�)�@"H1� 4@=|D���!?}�Lk���@�&����ٿ�*c�)�@"H1� 4@=|D���!?}�Lk���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@́��Ðٿ�(�-4�@��1�4@p�z}ܐ!?�TM]���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@'����ٿA��k��@�;��4@��wZ�!?�9���@;��AN�ٿ����&�@t��}44@� �V�!?�Wq����@�7�u�ٿ�T��@���� 4@�3��!?�U0���@l�
�!�ٿ%;���@SY.�4@��-"�!?e /���@l�
�!�ٿ%;���@SY.�4@��-"�!?e /���@/9v���ٿCm���@Ķ4@i�T��!?��	q��@/9v���ٿCm���@Ķ4@i�T��!?��	q��@/9v���ٿCm���@Ķ4@i�T��!?��	q��@/9v���ٿCm���@Ķ4@i�T��!?��	q��@/9v���ٿCm���@Ķ4@i�T��!?��	q��@�b1�ٿ���JE��@���#J4@?�?��!?mؠ\���@�(ɻ�ٿ7r�@�@�~��4@��x�"�!?�Z�Q��@�(ɻ�ٿ7r�@�@�~��4@��x�"�!?�Z�Q��@�(ɻ�ٿ7r�@�@�~��4@��x�"�!?�Z�Q��@�(ɻ�ٿ7r�@�@�~��4@��x�"�!?�Z�Q��@^�B���ٿ�NT�]��@TsB-�4@�%noa�!?)�~$�@^�B���ٿ�NT�]��@TsB-�4@�%noa�!?)�~$�@?�k��ٿ*�q`��@�ET�3@=���!�!?k�Cܼ�@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@�����ٿ� f�r=�@�=s'�3@�R��!?�6�1��@?����ٿ��/�`��@#m!!Q 4@�^��E�!?�J�+W>�@?����ٿ��/�`��@#m!!Q 4@�^��E�!?�J�+W>�@?����ٿ��/�`��@#m!!Q 4@�^��E�!?�J�+W>�@���m�ٿ0��ai��@�e��84@���'�!?^��hz�@���m�ٿ0��ai��@�e��84@���'�!?^��hz�@�T���ٿEM�����@ؾ|�14@�%B>^�!?Ӣ����@'D��R�ٿԢm���@�o��t4@h��(�!?(�	9��@����ٿX� �V<�@��v^4@��``�!?/^���@����ٿX� �V<�@��v^4@��``�!?/^���@����ٿX� �V<�@��v^4@��``�!?/^���@jٿ���$x��@o�+d� 4@V2& ��!?�_Ǡ�`�@jٿ���$x��@o�+d� 4@V2& ��!?�_Ǡ�`�@jٿ���$x��@o�+d� 4@V2& ��!?�_Ǡ�`�@x����ٿ�`����@#gд4@��%��!?�(�S|�@ȅ[�ӈٿe�-Z��@t{e >�3@���lt�!?�M�ij��@ȅ[�ӈٿe�-Z��@t{e >�3@���lt�!?�M�ij��@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@�����ٿ�;8����@H��3@�{*���!?���s�s�@��A��ٿ�+q�|*�@@̲�)4@8R�d��!?��&3���@��A��ٿ�+q�|*�@@̲�)4@8R�d��!?��&3���@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�B_�ٿ��mt���@�4@4@a���!?6Q�GR��@�"j}�ٿ��8$���@m�v�4@�w�ڰ�!?>�U2�@�"j}�ٿ��8$���@m�v�4@�w�ڰ�!?>�U2�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�P��ڊٿϫ���@�K+4@)�P���!?P-�!tO�@�I�<�ٿRazc��@����s4@���!?�=��:q�@�I�<�ٿRazc��@����s4@���!?�=��:q�@�I�<�ٿRazc��@����s4@���!?�=��:q�@�I�<�ٿRazc��@����s4@���!?�=��:q�@�I�<�ٿRazc��@����s4@���!?�=��:q�@$�
�ٿ�E�M;��@�e�/ 4@�,����!?�a��i�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@Њ&��ٿaSn��^�@�
19 4@~a��ܐ!?/��Z�@���]Ћٿ�%9�!C�@���*�4@�q����!?���V�@���]Ћٿ�%9�!C�@���*�4@�q����!?���V�@���]Ћٿ�%9�!C�@���*�4@�q����!?���V�@���]Ћٿ�%9�!C�@���*�4@�q����!?���V�@���]Ћٿ�%9�!C�@���*�4@�q����!?���V�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@��<�ٿ'���o��@���گ4@��ʐ!?e!ѧW�@K&�ٿsa���@�8��4@�p��!?���fZ�@K&�ٿsa���@�8��4@�p��!?���fZ�@K&�ٿsa���@�8��4@�p��!?���fZ�@���ח�ٿ���\M�@�3���4@S�����!?�vQu�@���ח�ٿ���\M�@�3���4@S�����!?�vQu�@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@D˔E�ٿb�
��)�@(���4@�y �!?�3��@��>�ٿ�&Q�<�@��O4@;�%���!?tj]��@��>�ٿ�&Q�<�@��O4@;�%���!?tj]��@��>�ٿ�&Q�<�@��O4@;�%���!?tj]��@��>�ٿ�&Q�<�@��O4@;�%���!?tj]��@��>�ٿ�&Q�<�@��O4@;�%���!?tj]��@�����ٿ���w���@�ֳD�4@���}e�!?��*=���@�����ٿ���w���@�ֳD�4@���}e�!?��*=���@�����ٿ���w���@�ֳD�4@���}e�!?��*=���@�����ٿ���w���@�ֳD�4@���}e�!?��*=���@�����ٿ���w���@�ֳD�4@���}e�!?��*=���@$L֊�ٿ��s&Ӗ�@���K@4@������!?��%����@$L֊�ٿ��s&Ӗ�@���K@4@������!?��%����@��q��ٿ��.�&�@���4@z����!?�R��F�@��q��ٿ��.�&�@���4@z����!?�R��F�@��q��ٿ��.�&�@���4@z����!?�R��F�@��q��ٿ��.�&�@���4@z����!?�R��F�@�c��ٿ�����@* %R4@H����!?�74|�@�c��ٿ�����@* %R4@H����!?�74|�@�c��ٿ�����@* %R4@H����!?�74|�@�c��ٿ�����@* %R4@H����!?�74|�@��^�ʂٿ�rqb��@ؗ4@+c���!?̻���@��^�ʂٿ�rqb��@ؗ4@+c���!?̻���@��^�ʂٿ�rqb��@ؗ4@+c���!?̻���@��^�ʂٿ�rqb��@ؗ4@+c���!?̻���@��^�ʂٿ�rqb��@ؗ4@+c���!?̻���@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@����ٿ���d��@��|��4@C�w��!?��K'�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@kG��{ٿ�Ni���@�"�B4@�%�	�!?�"<^�@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@#S^0�ٿ$���޶�@X'��4@&k��Ր!?�����@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@
�'E8�ٿ�F����@�S�C4@�dI8͐!?�t��i;�@n�m�'�ٿ�f �=��@(��|�4@|�Q���!?���I�G�@��>	�ٿ5o ��@`�ח�4@<|����!?c�Vj��@��>	�ٿ5o ��@`�ח�4@<|����!?c�Vj��@��>	�ٿ5o ��@`�ח�4@<|����!?c�Vj��@��>	�ٿ5o ��@`�ח�4@<|����!?c�Vj��@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�XC�߁ٿ��,���@�t�4@������!?��%(݆�@�v.��ٿUN.I:p�@���]4@Jp�!?�윻'�@Z�S�B�ٿ]� �-�@ ����4@��a�|�!?6��;��@Z�S�B�ٿ]� �-�@ ����4@��a�|�!?6��;��@Z�S�B�ٿ]� �-�@ ����4@��a�|�!?6��;��@Y/��ٿ |�5��@��Q�4@gm��\�!?��ۖf�@Y/��ٿ |�5��@��Q�4@gm��\�!?��ۖf�@Y/��ٿ |�5��@��Q�4@gm��\�!?��ۖf�@���0~ٿ�y�<٨�@�f��4@�6����!?̾��T�@���0~ٿ�y�<٨�@�f��4@�6����!?̾��T�@���Eԃٿ�GΑ��@������3@�jo6��!?Ɗ����@���Eԃٿ�GΑ��@������3@�jo6��!?Ɗ����@x�߿�ٿ�e�D�&�@�9�X4@�8��ϐ!?����@x�߿�ٿ�e�D�&�@�9�X4@�8��ϐ!?����@x�߿�ٿ�e�D�&�@�9�X4@�8��ϐ!?����@x�߿�ٿ�e�D�&�@�9�X4@�8��ϐ!?����@��W��ٿ]��U �@��I�4@��w���!?�f�k�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@k[����ٿ:FoH�@�@ WxmG4@��A��!?ͯ�7�c�@W]��ٿ'GL�M�@p#4�4@��
+�!?E��,��@��ps�ٿ��Ũ��@ha�K� 4@����!?:�w��
�@��ps�ٿ��Ũ��@ha�K� 4@����!?:�w��
�@��ps�ٿ��Ũ��@ha�K� 4@����!?:�w��
�@6��2>�ٿ����@��@�4@�Y���!?!�C�t�@6��2>�ٿ����@��@�4@�Y���!?!�C�t�@6��2>�ٿ����@��@�4@�Y���!?!�C�t�@6��2>�ٿ����@��@�4@�Y���!?!�C�t�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@������ٿ�����{�@��P<4@���ju�!?�s��V�@��t��ٿH�H�� �@�RBM 4@2��p��!?Y��֙�@��t��ٿH�H�� �@�RBM 4@2��p��!?Y��֙�@��t��ٿH�H�� �@�RBM 4@2��p��!?Y��֙�@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�Ol�&�ٿJ�?��@H�\t�3@x^Ԑ!?���L��@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@�G)�ٿ�6��1��@���G4@<)~!!�!?$�Ý�!�@G���ٿ2g+���@�����4@z�ǒ�!?ѥ�Q�M�@G���ٿ2g+���@�����4@z�ǒ�!?ѥ�Q�M�@���}ٿ ��q���@\���4@�&�ې!?�(�x�@7�D��ٿ��p����@��r�4@	)�3�!?���@7�D��ٿ��p����@��r�4@	)�3�!?���@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�St��ٿ�n ���@�r�9R4@�lz��!?`��t"��@�Mt]�ٿ�B�V~�@H7��� 4@g��t�!?���Pb9�@�Mt]�ٿ�B�V~�@H7��� 4@g��t�!?���Pb9�@�Mt]�ٿ�B�V~�@H7��� 4@g��t�!?���Pb9�@�Mt]�ٿ�B�V~�@H7��� 4@g��t�!?���Pb9�@�Mt]�ٿ�B�V~�@H7��� 4@g��t�!?���Pb9�@�B�K�ٿb�j���@v�=4@�M;��!?�� ���@��W�1�ٿD��{C�@b��3@f��ې!?]�uւ�@�G��ٿ����mq�@ � ��3@�ٔ�Ӑ!?b�����@�G��ٿ����mq�@ � ��3@�ٔ�Ӑ!?b�����@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@w@J�ٿ�9�w���@Z��2 4@��ˀ�!?zR��'�@�sc��ٿcC�� ��@*��,�4@�&w�!?��7?!�@�sc��ٿcC�� ��@*��,�4@�&w�!?��7?!�@�sc��ٿcC�� ��@*��,�4@�&w�!?��7?!�@�sc��ٿcC�� ��@*��,�4@�&w�!?��7?!�@��G�ٿ����#��@���� 4@3c<��!?pK��k�@^�!_�ٿ��Y����@�s�f4@�9	���!?i�I�u��@���ٿ�����P�@rKo�24@T��`�!?�D��Y�@�V�e|ٿ����� �@A��4@����Ð!?�uXZ���@^[��zٿ�9���@� �4@a�#0��!?��{s,�@^[��zٿ�9���@� �4@a�#0��!?��{s,�@餬~ٿJ'Y��@3#��W4@���}r�!?7��9�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@\�xI��ٿL��h��@<�
��4@�)?�w�!?�+-&�@�ȭ�V�ٿ��=�V5�@�V�`�4@�5o��!?ʓA�^�@�ȭ�V�ٿ��=�V5�@�V�`�4@�5o��!?ʓA�^�@�ȭ�V�ٿ��=�V5�@�V�`�4@�5o��!?ʓA�^�@�ȭ�V�ٿ��=�V5�@�V�`�4@�5o��!?ʓA�^�@�ȭ�V�ٿ��=�V5�@�V�`�4@�5o��!?ʓA�^�@͈)�܁ٿ�eՋ-t�@Όہw4@���hؐ!?��yo�A�@͈)�܁ٿ�eՋ-t�@Όہw4@���hؐ!?��yo�A�@͈)�܁ٿ�eՋ-t�@Όہw4@���hؐ!?��yo�A�@��v́ٿuީ����@� /�4@�٧�!?���1�'�@��v́ٿuީ����@� /�4@�٧�!?���1�'�@��v́ٿuީ����@� /�4@�٧�!?���1�'�@��v́ٿuީ����@� /�4@�٧�!?���1�'�@��v́ٿuީ����@� /�4@�٧�!?���1�'�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@ �~|��ٿ��!X��@@���4@�J�O��!?^Ҫ��~�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@��}���ٿ�������@�H�e\ 4@���o!?�Êp0�@|҂Y��ٿ��K���@-�Y�4@��HƳ�!?�MC�-�@�M:�|ٿ,�����@z����4@��%��!?GM0����@�M:�|ٿ,�����@z����4@��%��!?GM0����@A���zٿ&�n`���@��y�4@b�����!?����V�@7Q
��zٿ��{ZYI�@E��T4@K#hƐ!?���^tm�@jc$H�ٿ��ķ���@_�.9G4@�U�p�!?��^��G�@jc$H�ٿ��ķ���@_�.9G4@�U�p�!?��^��G�@jc$H�ٿ��ķ���@_�.9G4@�U�p�!?��^��G�@�/�{}ٿ��H�-I�@�� �44@L���!?�]�����@��F�!|ٿN�\mh��@�y	 4@�}���!?����I��@��F�!|ٿN�\mh��@�y	 4@�}���!?����I��@��F�!|ٿN�\mh��@�y	 4@�}���!?����I��@��F�!|ٿN�\mh��@�y	 4@�}���!?����I��@�`�zٿ�FB��@H�N�4@�m����!?�h���@�`�zٿ�FB��@H�N�4@�m����!?�h���@�`�zٿ�FB��@H�N�4@�m����!?�h���@�`�zٿ�FB��@H�N�4@�m����!?�h���@�`�zٿ�FB��@H�N�4@�m����!?�h���@����zٿT �4��@;�u5e4@&���!?Y/����@q�2_>ٿE`����@;:��4@�lP�!?��fB͒�@q�2_>ٿE`����@;:��4@�lP�!?��fB͒�@q�2_>ٿE`����@;:��4@�lP�!?��fB͒�@q�2_>ٿE`����@;:��4@�lP�!?��fB͒�@q�2_>ٿE`����@;:��4@�lP�!?��fB͒�@�x]�ٿHp��#�@ک�;4@'�`��!?�7͵���@�x]�ٿHp��#�@ک�;4@'�`��!?�7͵���@���ٿ9����@ǩ+ɽ4@�ε�!?�݈o��@���ٿ9����@ǩ+ɽ4@�ε�!?�݈o��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@"��#�ٿ*���*�@��@4@íJK �!?�HG>Y��@w���ٿ��?"��@�kIo� 4@�{�ː!?��ܰ�@[��Q�ٿ� �:���@M��JP�3@̎��m�!?�MO� ��@[��Q�ٿ� �:���@M��JP�3@̎��m�!?�MO� ��@[��Q�ٿ� �:���@M��JP�3@̎��m�!?�MO� ��@[��Q�ٿ� �:���@M��JP�3@̎��m�!?�MO� ��@[��Q�ٿ� �:���@M��JP�3@̎��m�!?�MO� ��@9$���ٿN��&��@)	 n;4@呖!��!?��L�.�@9$���ٿN��&��@)	 n;4@呖!��!?��L�.�@��`"�ٿF\�xG��@u��O�4@ Lk`�!?������@��`"�ٿF\�xG��@u��O�4@ Lk`�!?������@��Zh�ٿo�'��Z�@�Wti�	4@-�;�!?��RL]�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@/'R�΅ٿ��Z�v�@;^��]4@U,��!?�ݺ��v�@�5�B�ٿC*��9�@+�3#<4@�=m�(�!?Ǉ��F��@�5�B�ٿC*��9�@+�3#<4@�=m�(�!?Ǉ��F��@�5�B�ٿC*��9�@+�3#<4@�=m�(�!?Ǉ��F��@�5�B�ٿC*��9�@+�3#<4@�=m�(�!?Ǉ��F��@r����ٿ���d�@�&��4@��B�Ӑ!?�Ų6D��@r����ٿ���d�@�&��4@��B�Ӑ!?�Ų6D��@r����ٿ���d�@�&��4@��B�Ӑ!?�Ų6D��@r����ٿ���d�@�&��4@��B�Ӑ!?�Ų6D��@�@x�ٿY�K�VR�@
1ğ�4@.*tD��!?�]2�V�@�@x�ٿY�K�VR�@
1ğ�4@.*tD��!?�]2�V�@�@x�ٿY�K�VR�@
1ğ�4@.*tD��!?�]2�V�@�@x�ٿY�K�VR�@
1ğ�4@.*tD��!?�]2�V�@`�U�o�ٿ��awn�@�㈨4@�+L��!?�S�r��@`�U�o�ٿ��awn�@�㈨4@�+L��!?�S�r��@`�U�o�ٿ��awn�@�㈨4@�+L��!?�S�r��@`�U�o�ٿ��awn�@�㈨4@�+L��!?�S�r��@0�N/ۉٿ�ؿ^��@���F�4@�v;��!? �n��!�@0�N/ۉٿ�ؿ^��@���F�4@�v;��!? �n��!�@0�N/ۉٿ�ؿ^��@���F�4@�v;��!? �n��!�@�$���}ٿ�$���@�O� 4@�Ṅ�!?ӻ=j���@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@k���}ٿK�?�m��@��7�4@�E{�Ր!?'%�s)��@��1�ٿ�V7.���@s�k�4@ti|���!?�s����@��1�ٿ�V7.���@s�k�4@ti|���!?�s����@��1�ٿ�V7.���@s�k�4@ti|���!?�s����@�x��ٿ�o�o���@g�+U4@�h��!?��H�y�@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@:�k�Y�ٿ�����@MVw�4@���ǐ!?�tR4P��@98�5��ٿ�b0oN��@�7�4@'H�Ͷ�!?u~_��@98�5��ٿ�b0oN��@�7�4@'H�Ͷ�!?u~_��@98�5��ٿ�b0oN��@�7�4@'H�Ͷ�!?u~_��@���;s�ٿϧ��pr�@���P4@�?f[��!?�&�!y��@���;s�ٿϧ��pr�@���P4@�?f[��!?�&�!y��@���;s�ٿϧ��pr�@���P4@�?f[��!?�&�!y��@���;s�ٿϧ��pr�@���P4@�?f[��!?�&�!y��@�'{T��ٿ���K�@N���c4@�Vx~�!?2U\3���@�'{T��ٿ���K�@N���c4@�Vx~�!?2U\3���@�'{T��ٿ���K�@N���c4@�Vx~�!?2U\3���@�'{T��ٿ���K�@N���c4@�Vx~�!?2U\3���@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�+В��ٿܾ�Ѭa�@d���4@;�� -�!?:�ͻ6��@�%�v�ٿdDo�|�@e��q4@�A��!?���#��@��i�ٿ�-��۴�@bxx�4@���뻐!?	����@��i�ٿ�-��۴�@bxx�4@���뻐!?	����@��i�ٿ�-��۴�@bxx�4@���뻐!?	����@f��D�ٿ�$�)r�@�ML	:4@��:��!?�M��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@��yc�ٿBi�7{�@bq��R 4@�� ��!?��f��@����ٿ2'�s�N�@&�X���3@�����!?�I�/n��@�oSџ�ٿ�NS˫�@�����3@�� ��!?��9��W�@�oSџ�ٿ�NS˫�@�����3@�� ��!?��9��W�@6���ٿb�+}�@ۆ��4@��Լʐ!?y&�6��@nAؑ�ٿB�5R�z�@��L��4@d�1W��!?u<'�C��@����s�ٿ������@(�	��4@�|^|��!?��xJd�@����s�ٿ������@(�	��4@�|^|��!?��xJd�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@F�g �ٿa�)͙n�@ژ�
#4@ݡ�ﺐ!?]��݈�@~]ٝ��ٿ*��Ơ�@n��� 4@�ʝ���!?
wl��@~]ٝ��ٿ*��Ơ�@n��� 4@�ʝ���!?
wl��@~]ٝ��ٿ*��Ơ�@n��� 4@�ʝ���!?
wl��@��S�~ٿ��Ŭ�@u���4@FT�T��!?.�!�p�@��S�~ٿ��Ŭ�@u���4@FT�T��!?.�!�p�@��S�~ٿ��Ŭ�@u���4@FT�T��!?.�!�p�@��S�~ٿ��Ŭ�@u���4@FT�T��!?.�!�p�@��S�~ٿ��Ŭ�@u���4@FT�T��!?.�!�p�@�ݵ���ٿ��4 ��@�%��4@��>��!?�uN��e�@�ݵ���ٿ��4 ��@�%��4@��>��!?�uN��e�@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@����Z�ٿ��NM���@'���:4@D���!?dA��"��@W<�Q�ٿȅRT[�@M����4@Y!��ݐ!?\��zb�@���lZ�ٿ����@jx� 4@���"�!?��]��X�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@� ���ٿ�E��!��@|���4@���"�!?D�X�5�@
�'���ٿi�r�b�@:rVz#4@8�ὐ!?b�s�Փ�@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@���47�ٿ̉��/�@9O���4@�f~J��!?�[տs��@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@ ��o�ٿ=9��|@�@��,��4@�rV6��!?-AE�!�@�4Ì��ٿRh'�3e�@Ӆ p
4@.1�v�!?Q��T_�@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�3����ٿR�P�0��@�U4@��3�Ր!?�r3���@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�/��W�ٿ�1����@��\;�
4@��|Ґ!?��o[�@�s;�ٿ����l�@��"�4@F$sT��!?q��P�@�s;�ٿ����l�@��"�4@F$sT��!?q��P�@�s;�ٿ����l�@��"�4@F$sT��!?q��P�@�s;�ٿ����l�@��"�4@F$sT��!?q��P�@�s;�ٿ����l�@��"�4@F$sT��!?q��P�@,m�k5�ٿz��.$��@�=�	4@��l���!?�7�-j�@,m�k5�ٿz��.$��@�=�	4@��l���!?�7�-j�@,m�k5�ٿz��.$��@�=�	4@��l���!?�7�-j�@,m�k5�ٿz��.$��@�=�	4@��l���!?�7�-j�@,m�k5�ٿz��.$��@�=�	4@��l���!?�7�-j�@Aa�ٿ��Ws��@CPp�.4@^���!?�><���@Aa�ٿ��Ws��@CPp�.4@^���!?�><���@Aa�ٿ��Ws��@CPp�.4@^���!?�><���@Aa�ٿ��Ws��@CPp�.4@^���!?�><���@Aa�ٿ��Ws��@CPp�.4@^���!?�><���@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@G�&rޅٿ��,6V�@�\<t�4@3�h��!?�kBOk�@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@p5.Âٿ���l�@6X��4@���)Ɛ!?�i}��@�g���ٿ��Rg��@Tj_R4@㼋�!?
2����@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@D�?��ٿ�<�Ѝ��@����4@�}��!?A4��}�@�PpІٿ�O�`���@_t�4@����!?�II�@�PpІٿ�O�`���@_t�4@����!?�II�@�PpІٿ�O�`���@_t�4@����!?�II�@J@�i�ٿ�+�ӯh�@��eW4@.֫��!?�S�Ŀ�@J@�i�ٿ�+�ӯh�@��eW4@.֫��!?�S�Ŀ�@J@�i�ٿ�+�ӯh�@��eW4@.֫��!?�S�Ŀ�@J@�i�ٿ�+�ӯh�@��eW4@.֫��!?�S�Ŀ�@x�5��ٿ��jl8�@yr��4@���̐!?��)r|��@x�5��ٿ��jl8�@yr��4@���̐!?��)r|��@x�5��ٿ��jl8�@yr��4@���̐!?��)r|��@x�5��ٿ��jl8�@yr��4@���̐!?��)r|��@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@	1Z྄ٿ���Ҷ�@9��4@������!?��q"���@�B'=�ٿ���ҽ3�@"(vD4@t*:Q��!?�h�m��@�Ų��ٿG��4�"�@ǵ%3)4@�_�\1�!?�35�q�@�Ų��ٿG��4�"�@ǵ%3)4@�_�\1�!?�35�q�@�Ų��ٿG��4�"�@ǵ%3)4@�_�\1�!?�35�q�@�Ų��ٿG��4�"�@ǵ%3)4@�_�\1�!?�35�q�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@`��ٿ�6����@ -6��4@9N�	�!?�7T�_�@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@;h����ٿ�"h{ښ�@v�O#4@ެ=:�!?X�r���@T4Ӽ��ٿ���M?�@9\`n�4@����!?�����@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@?�!�ٿ��j7S�@J���4@|j��א!?�#2�F��@�9�$�ٿ0Ԭ]��@�����3@�ק���!?P�s��@�9�$�ٿ0Ԭ]��@�����3@�ק���!?P�s��@�9�$�ٿ0Ԭ]��@�����3@�ק���!?P�s��@��H�!�ٿS[��Q��@��L��3@v�,O�!?�gB��@��H�!�ٿS[��Q��@��L��3@v�,O�!?�gB��@��H�!�ٿS[��Q��@��L��3@v�,O�!?�gB��@g���ٿ6	�+a��@��`�'4@;�1�T�!?`�h���@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@�6`��ٿ�d1��@z���4@w�C�!?�~Fn\�@���XE�ٿ�:]�X�@b%wƺ	4@�ڈ#��!?����5�@\�[_�ٿqT�5�@��!o�4@Вe���!?J G3+��@\�[_�ٿqT�5�@��!o�4@Вe���!?J G3+��@\�[_�ٿqT�5�@��!o�4@Вe���!?J G3+��@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@�B����ٿ]��I�@+�
��4@��C�!?�v���l�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@����ٿMu�ȍ[�@��B�4@@�t���!?��TQf�@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��$��ٿ溾h���@��4*4@���-��!?�f%/R��@��1���ٿqđ\��@�?�Y�4@�b��z�!?��5��@��1���ٿqđ\��@�?�Y�4@�b��z�!?��5��@��1���ٿqđ\��@�?�Y�4@�b��z�!?��5��@��1���ٿqđ\��@�?�Y�4@�b��z�!?��5��@��1���ٿqđ\��@�?�Y�4@�b��z�!?��5��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�� ��ٿ5�}���@v�<04@5r��!?%f{��@�0=K�ٿ,Z��@��B7� 4@���N�!?3Å��@`�1Uk�ٿ@��.���@�M�3@j�W�!?��P7��@`�1Uk�ٿ@��.���@�M�3@j�W�!?��P7��@��+y�ٿ"}���:�@*���
�3@��~ϐ!?O%-�p��@�N��ٿ��J����@��Gc*�3@��&�ߐ!?cyo����@r�B&�ٿ��q���@���+4@��8��!?芷;o��@r�B&�ٿ��q���@���+4@��8��!?芷;o��@g�ph͇ٿ�	ܔ��@6�ŏ�4@o��ە�!?n;��@g�ph͇ٿ�	ܔ��@6�ŏ�4@o��ە�!?n;��@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@���ٿ�R&X:��@�S4@��!?����s�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@=�K�ٿ����"��@�f`ƶ4@��E=��!?p���!�@� 6+\�ٿ������@�x�np4@K��׈�!?��C1w�@� 6+\�ٿ������@�x�np4@K��׈�!?��C1w�@� 6+\�ٿ������@�x�np4@K��׈�!?��C1w�@� 6+\�ٿ������@�x�np4@K��׈�!?��C1w�@� 6+\�ٿ������@�x�np4@K��׈�!?��C1w�@@��ٿ�3]����@�	���4@�hؐ�!?�}�X���@@��ٿ�3]����@�	���4@�hؐ�!?�}�X���@@��ٿ�3]����@�	���4@�hؐ�!?�}�X���@	�D��ٿ��Y֨�@ҵCgw4@����!?���	j�@	�D��ٿ��Y֨�@ҵCgw4@����!?���	j�@t�~�o�ٿ��%�?��@�����4@[S��!?�I.ǻ�@t�~�o�ٿ��%�?��@�����4@[S��!?�I.ǻ�@t�~�o�ٿ��%�?��@�����4@[S��!?�I.ǻ�@t�~�o�ٿ��%�?��@�����4@[S��!?�I.ǻ�@t�~�o�ٿ��%�?��@�����4@[S��!?�I.ǻ�@7Uxvb�ٿ��σ�]�@T�ɲ,4@�y[:�!?�=: j�@7Uxvb�ٿ��σ�]�@T�ɲ,4@�y[:�!?�=: j�@7Uxvb�ٿ��σ�]�@T�ɲ,4@�y[:�!?�=: j�@`��솈ٿI��[�O�@_f����3@vi�QƐ!?#�nԑ,�@`��솈ٿI��[�O�@_f����3@vi�QƐ!?#�nԑ,�@,ٿ0�ٿ9]�8ا�@��& R4@���!?�,FD}�@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�"���ٿ�O3TQ��@��f�
4@7Ʀ�!?)]ި���@�Cl}�ٿ"~�ܻ��@�p��4@�!&�!?5?�p�d�@�Cl}�ٿ"~�ܻ��@�p��4@�!&�!?5?�p�d�@99>��ٿ��4)�@|��� 4@<����!?�)�����@��oVD�ٿ 
���^�@�ЮJ�4@�'�/�!?�ݮ�z��@��oVD�ٿ 
���^�@�ЮJ�4@�'�/�!?�ݮ�z��@��oVD�ٿ 
���^�@�ЮJ�4@�'�/�!?�ݮ�z��@��oVD�ٿ 
���^�@�ЮJ�4@�'�/�!?�ݮ�z��@-� u�ٿ���1Q�@_��� 4@!����!?�/V��@-� u�ٿ���1Q�@_��� 4@!����!?�/V��@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@��{˷�ٿ�8�F��@��D�4@\K/��!?{Ƃ�>o�@[Xh�zٿ����@;�&�4@9y���!?���o�g�@�$e�^~ٿ�I����@1˱�i4@��R\�!?k�Xx���@�$e�^~ٿ�I����@1˱�i4@��R\�!?k�Xx���@�$e�^~ٿ�I����@1˱�i4@��R\�!?k�Xx���@��gk|ٿ��q��@nY04@����!?d��5|#�@��gk|ٿ��q��@nY04@����!?d��5|#�@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@w_T�X�ٿ�m!^:�@�R�q�4@iiܐ!?�9���@���ٿ�ZnI'`�@�-�4@�kx֤�!?�����@���ٿ�ZnI'`�@�-�4@�kx֤�!?�����@ui 	Çٿ�+o�I�@�}��4@���Z��!?E5^�-�@-�#�J�ٿ�����@�9$�a 4@��*U��!?�����@�p��͉ٿ�7�u��@�y�u@�3@D��/��!?_>���j�@�p��͉ٿ�7�u��@�y�u@�3@D��/��!?_>���j�@�c�P��ٿk�wP�)�@�,y�l4@����!?0��?���@�c�P��ٿk�wP�)�@�,y�l4@����!?0��?���@�c�P��ٿk�wP�)�@�,y�l4@����!?0��?���@�c�P��ٿk�wP�)�@�,y�l4@����!?0��?���@�c�P��ٿk�wP�)�@�,y�l4@����!?0��?���@�N��ٿ��Zu4A�@
�<�4@m� �!?'���^m�@�N��ٿ��Zu4A�@
�<�4@m� �!?'���^m�@�N��ٿ��Zu4A�@
�<�4@m� �!?'���^m�@�N��ٿ��Zu4A�@
�<�4@m� �!?'���^m�@�Gh�	�ٿ�^����@t���4@�ǭF�!?���c��@�Gh�	�ٿ�^����@t���4@�ǭF�!?���c��@��O��ٿ��)}3�@���4@����!?�N��A�@��O��ٿ��)}3�@���4@����!?�N��A�@��O��ٿ��)}3�@���4@����!?�N��A�@t��G��ٿzM�l��@g�y��4@t&��ِ!?hp�:W�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�2F �ٿf������@^|V4@�ȇt��!?�K�h	�@�3i,��ٿ�躜#:�@���}4@����Ԑ!?-��7m�@�3i,��ٿ�躜#:�@���}4@����Ԑ!?-��7m�@m\�}�ٿ޼ʹ�_�@�;���3@z&u�Ґ!?�i!�@m\�}�ٿ޼ʹ�_�@�;���3@z&u�Ґ!?�i!�@>���O�ٿmc��RU�@����3@��ڔ��!?猣-��@>���O�ٿmc��RU�@����3@��ڔ��!?猣-��@/�X؈ٿ㩆�	��@fp�]I4@�u���!?�?K�y�@/�X؈ٿ㩆�	��@fp�]I4@�u���!?�?K�y�@/�X؈ٿ㩆�	��@fp�]I4@�u���!?�?K�y�@/�X؈ٿ㩆�	��@fp�]I4@�u���!?�?K�y�@5�+G݅ٿQ��i�e�@]_��.4@Z����!?o���Y�@�] �ٿ����h�@wJ�! 4@R���Ґ!?�m=�%�@�] �ٿ����h�@wJ�! 4@R���Ґ!?�m=�%�@O[t%)�ٿ"�hNf��@W���4@�k��q�!?4�	 ��@O[t%)�ٿ"�hNf��@W���4@�k��q�!?4�	 ��@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@f�ZQƎٿ��&����@`��E4@;�B�!?�A�����@�)�-��ٿ/�Hն��@'��x�4@��[ϒ�!?��hf�_�@��ٿ �3�_��@�]��4@O�ʣ��!?�F��>�@��ٿ �3�_��@�]��4@O�ʣ��!?�F��>�@��ٿ �3�_��@�]��4@O�ʣ��!?�F��>�@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@B�#���ٿ-��$���@���4�4@�����!?�����@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@F�����ٿ/ܚU�'�@^L�f4@�����!?s-�!��@��GW�ٿu������@���4@�{�ې!?ϥ�}q�@Wg李ٿy�v���@Ԕ�C4@,	�I�!?uN���@s�wl�ٿD0[�/�@�c��y4@V�Q��!?D	a�S�@{^�L.�ٿ�;�w�Z�@9�-64@`Ч�!?����]�@{^�L.�ٿ�;�w�Z�@9�-64@`Ч�!?����]�@{^�L.�ٿ�;�w�Z�@9�-64@`Ч�!?����]�@�:� �ٿV��h,��@+�S�d4@�Q��ސ!?��Wu?��@�:� �ٿV��h,��@+�S�d4@�Q��ސ!?��Wu?��@�:� �ٿV��h,��@+�S�d4@�Q��ސ!?��Wu?��@��X��ٿ�gO�r�@"�0w14@�$����!?[�����@F�Ŝ7�ٿ��{���@p�ӥ4@-��@�!?����A�@���8�zٿ	�ˢx��@���φ4@��m�9�!?�oyJb�@���8�zٿ	�ˢx��@���φ4@��m�9�!?�oyJb�@���8�zٿ	�ˢx��@���φ4@��m�9�!?�oyJb�@���8�zٿ	�ˢx��@���φ4@��m�9�!?�oyJb�@���8�zٿ	�ˢx��@���φ4@��m�9�!?�oyJb�@ �Y[��ٿhd�]@��@�ڐ��4@��r�!?��DOi �@������ٿ@N=�H�@��K�&4@%�'�y�!?L�����@����ٿY}WZ�0�@�	:�4@s���#�!?t���*9�@����ٿY}WZ�0�@�	:�4@s���#�!?t���*9�@�.��}ٿ��D5��@|4�
4@τ���!?��-�1�@^2���ٿ`K����@�N94@�ݨ ސ!?%n|��	�@^2���ٿ`K����@�N94@�ݨ ސ!?%n|��	�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@�c�ٿ���D6��@_@��4@D֯�n�!?��3E13�@��/�i�ٿ�N�#�A�@{�6�P4@��f���!?׎���P�@����ٿ�������@~��6�4@���餐!?�!>7�@����ٿ�������@~��6�4@���餐!?�!>7�@����ٿ�������@~��6�4@���餐!?�!>7�@����ٿ�������@~��6�4@���餐!?�!>7�@����ٿ�������@~��6�4@���餐!?�!>7�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@L���ٿf�6\���@���b4@.Qs'�!?ؑ�Y$�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@�so�׆ٿ˩~2�)�@ݧ�Շ4@�_Vǐ!?v͊{�@7r���ٿ�9�k�@ ��B4@}�EV��!?Q-/tN0�@7r���ٿ�9�k�@ ��B4@}�EV��!?Q-/tN0�@7r���ٿ�9�k�@ ��B4@}�EV��!?Q-/tN0�@��/��ٿ��2gO��@��A��4@�����!?0ə�_�@��/��ٿ��2gO��@��A��4@�����!?0ə�_�@��/��ٿ��2gO��@��A��4@�����!?0ə�_�@��/��ٿ��2gO��@��A��4@�����!?0ə�_�@t؜���ٿ)�"`���@|� �V4@������!?�H��Y�@?���ٿ�PaM���@��}�=4@�S�Qg�!?�x��@?���ٿ�PaM���@��}�=4@�S�Qg�!?�x��@?���ٿ�PaM���@��}�=4@�S�Qg�!?�x��@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@d����ٿ�Gy�ߚ�@е�I;4@��ʐ!?�7�X�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@���ՀٿW���s�@�|��x4@a�.vŐ!?fd=J�=�@�j�[ӆٿi�A���@p�>H4@t��!��!?��0"&�@�j�[ӆٿi�A���@p�>H4@t��!��!?��0"&�@�j�[ӆٿi�A���@p�>H4@t��!��!?��0"&�@�j�[ӆٿi�A���@p�>H4@t��!��!?��0"&�@Ď��ٿ���FMJ�@/�KR�4@���X�!?S��*�@�$���ٿ���t���@0��� 4@P�W��!?6�Qa�@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@7���|ٿ�Гg6��@|x0�c4@� &��!?��	���@e�Sbm�ٿ���Z�5�@r�-�4@ y6ؐ�!?~(0q�@e�Sbm�ٿ���Z�5�@r�-�4@ y6ؐ�!?~(0q�@	C��ٿ��sq�@A)��4@*����!?c�����@	C��ٿ��sq�@A)��4@*����!?c�����@	C��ٿ��sq�@A)��4@*����!?c�����@	C��ٿ��sq�@A)��4@*����!?c�����@���Jڄٿv/+3Ų�@�]J>4@�$���!?DQ@�N]�@[�	�ٿpy\�@�~��4@m8c��!?f�1�R�@[�	�ٿpy\�@�~��4@m8c��!?f�1�R�@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@앸�*�ٿ�~���@��d��4@e�>��!?���Q��@ R�*׈ٿ��
j]�@ٌ]�G4@̷<��!?`�GN���@ R�*׈ٿ��
j]�@ٌ]�G4@̷<��!?`�GN���@�y�S�ٿ<}]��!�@g�' 4@���G�!?/�YZa�@�5c4�ٿ��I)m�@��f^�4@z���!�!?UkSc��@���ٿ��29��@���a�4@ c�!?[\��d�@���ٿ��29��@���a�4@ c�!?[\��d�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�_��ٿ�Ӎ��V�@0�BXs4@��f��!?,>h��Q�@�jOh��ٿ%��+^��@�P�4@Iq���!?�+����@�jOh��ٿ%��+^��@�P�4@Iq���!?�+����@�jOh��ٿ%��+^��@�P�4@Iq���!?�+����@�$���ٿ	�]�=�@�Yfd4@���M��!?������@�$���ٿ	�]�=�@�Yfd4@���M��!?������@�$���ٿ	�]�=�@�Yfd4@���M��!?������@426��ٿv��ᛢ�@$�x�.4@w�BX��!?.�fgQr�@426��ٿv��ᛢ�@$�x�.4@w�BX��!?.�fgQr�@426��ٿv��ᛢ�@$�x�.4@w�BX��!?.�fgQr�@S�G��ٿ8��Q��@�Ŝ4@����!?VN�7�@i��Z��ٿ���ڂ�@�U}r4@-����!?�2��n�@i��Z��ٿ���ڂ�@�U}r4@-����!?�2��n�@i��Z��ٿ���ڂ�@�U}r4@-����!?�2��n�@i��Z��ٿ���ڂ�@�U}r4@-����!?�2��n�@i��Z��ٿ���ڂ�@�U}r4@-����!?�2��n�@=D�9׋ٿ�`�
��@����4@�aH~�!?������@=D�9׋ٿ�`�
��@����4@�aH~�!?������@���ٿ=�^,��@G�i�4@�Eu�ʐ!?���v�(�@���ٿ=�^,��@G�i�4@�Eu�ʐ!?���v�(�@���ٿ=�^,��@G�i�4@�Eu�ʐ!?���v�(�@���ٿ=�^,��@G�i�4@�Eu�ʐ!?���v�(�@�f���ٿ�qi(d��@��%�4@U��:��!?)�t��@�f���ٿ�qi(d��@��%�4@U��:��!?)�t��@���%�ٿ\��.bP�@�.�4@aE����!?h�Z�F��@���%�ٿ\��.bP�@�.�4@aE����!?h�Z�F��@r &��ٿ����}�@f���F4@�wE֐!?4�M"��@r &��ٿ����}�@f���F4@�wE֐!?4�M"��@!�%K�ٿ���"�@�嬫|4@��9yd�!?(�UpZM�@!�%K�ٿ���"�@�嬫|4@��9yd�!?(�UpZM�@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@yƾɦ�ٿ��Ep�@�O4�#4@3a�א!?~`�J��@!�t
�ٿo�~�j<�@Yx*�4@��')��!?\ӊ�@!�t
�ٿo�~�j<�@Yx*�4@��')��!?\ӊ�@�-W�&�ٿ̯�&Kf�@e�%�E4@f ���!?�v� �@�-W�&�ٿ̯�&Kf�@e�%�E4@f ���!?�v� �@�-W�&�ٿ̯�&Kf�@e�%�E4@f ���!?�v� �@�-W�&�ٿ̯�&Kf�@e�%�E4@f ���!?�v� �@�-W�&�ٿ̯�&Kf�@e�%�E4@f ���!?�v� �@v��N�ٿ��~W[�@пH!�4@f���!?����lR�@v��N�ٿ��~W[�@пH!�4@f���!?����lR�@v��N�ٿ��~W[�@пH!�4@f���!?����lR�@v��N�ٿ��~W[�@пH!�4@f���!?����lR�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@�jo`�ٿ4S�~�@�P(:*4@M�0�ؐ!?�]�{"�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@������ٿ�G]U_��@�R��4@�Z����!?�����\�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@n�|��ٿ�6��ȃ�@=>P�4@������!?ʺ|ax�@U�u#�ٿ4D�1�@��q�4@�'Pɑ�!?�g%5�0�@���ٿes�OD�@���H4@��Ɛ!?�T�#�@���،ٿ�焩��@����4@MQ���!?��U�u�@���،ٿ�焩��@����4@MQ���!?��U�u�@ ��$�ٿ���t:��@_D��4@y�JTi�!?��j,�b�@ ��$�ٿ���t:��@_D��4@y�JTi�!?��j,�b�@ ��$�ٿ���t:��@_D��4@y�JTi�!?��j,�b�@ ��$�ٿ���t:��@_D��4@y�JTi�!?��j,�b�@ ��$�ٿ���t:��@_D��4@y�JTi�!?��j,�b�@~���m�ٿ��业�@��	��4@`�~�!?0��6��@~���m�ٿ��业�@��	��4@`�~�!?0��6��@�w~�{ٿ��@���@���4@��ԙ�!?�)"����@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@���xٿ�S3�[��@���,`4@�Nm���!?x�6�m�@��xٿ� ��u�@H��ɖ4@2M���!?�}�^���@'���r|ٿ�j��@xF��]4@Ǟ^)��!?V	"b���@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@�@��r�ٿ`��M_�@!�a_�4@#���!?�L}=pT�@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@N�q�ٿ����� �@ n��24@HX�א!?C#����@�@���ٿ"��Q�5�@�G�C�4@Q3���!?��4��@�@���ٿ"��Q�5�@�G�C�4@Q3���!?��4��@�@���ٿ"��Q�5�@�G�C�4@Q3���!?��4��@�@���ٿ"��Q�5�@�G�C�4@Q3���!?��4��@�@���ٿ"��Q�5�@�G�C�4@Q3���!?��4��@] ��i�ٿ'���0��@��A8� 4@T
>��!?_w����@] ��i�ٿ'���0��@��A8� 4@T
>��!?_w����@˦l�}ٿ(�Gr���@�Ο� 4@U�n��!?���t���@R'KÓٿ݉��M�@FB�-m4@T����!?�I�B�@R'KÓٿ݉��M�@FB�-m4@T����!?�I�B�@R'KÓٿ݉��M�@FB�-m4@T����!?�I�B�@R'KÓٿ݉��M�@FB�-m4@T����!?�I�B�@R���z�ٿ^&���@��g��4@�5Cy�!?�2l��@R���z�ٿ^&���@��g��4@�5Cy�!?�2l��@R���z�ٿ^&���@��g��4@�5Cy�!?�2l��@R���z�ٿ^&���@��g��4@�5Cy�!?�2l��@R���z�ٿ^&���@��g��4@�5Cy�!?�2l��@;C�hҌٿR"\�b��@=�[ 4@V��wk�!?A�
��@;C�hҌٿR"\�b��@=�[ 4@V��wk�!?A�
��@;C�hҌٿR"\�b��@=�[ 4@V��wk�!?A�
��@:l�lg�ٿc|Rm��@�"<�4@4�jb�!?�㩵0<�@�W]��ٿb �3w�@�H</�3@�u��0�!?�N`W�@�W]��ٿb �3w�@�H</�3@�u��0�!?�N`W�@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@�l�ؘ�ٿ��1D��@�~�C 4@Fs=���!?�;FC��@}q���ٿAK���P�@Җ�4@aƢ֐!?������@}q���ٿAK���P�@Җ�4@aƢ֐!?������@}q���ٿAK���P�@Җ�4@aƢ֐!?������@}q���ٿAK���P�@Җ�4@aƢ֐!?������@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@n��L��ٿ�K���@ѡ��14@��,w��!?��k��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@u:���ٿP<�X[�@��ah4@�>�EȐ!?��gu ��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@5��9�ٿ��;'�@����4@� A��!?!�!�^��@A��(T�ٿB4���@ugl��4@О�u�!?0�����@�?�R
�ٿ)����D�@j��! 4@Ej$���!?=5BG(�@�?�R
�ٿ)����D�@j��! 4@Ej$���!?=5BG(�@�?�R
�ٿ)����D�@j��! 4@Ej$���!?=5BG(�@�?�R
�ٿ)����D�@j��! 4@Ej$���!?=5BG(�@�?�R
�ٿ)����D�@j��! 4@Ej$���!?=5BG(�@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@ظA�;�ٿ��)��7�@�*��4@�r"@�!?��|��@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@̞�l��ٿ{�����@,���4@���
�!?r�����@/�k%\ٿL������@��~"4@e�ۊg�!?��j�0��@/�k%\ٿL������@��~"4@e�ۊg�!?��j�0��@��^�c�ٿ!�x]���@J��4@���XU�!?B�	c��@��^�c�ٿ!�x]���@J��4@���XU�!?B�	c��@��^�c�ٿ!�x]���@J��4@���XU�!?B�	c��@��Z�ٿ��u���@���C4@pXFT�!?���[jA�@��=�ٿ��ǳ��@\�M��	4@��9�/�!?�>�ߓ�@��=�ٿ��ǳ��@\�M��	4@��9�/�!?�>�ߓ�@��=�ٿ��ǳ��@\�M��	4@��9�/�!?�>�ߓ�@��=�ٿ��ǳ��@\�M��	4@��9�/�!?�>�ߓ�@Y��G��ٿJ2�zr�@��B]4@�
;8�!?������@Y��G��ٿJ2�zr�@��B]4@�
;8�!?������@Y��G��ٿJ2�zr�@��B]4@�
;8�!?������@��K�-}ٿ������@Z�L��4@�o~�?�!?U|tA1�@��K�-}ٿ������@Z�L��4@�o~�?�!?U|tA1�@��K�-}ٿ������@Z�L��4@�o~�?�!?U|tA1�@��K�-}ٿ������@Z�L��4@�o~�?�!?U|tA1�@��K�-}ٿ������@Z�L��4@�o~�?�!?U|tA1�@q��Grٿ4�
����@ViB�	4@�'���!?�BL}ת�@q��Grٿ4�
����@ViB�	4@�'���!?�BL}ת�@q��Grٿ4�
����@ViB�	4@�'���!?�BL}ת�@{�G�RuٿD^����@G}�Ԛ4@����!?�N_����@{�G�RuٿD^����@G}�Ԛ4@����!?�N_����@{�G�RuٿD^����@G}�Ԛ4@����!?�N_����@{�G�RuٿD^����@G}�Ԛ4@����!?�N_����@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@=+*wٿa?��M��@�V�k?	4@�����!? m���}�@�V�K�~ٿ�Q�#r�@`��m�
4@���!?��&PiK�@�V�K�~ٿ�Q�#r�@`��m�
4@���!?��&PiK�@�g q�{ٿ�mw{�j�@�=�U�
4@~��)�!?�J�W��@�g q�{ٿ�mw{�j�@�=�U�
4@~��)�!?�J�W��@�g q�{ٿ�mw{�j�@�=�U�
4@~��)�!?�J�W��@�g q�{ٿ�mw{�j�@�=�U�
4@~��)�!?�J�W��@�H��^}ٿ��u��v�@v�� �4@Z�*}*�!?{m�$��@�H��^}ٿ��u��v�@v�� �4@Z�*}*�!?{m�$��@�w�n}ٿ��� ��@�t�]�4@A�L���!?�Sb�Ҽ�@�YB[�ٿ��i��@����4@��MV�!?%H���@�YB[�ٿ��i��@����4@��MV�!?%H���@[;��ٿ�^ۨ���@���4@hPI,q�!?]�N��@[;��ٿ�^ۨ���@���4@hPI,q�!?]�N��@[;��ٿ�^ۨ���@���4@hPI,q�!?]�N��@[;��ٿ�^ۨ���@���4@hPI,q�!?]�N��@�*��ٿ�ita�@��}�4@��I�Ȑ!?����@��s�ٿ�1�Xm�@g<�� 4@T�yƐ!?�hP�@���~ٿ��0�H��@n}�,�4@}{t��!?Iu� �@���~ٿ��0�H��@n}�,�4@}{t��!?Iu� �@�̵I��ٿ����@����T4@w0@#D�!?S�(�G�@�̵I��ٿ����@����T4@w0@#D�!?S�(�G�@߿��*�ٿ`7��@ ��d4@��B�}�!?��g�_��@߿��*�ٿ`7��@ ��d4@��B�}�!?��g�_��@߿��*�ٿ`7��@ ��d4@��B�}�!?��g�_��@߿��*�ٿ`7��@ ��d4@��B�}�!?��g�_��@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�*ZJ�ٿl�&��@3���K4@;r�ڐ!?o�0�ij�@�JPk_�ٿ�6���@<O�C4@��
Ȑ!?jx�c|�@���O��ٿ��ޞ��@$��q4@ �ћ�!??�h/��@���O��ٿ��ޞ��@$��q4@ �ћ�!??�h/��@���O��ٿ��ޞ��@$��q4@ �ћ�!??�h/��@���O��ٿ��ޞ��@$��q4@ �ћ�!??�h/��@���O��ٿ��ޞ��@$��q4@ �ћ�!??�h/��@���»�ٿ�DW���@ ���4@�5�緐!?��t�>�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@=�}ςٿ��+��_�@�C�z�4@��̾��!?�V�S�-�@� ʖ;�ٿ�Jx���@�@��4@ЏD�R�!?�P��J�@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@P5�ٿ������@��e�	4@+.�А!?�-��}��@�~F���ٿ�j:���@Z�4@k;���!?׍f�.�@�~F���ٿ�j:���@Z�4@k;���!?׍f�.�@�~F���ٿ�j:���@Z�4@k;���!?׍f�.�@�~F���ٿ�j:���@Z�4@k;���!?׍f�.�@�~F���ٿ�j:���@Z�4@k;���!?׍f�.�@��wx�ٿ��h[r��@_/8�4@����!?��3��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@�9OZ�ٿP�@h���@h]�J�4@h��@��!?��'H��@5/te�ٿ13-����@ޚ�c4@F脐!?�����@5/te�ٿ13-����@ޚ�c4@F脐!?�����@¸�4�ٿ�(����@fP�qc4@�!~Ɛ!?��I�-�@¸�4�ٿ�(����@fP�qc4@�!~Ɛ!?��I�-�@¸�4�ٿ�(����@fP�qc4@�!~Ɛ!?��I�-�@���w�ٿp(�B�@h:���4@�����!?`��$c��@.�����ٿo;�U�@�6I�4@�=Y��!?*ˤ��@.�����ٿo;�U�@�6I�4@�=Y��!?*ˤ��@.�����ٿo;�U�@�6I�4@�=Y��!?*ˤ��@.�����ٿo;�U�@�6I�4@�=Y��!?*ˤ��@���^�ٿ@aIhܘ�@t�!;J4@�1�9!?1U�Lɓ�@���^�ٿ@aIhܘ�@t�!;J4@�1�9!?1U�Lɓ�@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@�򟄍�ٿ�!��p��@�/6�4@ޢ�!?1d>4���@E�0���ٿ�;AT���@sR��4@�:ZQ��!?
���Jw�@E�0���ٿ�;AT���@sR��4@�:ZQ��!?
���Jw�@E�0���ٿ�;AT���@sR��4@�:ZQ��!?
���Jw�@��.��ٿ��kx��@�ȝ�4@|��2��!?	�4�)��@��.��ٿ��kx��@�ȝ�4@|��2��!?	�4�)��@��.��ٿ��kx��@�ȝ�4@|��2��!?	�4�)��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@��A�ٿ���^��@6B��4@��nߐ!?��M`��@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@�ܕ5�ٿP�ȓ��@U(|@�4@.q��Ő!?�0��4|�@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@-Z�|ٿ�vp���@�1��M4@��^��!?�'8@��@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@ �T���ٿ���Է��@Q��[�4@��R%��!?x5����@N�J|��ٿ�
Hre�@���4@�?�_|�!?x��Ip�@N�J|��ٿ�
Hre�@���4@�?�_|�!?x��Ip�@N�J|��ٿ�
Hre�@���4@�?�_|�!?x��Ip�@N�J|��ٿ�
Hre�@���4@�?�_|�!?x��Ip�@N�J|��ٿ�
Hre�@���4@�?�_|�!?x��Ip�@��l�ٿ�.O��v�@w�.�4@8^kw��!?^b�<���@��l�ٿ�.O��v�@w�.�4@8^kw��!?^b�<���@��l�ٿ�.O��v�@w�.�4@8^kw��!?^b�<���@��l�ٿ�.O��v�@w�.�4@8^kw��!?^b�<���@��l�ٿ�.O��v�@w�.�4@8^kw��!?^b�<���@���ѝ|ٿψ�m
�@�WX(�4@6Kdd��!?�Rr���@���ѝ|ٿψ�m
�@�WX(�4@6Kdd��!?�Rr���@���ѝ|ٿψ�m
�@�WX(�4@6Kdd��!?�Rr���@���ѝ|ٿψ�m
�@�WX(�4@6Kdd��!?�Rr���@7�c3��ٿ��h����@=8ڈ�4@��~͐!?���@7�c3��ٿ��h����@=8ڈ�4@��~͐!?���@7�c3��ٿ��h����@=8ڈ�4@��~͐!?���@7�c3��ٿ��h����@=8ڈ�4@��~͐!?���@7�c3��ٿ��h����@=8ڈ�4@��~͐!?���@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@b����ٿya��z]�@����N4@��S�!?�Q�8J*�@�_$H�ٿ��^C�@g����4@� ��!?[�l���@�_$H�ٿ��^C�@g����4@� ��!?[�l���@�����ٿ��2x��@ڏG��4@�x�1��!?0]�����@�����ٿ��2x��@ڏG��4@�x�1��!?0]�����@�����ٿ��2x��@ڏG��4@�x�1��!?0]�����@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@uܨCԊٿw�'��#�@�>��4@Asn��!?�qݮN)�@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@��M�	�ٿ�)����@J�ڪ4@��r!?Z� ���@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@���l�ٿ~�B����@ߜwE4@�֯��!?�g�ʋ��@�ΚN��ٿ{����@��54@#�_�z�!?��?�@�ΚN��ٿ{����@��54@#�_�z�!?��?�@�ΚN��ٿ{����@��54@#�_�z�!?��?�@�ΚN��ٿ{����@��54@#�_�z�!?��?�@�(+(��ٿ���2�I�@�*���4@�k^g��!?E�f�3j�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@�!��ٿ������@lvͼ}4@�v���!?\�Q!�@n~���ٿ����@�W�4@UR,��!?�I�����@n~���ٿ����@�W�4@UR,��!?�I�����@n~���ٿ����@�W�4@UR,��!?�I�����@n~���ٿ����@�W�4@UR,��!?�I�����@n~���ٿ����@�W�4@UR,��!?�I�����@5J�荊ٿ�N*��x�@��#�3@��y��!?<�����@�c�bȇٿ��Χ���@�O�Rz4@|>T�:�!?ft7�Ȉ�@�c�bȇٿ��Χ���@�O�Rz4@|>T�:�!?ft7�Ȉ�@��L�U�ٿ��q?��@cl��4@�]q�!?�"ǳL|�@��L�U�ٿ��q?��@cl��4@�]q�!?�"ǳL|�@��L�U�ٿ��q?��@cl��4@�]q�!?�"ǳL|�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@��O��ٿ=������@�۲ 4@�)X�!?�*r½�@���o�ٿWM�+ ��@p%�g4@�s���!?#�L�7�@���o�ٿWM�+ ��@p%�g4@�s���!?#�L�7�@�l�щٿ�67��.�@�r�.� 4@��Q��!?2<�Y9��@����?}ٿ�&㢪�@��K�k4@��n��!??7i�@����?}ٿ�&㢪�@��K�k4@��n��!??7i�@��o"(�ٿ��޵���@m�O��	4@��w���!?#~��N�@��o"(�ٿ��޵���@m�O��	4@��w���!?#~��N�@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@g��ɳ�ٿ��|h��@�=Ze4@��ʦ��!?�Ϡ��@;���ٿ��H���@c�#S=4@_��$�!?4�Y���@Ix~��ٿ��Ej�=�@�:g�4@:����!?�^�U��@����ٿ{~���@���4@t�i��!?U�b��s�@��_ �ٿh��Q��@�Q�*4@�L�.��!?"~��Ie�@��_ �ٿh��Q��@�Q�*4@�L�.��!?"~��Ie�@��_ �ٿh��Q��@�Q�*4@�L�.��!?"~��Ie�@��_ �ٿh��Q��@�Q�*4@�L�.��!?"~��Ie�@�d͊Èٿ{t�9��@s��� 
4@����!?�Do��@"�B��ٿⵧfR��@�|�o4@��?@�!?,����@"�B��ٿⵧfR��@�|�o4@��?@�!?,����@"�B��ٿⵧfR��@�|�o4@��?@�!?,����@(� ��ٿ`f:�#c�@�I���4@���P��!?�{�4Z�@(� ��ٿ`f:�#c�@�I���4@���P��!?�{�4Z�@(� ��ٿ`f:�#c�@�I���4@���P��!?�{�4Z�@(� ��ٿ`f:�#c�@�I���4@���P��!?�{�4Z�@(� ��ٿ`f:�#c�@�I���4@���P��!?�{�4Z�@�
(�%}ٿQJb��@A�v]�4@��Oq�!?4�:yro�@�
(�%}ٿQJb��@A�v]�4@��Oq�!?4�:yro�@�
(�%}ٿQJb��@A�v]�4@��Oq�!?4�:yro�@�T`�ٿ%�;���@s�
1�4@W��!u�!?k6��@�T`�ٿ%�;���@s�
1�4@W��!u�!?k6��@�T`�ٿ%�;���@s�
1�4@W��!u�!?k6��@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@������ٿV����@�S��4@��� ��!?/�v��D�@�p[谇ٿٯ�ft9�@T
ڞ24@�H?�	�!?G_�~���@�p[谇ٿٯ�ft9�@T
ڞ24@�H?�	�!?G_�~���@�p[谇ٿٯ�ft9�@T
ڞ24@�H?�	�!?G_�~���@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@�2�w��ٿf�5O�@�1\��4@zN6H͐!?�	�4�1�@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@eO��x�ٿ�o;��@����
4@�T� �!?�o@�c��@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@)��~�ٿل�w��@�T��x4@rR�*�!?�����;�@9�WՑٿ<�Ð��@qXg4@0���!?�������@9�WՑٿ<�Ð��@qXg4@0���!?�������@9�WՑٿ<�Ð��@qXg4@0���!?�������@9�WՑٿ<�Ð��@qXg4@0���!?�������@9�WՑٿ<�Ð��@qXg4@0���!?�������@9�WՑٿ<�Ð��@qXg4@0���!?�������@L�{,ٿИ�P�@7AP�4@j�
��!?	=J���@L�{,ٿИ�P�@7AP�4@j�
��!?	=J���@L�{,ٿИ�P�@7AP�4@j�
��!?	=J���@L�{,ٿИ�P�@7AP�4@j�
��!?	=J���@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@��x�S�ٿ;8�w��@�W�4@�BQ�n�!?P �����@#�nž�ٿ�<9z\�@���˼4@���G��!?�2�5`�@��򑏆ٿ��3�@�e���4@�N79�!?
iqW���@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�,O�ٿ-���%��@~V+E4@c�V���!?��yڢ[�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@�媨t�ٿ�f'r��@TΏ�4@���!?WJa�R�@����r�ٿ�KlަZ�@��q4@НH,�!?�v!��@����r�ٿ�KlަZ�@��q4@НH,�!?�v!��@_n�r��ٿ]X�gaX�@�a蚛	4@ū�f�!?��DH��@_n�r��ٿ]X�gaX�@�a蚛	4@ū�f�!?��DH��@_n�r��ٿ]X�gaX�@�a蚛	4@ū�f�!?��DH��@<BI��ٿ�R=
�@�^TWA4@@¾�!?� �R{k�@<BI��ٿ�R=
�@�^TWA4@@¾�!?� �R{k�@<BI��ٿ�R=
�@�^TWA4@@¾�!?� �R{k�@�z��~ٿ�G�
v��@�����4@���]�!?M�"Xr�@�z��~ٿ�G�
v��@�����4@���]�!?M�"Xr�@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@F�W,}ٿ��|��@�^zʣ4@0u�r�!?a�+h��@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@T j.5�ٿ���b���@2F�
4@��4�h�!?�������@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@_�'��ٿ^���H��@# ӹ*4@��\Ẑ!?4�}l�@T�4�ٿ��t	c�@�1�Μ4@cTh��!?��KVc�@T�4�ٿ��t	c�@�1�Μ4@cTh��!?��KVc�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@%^�*n�ٿ�a�7��@󾇼?4@K�,�!?Ρ�?D�@